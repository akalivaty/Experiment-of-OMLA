//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 0 0 1 0 1 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n203), .A2(KEYINPUT96), .A3(KEYINPUT16), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT96), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n205), .B1(new_n206), .B2(G1gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n202), .A2(new_n204), .A3(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n208), .B1(G1gat), .B2(new_n202), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT97), .B1(new_n202), .B2(G1gat), .ZN(new_n210));
  INV_X1    g009(.A(G8gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n209), .B(new_n212), .ZN(new_n213));
  XOR2_X1   g012(.A(G43gat), .B(G50gat), .Z(new_n214));
  INV_X1    g013(.A(KEYINPUT15), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n216), .B(KEYINPUT94), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n214), .A2(new_n215), .ZN(new_n218));
  INV_X1    g017(.A(G29gat), .ZN(new_n219));
  AND3_X1   g018(.A1(new_n219), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT14), .B(G29gat), .ZN(new_n221));
  INV_X1    g020(.A(G36gat), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NOR3_X1   g022(.A1(new_n217), .A2(new_n218), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n218), .A2(new_n223), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n225), .B(KEYINPUT93), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT95), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT17), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n229), .A2(KEYINPUT17), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n213), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT98), .ZN(new_n235));
  INV_X1    g034(.A(new_n227), .ZN(new_n236));
  AOI22_X1  g035(.A1(new_n234), .A2(new_n235), .B1(new_n213), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G229gat), .A2(G233gat), .ZN(new_n238));
  XOR2_X1   g037(.A(new_n238), .B(KEYINPUT99), .Z(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n213), .ZN(new_n241));
  INV_X1    g040(.A(new_n233), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n229), .A2(KEYINPUT17), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT98), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n237), .A2(new_n240), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT18), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n237), .A2(new_n245), .A3(KEYINPUT18), .A4(new_n240), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n227), .B(new_n213), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n239), .B(KEYINPUT13), .Z(new_n251));
  OR2_X1    g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n248), .A2(new_n249), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT92), .ZN(new_n254));
  XNOR2_X1  g053(.A(G113gat), .B(G141gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(G197gat), .ZN(new_n256));
  XOR2_X1   g055(.A(KEYINPUT11), .B(G169gat), .Z(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XOR2_X1   g057(.A(new_n258), .B(KEYINPUT12), .Z(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n253), .A2(new_n254), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n260), .B1(new_n253), .B2(new_n254), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT36), .ZN(new_n266));
  NAND2_X1  g065(.A1(G227gat), .A2(G233gat), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(G120gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(G113gat), .ZN(new_n270));
  INV_X1    g069(.A(G113gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(G120gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT1), .ZN(new_n274));
  XNOR2_X1  g073(.A(G127gat), .B(G134gat), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n273), .B(new_n274), .C1(new_n275), .C2(KEYINPUT74), .ZN(new_n276));
  INV_X1    g075(.A(G127gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(G134gat), .ZN(new_n278));
  INV_X1    g077(.A(G134gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(G127gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n274), .A2(KEYINPUT74), .ZN(new_n282));
  XNOR2_X1  g081(.A(G113gat), .B(G120gat), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n281), .B(new_n282), .C1(new_n283), .C2(KEYINPUT1), .ZN(new_n284));
  AND2_X1   g083(.A1(new_n276), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT24), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT65), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT65), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n286), .A2(new_n290), .A3(new_n287), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND4_X1  g091(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT64), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT66), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n297), .B1(G183gat), .B2(G190gat), .ZN(new_n298));
  INV_X1    g097(.A(G183gat), .ZN(new_n299));
  INV_X1    g098(.A(G190gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n299), .A2(new_n300), .A3(KEYINPUT66), .ZN(new_n301));
  AND4_X1   g100(.A1(new_n293), .A2(new_n296), .A3(new_n298), .A4(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G169gat), .A2(G176gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT23), .ZN(new_n304));
  INV_X1    g103(.A(G169gat), .ZN(new_n305));
  INV_X1    g104(.A(G176gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT68), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(new_n306), .ZN(new_n310));
  NAND2_X1  g109(.A1(KEYINPUT68), .A2(G176gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n310), .A2(KEYINPUT23), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n305), .A2(KEYINPUT67), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT67), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G169gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n308), .B1(new_n312), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT69), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n292), .A2(new_n302), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OAI211_X1 g118(.A(KEYINPUT69), .B(new_n308), .C1(new_n312), .C2(new_n316), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT25), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT25), .ZN(new_n322));
  INV_X1    g121(.A(new_n307), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n322), .B1(new_n323), .B2(KEYINPUT23), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n288), .B(new_n294), .C1(G183gat), .C2(G190gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n324), .A2(new_n308), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT70), .B1(new_n321), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n317), .A2(new_n318), .ZN(new_n329));
  AND3_X1   g128(.A1(new_n296), .A2(new_n298), .A3(new_n301), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n330), .A2(new_n292), .A3(new_n293), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n329), .A2(new_n331), .A3(new_n320), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(new_n322), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT70), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(new_n334), .A3(new_n326), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n328), .A2(new_n335), .ZN(new_n336));
  AOI22_X1  g135(.A1(new_n323), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n337));
  OR2_X1    g136(.A1(new_n323), .A2(KEYINPUT26), .ZN(new_n338));
  INV_X1    g137(.A(new_n303), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT28), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT27), .ZN(new_n342));
  OAI21_X1  g141(.A(KEYINPUT71), .B1(new_n342), .B2(G183gat), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT71), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n344), .A2(new_n299), .A3(KEYINPUT27), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n343), .A2(new_n345), .A3(new_n300), .ZN(new_n346));
  OR2_X1    g145(.A1(KEYINPUT72), .A2(KEYINPUT27), .ZN(new_n347));
  NAND2_X1  g146(.A1(KEYINPUT72), .A2(KEYINPUT27), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n299), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n341), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT27), .B(G183gat), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n351), .A2(KEYINPUT28), .A3(new_n300), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT73), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT73), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n350), .A2(new_n355), .A3(new_n352), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n340), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n285), .B1(new_n336), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n276), .A2(new_n284), .ZN(new_n360));
  AOI211_X1 g159(.A(new_n360), .B(new_n357), .C1(new_n328), .C2(new_n335), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n268), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT32), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT75), .B(KEYINPUT33), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  XOR2_X1   g165(.A(G15gat), .B(G43gat), .Z(new_n367));
  XNOR2_X1  g166(.A(G71gat), .B(G99gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n363), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n369), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n362), .B(KEYINPUT32), .C1(new_n365), .C2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n334), .B1(new_n333), .B2(new_n326), .ZN(new_n374));
  AOI211_X1 g173(.A(KEYINPUT70), .B(new_n327), .C1(new_n332), .C2(new_n322), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n358), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n360), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n358), .B(new_n285), .C1(new_n374), .C2(new_n375), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n377), .A2(new_n267), .A3(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(KEYINPUT76), .B(KEYINPUT34), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(KEYINPUT76), .A2(KEYINPUT34), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n377), .A2(new_n267), .A3(new_n378), .A4(new_n382), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n373), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n372), .A3(new_n384), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT77), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT77), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n370), .A2(new_n384), .A3(new_n389), .A4(new_n372), .ZN(new_n390));
  AND3_X1   g189(.A1(new_n388), .A2(KEYINPUT78), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT78), .B1(new_n388), .B2(new_n390), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n266), .B(new_n386), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(G155gat), .A2(G162gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT2), .ZN(new_n395));
  INV_X1    g194(.A(G141gat), .ZN(new_n396));
  INV_X1    g195(.A(G148gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(G141gat), .A2(G148gat), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n395), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT80), .ZN(new_n401));
  XNOR2_X1  g200(.A(G155gat), .B(G162gat), .ZN(new_n402));
  AND3_X1   g201(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n402), .B1(new_n400), .B2(new_n401), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT4), .B1(new_n405), .B2(new_n360), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n400), .A2(new_n401), .ZN(new_n407));
  INV_X1    g206(.A(new_n402), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT4), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(new_n285), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n406), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT3), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT81), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n360), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n409), .A2(KEYINPUT3), .A3(new_n410), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n276), .A2(new_n284), .A3(KEYINPUT81), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n416), .A2(new_n418), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT5), .ZN(new_n422));
  NAND2_X1  g221(.A1(G225gat), .A2(G233gat), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n414), .A2(new_n421), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT82), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n406), .A2(new_n425), .A3(new_n413), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n285), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n427), .A2(KEYINPUT82), .A3(KEYINPUT4), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n426), .A2(new_n428), .A3(new_n421), .A4(new_n423), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n418), .A2(new_n405), .A3(new_n420), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n427), .ZN(new_n431));
  INV_X1    g230(.A(new_n423), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n422), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n429), .A2(KEYINPUT83), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT83), .B1(new_n429), .B2(new_n433), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n424), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(G1gat), .B(G29gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n437), .B(KEYINPUT0), .ZN(new_n438));
  XNOR2_X1  g237(.A(G57gat), .B(G85gat), .ZN(new_n439));
  XOR2_X1   g238(.A(new_n438), .B(new_n439), .Z(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT6), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n424), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n433), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT83), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n429), .A2(KEYINPUT83), .A3(new_n433), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n445), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT6), .B1(new_n450), .B2(new_n440), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n444), .B1(new_n442), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(G197gat), .B(G204gat), .ZN(new_n454));
  INV_X1    g253(.A(G211gat), .ZN(new_n455));
  INV_X1    g254(.A(G218gat), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n454), .B1(KEYINPUT22), .B2(new_n457), .ZN(new_n458));
  XOR2_X1   g257(.A(G211gat), .B(G218gat), .Z(new_n459));
  XNOR2_X1  g258(.A(new_n458), .B(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n358), .B1(new_n321), .B2(new_n327), .ZN(new_n462));
  NAND2_X1  g261(.A1(G226gat), .A2(G233gat), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT29), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n464), .B1(new_n376), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT79), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n357), .B1(new_n328), .B2(new_n335), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n463), .B1(new_n470), .B2(KEYINPUT29), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n471), .A2(KEYINPUT79), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n461), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n470), .A2(new_n464), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n462), .A2(new_n466), .A3(new_n463), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n460), .ZN(new_n477));
  XNOR2_X1  g276(.A(G8gat), .B(G36gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(G64gat), .B(G92gat), .ZN(new_n479));
  XOR2_X1   g278(.A(new_n478), .B(new_n479), .Z(new_n480));
  NAND3_X1  g279(.A1(new_n473), .A2(new_n477), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT30), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n473), .A2(KEYINPUT30), .A3(new_n477), .A4(new_n480), .ZN(new_n484));
  INV_X1    g283(.A(new_n480), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n471), .A2(KEYINPUT79), .B1(new_n464), .B2(new_n462), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n467), .A2(new_n468), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n460), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n477), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n485), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n453), .A2(new_n483), .A3(new_n484), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n460), .A2(new_n466), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n411), .B1(new_n492), .B2(new_n415), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n460), .B1(new_n416), .B2(new_n466), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(G78gat), .B(G106gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n495), .B(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(G228gat), .A2(G233gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n498), .B(G22gat), .ZN(new_n499));
  XOR2_X1   g298(.A(KEYINPUT31), .B(G50gat), .Z(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n497), .A2(new_n501), .ZN(new_n503));
  OR2_X1    g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n491), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n388), .A2(new_n390), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(new_n386), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT36), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n393), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n490), .A2(new_n484), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n486), .A2(new_n487), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n489), .B1(new_n511), .B2(new_n461), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT30), .B1(new_n512), .B2(new_n480), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT84), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT87), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT84), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n483), .A2(new_n516), .A3(new_n484), .A4(new_n490), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n414), .A2(new_n421), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(new_n432), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT39), .B1(new_n431), .B2(new_n432), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT85), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(new_n519), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n520), .A2(new_n521), .ZN(new_n524));
  OAI221_X1 g323(.A(new_n440), .B1(KEYINPUT39), .B2(new_n519), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT40), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n525), .A2(new_n526), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n450), .A2(KEYINPUT86), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT86), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n440), .B1(new_n436), .B2(new_n530), .ZN(new_n531));
  AOI211_X1 g330(.A(new_n527), .B(new_n528), .C1(new_n529), .C2(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n514), .A2(new_n515), .A3(new_n517), .A4(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n504), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n440), .B(new_n424), .C1(new_n434), .C2(new_n435), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n443), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n536), .B1(new_n531), .B2(new_n529), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT88), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n444), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n460), .B1(new_n469), .B2(new_n472), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT37), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n541), .B1(new_n476), .B2(new_n461), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT38), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(KEYINPUT89), .B(KEYINPUT37), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n473), .A2(new_n477), .A3(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n543), .A2(new_n485), .A3(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n441), .B1(new_n450), .B2(KEYINPUT86), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n436), .A2(new_n530), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n451), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT88), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n539), .A2(new_n546), .A3(new_n481), .A4(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT38), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n480), .B1(new_n512), .B2(new_n544), .ZN(new_n553));
  OAI21_X1  g352(.A(KEYINPUT37), .B1(new_n488), .B2(new_n489), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n534), .B1(new_n551), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n514), .A2(new_n517), .A3(new_n532), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n556), .B1(KEYINPUT87), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n509), .B1(new_n533), .B2(new_n558), .ZN(new_n559));
  OAI22_X1  g358(.A1(new_n549), .A2(KEYINPUT88), .B1(new_n443), .B2(new_n442), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n537), .A2(new_n538), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT90), .B(KEYINPUT35), .ZN(new_n563));
  NOR3_X1   g362(.A1(new_n562), .A2(new_n504), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT78), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n506), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n388), .A2(KEYINPUT78), .A3(new_n390), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n514), .A2(new_n517), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n564), .A2(new_n568), .A3(new_n386), .A4(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n506), .A2(new_n386), .A3(new_n534), .ZN(new_n571));
  OAI21_X1  g370(.A(KEYINPUT35), .B1(new_n571), .B2(new_n491), .ZN(new_n572));
  AND2_X1   g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT91), .B1(new_n559), .B2(new_n573), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n393), .A2(new_n505), .A3(new_n508), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n557), .A2(KEYINPUT87), .ZN(new_n576));
  OR2_X1    g375(.A1(new_n551), .A2(new_n555), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n576), .A2(new_n534), .A3(new_n577), .A4(new_n533), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT91), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n570), .A2(new_n572), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n265), .B1(new_n574), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G99gat), .A2(G106gat), .ZN(new_n584));
  INV_X1    g383(.A(G85gat), .ZN(new_n585));
  INV_X1    g384(.A(G92gat), .ZN(new_n586));
  AOI22_X1  g385(.A1(KEYINPUT8), .A2(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT104), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G85gat), .A2(G92gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT7), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(G99gat), .B(G106gat), .Z(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(KEYINPUT105), .ZN(new_n595));
  OR2_X1    g394(.A1(new_n592), .A2(new_n593), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n595), .B(new_n596), .Z(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n598), .B1(new_n242), .B2(new_n243), .ZN(new_n599));
  XNOR2_X1  g398(.A(G190gat), .B(G218gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT106), .ZN(new_n601));
  NAND3_X1  g400(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n603), .B1(new_n597), .B2(new_n236), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n600), .A2(KEYINPUT106), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT103), .ZN(new_n609));
  XNOR2_X1  g408(.A(G134gat), .B(G162gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n607), .B(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(KEYINPUT100), .B(G57gat), .Z(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(G64gat), .ZN(new_n616));
  INV_X1    g415(.A(G57gat), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n616), .B1(new_n617), .B2(G64gat), .ZN(new_n618));
  AND2_X1   g417(.A1(G71gat), .A2(G78gat), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n619), .A2(KEYINPUT9), .ZN(new_n620));
  NOR2_X1   g419(.A1(G71gat), .A2(G78gat), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n620), .B1(new_n623), .B2(KEYINPUT101), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n618), .B(new_n624), .C1(KEYINPUT101), .C2(new_n623), .ZN(new_n625));
  XNOR2_X1  g424(.A(G57gat), .B(G64gat), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT9), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n622), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT21), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(G231gat), .A2(G233gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(G127gat), .B(G155gat), .Z(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT20), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n633), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G183gat), .B(G211gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n241), .B1(new_n629), .B2(new_n630), .ZN(new_n639));
  XOR2_X1   g438(.A(KEYINPUT102), .B(KEYINPUT19), .Z(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n638), .A2(new_n642), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n614), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(G230gat), .ZN(new_n648));
  INV_X1    g447(.A(G233gat), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n629), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n651), .A2(new_n596), .A3(new_n594), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n652), .B1(new_n597), .B2(new_n651), .ZN(new_n653));
  OR2_X1    g452(.A1(new_n653), .A2(KEYINPUT10), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n597), .A2(KEYINPUT10), .A3(new_n651), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n650), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(G120gat), .B(G148gat), .Z(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT108), .ZN(new_n659));
  XNOR2_X1  g458(.A(G176gat), .B(G204gat), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n659), .B(new_n660), .Z(new_n661));
  AND2_X1   g460(.A1(new_n653), .A2(new_n650), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n661), .B1(new_n662), .B2(KEYINPUT107), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n657), .B(new_n663), .C1(KEYINPUT107), .C2(new_n662), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n661), .B(KEYINPUT109), .Z(new_n665));
  OAI21_X1  g464(.A(new_n665), .B1(new_n656), .B2(new_n662), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n647), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n583), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n669), .A2(new_n453), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(new_n203), .ZN(G1324gat));
  INV_X1    g470(.A(new_n569), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n583), .A2(new_n672), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n673), .A2(new_n647), .A3(new_n667), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT16), .B(G8gat), .Z(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n676), .B1(new_n211), .B2(new_n674), .ZN(new_n677));
  MUX2_X1   g476(.A(new_n676), .B(new_n677), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g477(.A(G15gat), .ZN(new_n679));
  AOI22_X1  g478(.A1(new_n566), .A2(new_n567), .B1(new_n373), .B2(new_n385), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n679), .B1(new_n669), .B2(new_n681), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n682), .B(KEYINPUT110), .Z(new_n683));
  AND2_X1   g482(.A1(new_n393), .A2(new_n508), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n669), .A2(new_n679), .A3(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n683), .A2(new_n685), .ZN(G1326gat));
  NOR2_X1   g485(.A1(new_n669), .A2(new_n534), .ZN(new_n687));
  XOR2_X1   g486(.A(KEYINPUT43), .B(G22gat), .Z(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1327gat));
  NOR2_X1   g488(.A1(new_n646), .A2(new_n667), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n264), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT112), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n614), .B1(new_n574), .B2(new_n582), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  AOI221_X4 g494(.A(KEYINPUT91), .B1(new_n570), .B2(new_n572), .C1(new_n575), .C2(new_n578), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n580), .B1(new_n579), .B2(new_n581), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n613), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n698), .A2(KEYINPUT112), .A3(KEYINPUT44), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n579), .A2(new_n581), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n613), .B(KEYINPUT113), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(new_n694), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n691), .B1(new_n700), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(G29gat), .B1(new_n705), .B2(new_n453), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n613), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n583), .A2(new_n219), .A3(new_n452), .A4(new_n708), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT111), .B(KEYINPUT45), .Z(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n706), .A2(new_n711), .ZN(G1328gat));
  OAI21_X1  g511(.A(G36gat), .B1(new_n705), .B2(new_n569), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n673), .A2(G36gat), .A3(new_n707), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT46), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(G1329gat));
  INV_X1    g515(.A(G43gat), .ZN(new_n717));
  INV_X1    g516(.A(new_n684), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n717), .B1(new_n704), .B2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT47), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n583), .A2(new_n717), .A3(new_n680), .A4(new_n708), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  OR3_X1    g521(.A1(new_n719), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n720), .B1(new_n719), .B2(new_n722), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(G1330gat));
  INV_X1    g524(.A(G50gat), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n726), .B1(new_n704), .B2(new_n504), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT48), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n504), .A2(new_n726), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT114), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n583), .A2(new_n708), .A3(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  OR3_X1    g531(.A1(new_n727), .A2(new_n728), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n728), .B1(new_n727), .B2(new_n732), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(G1331gat));
  AOI211_X1 g534(.A(new_n264), .B(new_n647), .C1(new_n579), .C2(new_n581), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n736), .A2(new_n667), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n452), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n738), .B(new_n615), .Z(G1332gat));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n672), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n740), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n741));
  XOR2_X1   g540(.A(KEYINPUT49), .B(G64gat), .Z(new_n742));
  OAI21_X1  g541(.A(new_n741), .B1(new_n740), .B2(new_n742), .ZN(G1333gat));
  INV_X1    g542(.A(G71gat), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n680), .A2(new_n667), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n736), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n737), .A2(new_n718), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n748), .B2(new_n744), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g549(.A1(new_n737), .A2(new_n504), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g551(.A1(new_n265), .A2(new_n645), .A3(new_n667), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n753), .B1(new_n700), .B2(new_n703), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(G85gat), .B1(new_n755), .B2(new_n453), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n701), .A2(new_n265), .A3(new_n645), .A4(new_n613), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n757), .B(KEYINPUT51), .Z(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n667), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n452), .A2(new_n585), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n756), .B1(new_n759), .B2(new_n760), .ZN(G1336gat));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n762));
  OR2_X1    g561(.A1(new_n762), .A2(KEYINPUT52), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(KEYINPUT52), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n586), .B1(new_n754), .B2(new_n672), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n672), .A2(new_n586), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n759), .A2(new_n766), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n763), .B(new_n764), .C1(new_n765), .C2(new_n767), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n693), .A2(new_n692), .A3(new_n694), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT112), .B1(new_n698), .B2(KEYINPUT44), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n703), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n753), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n771), .A2(new_n672), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(G92gat), .ZN(new_n774));
  OR2_X1    g573(.A1(new_n759), .A2(new_n766), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n774), .A2(new_n762), .A3(new_n775), .A4(KEYINPUT52), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n768), .A2(new_n776), .ZN(G1337gat));
  OAI21_X1  g576(.A(G99gat), .B1(new_n755), .B2(new_n684), .ZN(new_n778));
  INV_X1    g577(.A(G99gat), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n758), .A2(new_n779), .A3(new_n746), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(G1338gat));
  NAND3_X1  g580(.A1(new_n754), .A2(G106gat), .A3(new_n504), .ZN(new_n782));
  INV_X1    g581(.A(G106gat), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n783), .B1(new_n759), .B2(new_n534), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g584(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n782), .A2(new_n784), .A3(new_n786), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(G1339gat));
  INV_X1    g589(.A(KEYINPUT118), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n654), .A2(new_n650), .A3(new_n655), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n657), .A2(KEYINPUT54), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n661), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT54), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n794), .B1(new_n656), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n793), .A2(KEYINPUT55), .A3(new_n796), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n797), .A2(new_n664), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n654), .A2(new_n650), .A3(new_n655), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n800), .A2(new_n656), .A3(new_n795), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n654), .A2(new_n655), .ZN(new_n802));
  INV_X1    g601(.A(new_n650), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n802), .A2(new_n795), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n661), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n799), .B1(new_n801), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n798), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n264), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n240), .B1(new_n237), .B2(new_n245), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n250), .A2(new_n251), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n812), .B1(new_n809), .B2(new_n810), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n258), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n248), .A2(new_n249), .A3(new_n252), .A4(new_n260), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n667), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n702), .B1(new_n808), .B2(new_n817), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n702), .A2(new_n807), .A3(new_n816), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n645), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n668), .A2(new_n265), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n791), .B1(new_n822), .B2(new_n534), .ZN(new_n823));
  AOI211_X1 g622(.A(KEYINPUT118), .B(new_n504), .C1(new_n820), .C2(new_n821), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n672), .A2(new_n453), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n680), .ZN(new_n828));
  OAI21_X1  g627(.A(G113gat), .B1(new_n828), .B2(new_n265), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n571), .B1(new_n820), .B2(new_n821), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n826), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n264), .A2(new_n271), .ZN(new_n832));
  XOR2_X1   g631(.A(new_n832), .B(KEYINPUT119), .Z(new_n833));
  OAI21_X1  g632(.A(new_n829), .B1(new_n831), .B2(new_n833), .ZN(G1340gat));
  INV_X1    g633(.A(new_n831), .ZN(new_n835));
  AOI21_X1  g634(.A(G120gat), .B1(new_n835), .B2(new_n667), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n745), .A2(new_n269), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n836), .B1(new_n827), .B2(new_n837), .ZN(G1341gat));
  OAI21_X1  g637(.A(G127gat), .B1(new_n828), .B2(new_n645), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n835), .A2(new_n277), .A3(new_n646), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(G1342gat));
  OAI21_X1  g640(.A(G134gat), .B1(new_n828), .B2(new_n614), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n831), .A2(G134gat), .A3(new_n614), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(KEYINPUT56), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n844), .ZN(G1343gat));
  AND2_X1   g644(.A1(new_n684), .A2(new_n826), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n534), .B1(new_n820), .B2(new_n821), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n847), .A2(KEYINPUT57), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT120), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n806), .A2(new_n850), .ZN(new_n851));
  OAI211_X1 g650(.A(KEYINPUT120), .B(new_n799), .C1(new_n801), .C2(new_n805), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n263), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n853), .A2(new_n854), .A3(new_n261), .A4(new_n798), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n613), .B1(new_n855), .B2(new_n817), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n645), .B1(new_n856), .B2(new_n819), .ZN(new_n857));
  AOI211_X1 g656(.A(new_n849), .B(new_n534), .C1(new_n857), .C2(new_n821), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n846), .B1(new_n848), .B2(new_n858), .ZN(new_n859));
  OR3_X1    g658(.A1(new_n859), .A2(new_n396), .A3(new_n265), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n847), .A2(new_n846), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n396), .B1(new_n861), .B2(new_n265), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT58), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n860), .A2(KEYINPUT58), .A3(new_n862), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(G1344gat));
  AND2_X1   g666(.A1(new_n846), .A2(new_n667), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n847), .A2(new_n397), .A3(new_n868), .ZN(new_n869));
  XOR2_X1   g668(.A(new_n869), .B(KEYINPUT121), .Z(new_n870));
  NOR2_X1   g669(.A1(new_n397), .A2(KEYINPUT59), .ZN(new_n871));
  INV_X1    g670(.A(new_n667), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n871), .B1(new_n859), .B2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n873), .B(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT124), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n613), .A2(new_n806), .A3(new_n797), .A4(new_n664), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(KEYINPUT123), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n798), .A2(new_n880), .A3(new_n613), .A4(new_n806), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n879), .A2(new_n881), .A3(new_n816), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n877), .B1(new_n856), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n879), .A2(new_n881), .A3(new_n816), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n797), .A2(new_n664), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n885), .B1(new_n851), .B2(new_n852), .ZN(new_n886));
  AOI22_X1  g685(.A1(new_n264), .A2(new_n886), .B1(new_n816), .B2(new_n667), .ZN(new_n887));
  OAI211_X1 g686(.A(KEYINPUT124), .B(new_n884), .C1(new_n887), .C2(new_n613), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n883), .A2(new_n888), .A3(new_n645), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n534), .B1(new_n889), .B2(new_n821), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT125), .B1(new_n890), .B2(KEYINPUT57), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT125), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n884), .B1(new_n887), .B2(new_n613), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n646), .B1(new_n893), .B2(new_n877), .ZN(new_n894));
  AOI22_X1  g693(.A1(new_n894), .A2(new_n888), .B1(new_n265), .B2(new_n668), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n892), .B(new_n849), .C1(new_n895), .C2(new_n534), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n822), .A2(KEYINPUT57), .A3(new_n504), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n891), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n868), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n876), .B1(new_n899), .B2(G148gat), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n870), .B1(new_n875), .B2(new_n900), .ZN(G1345gat));
  OAI21_X1  g700(.A(G155gat), .B1(new_n859), .B2(new_n645), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n645), .A2(G155gat), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n902), .B1(new_n861), .B2(new_n903), .ZN(G1346gat));
  NAND2_X1  g703(.A1(new_n702), .A2(G162gat), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n859), .A2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(G162gat), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n907), .B1(new_n861), .B2(new_n614), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n906), .A2(new_n908), .ZN(G1347gat));
  NOR2_X1   g708(.A1(new_n569), .A2(new_n452), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n830), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT126), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n912), .A2(new_n264), .A3(new_n313), .A4(new_n315), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n680), .B(new_n910), .C1(new_n823), .C2(new_n824), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n914), .A2(new_n265), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT127), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n915), .A2(new_n916), .A3(G169gat), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n916), .B1(new_n915), .B2(G169gat), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n913), .B1(new_n918), .B2(new_n919), .ZN(G1348gat));
  AOI21_X1  g719(.A(G176gat), .B1(new_n912), .B2(new_n667), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n825), .A2(new_n910), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n745), .B1(new_n310), .B2(new_n311), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(G1349gat));
  OAI21_X1  g723(.A(G183gat), .B1(new_n914), .B2(new_n645), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n830), .A2(new_n351), .A3(new_n646), .A4(new_n910), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g727(.A1(new_n912), .A2(new_n300), .A3(new_n702), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n914), .A2(new_n614), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT61), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n930), .A2(new_n931), .A3(G190gat), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n931), .B1(new_n930), .B2(G190gat), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n929), .B1(new_n933), .B2(new_n934), .ZN(G1351gat));
  NAND2_X1  g734(.A1(new_n684), .A2(new_n910), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n847), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(G197gat), .B1(new_n938), .B2(new_n264), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n898), .A2(new_n937), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n264), .A2(G197gat), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(G1352gat));
  OAI21_X1  g742(.A(G204gat), .B1(new_n940), .B2(new_n872), .ZN(new_n944));
  INV_X1    g743(.A(G204gat), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n938), .A2(new_n945), .A3(new_n667), .ZN(new_n946));
  XOR2_X1   g745(.A(new_n946), .B(KEYINPUT62), .Z(new_n947));
  NAND2_X1  g746(.A1(new_n944), .A2(new_n947), .ZN(G1353gat));
  NAND3_X1  g747(.A1(new_n938), .A2(new_n455), .A3(new_n646), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n898), .A2(new_n646), .A3(new_n937), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n950), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n951));
  AOI21_X1  g750(.A(KEYINPUT63), .B1(new_n950), .B2(G211gat), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(G1354gat));
  OAI21_X1  g752(.A(G218gat), .B1(new_n940), .B2(new_n614), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n938), .A2(new_n456), .A3(new_n702), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1355gat));
endmodule


