

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U552 ( .A1(G8), .A2(n703), .ZN(n749) );
  OR2_X1 U553 ( .A1(n731), .A2(n730), .ZN(n732) );
  OR2_X1 U554 ( .A1(n752), .A2(n729), .ZN(n730) );
  NOR2_X1 U555 ( .A1(n584), .A2(n537), .ZN(n801) );
  NOR2_X1 U556 ( .A1(n684), .A2(n683), .ZN(n685) );
  INV_X1 U557 ( .A(KEYINPUT29), .ZN(n696) );
  XNOR2_X1 U558 ( .A(n697), .B(n696), .ZN(n700) );
  NOR2_X1 U559 ( .A1(n749), .A2(G1966), .ZN(n717) );
  INV_X1 U560 ( .A(KEYINPUT64), .ZN(n738) );
  XNOR2_X1 U561 ( .A(KEYINPUT13), .B(KEYINPUT72), .ZN(n674) );
  XNOR2_X1 U562 ( .A(n675), .B(n674), .ZN(n676) );
  NOR2_X1 U563 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  NOR2_X1 U564 ( .A1(G2105), .A2(n523), .ZN(n890) );
  AND2_X1 U565 ( .A1(n733), .A2(n732), .ZN(n759) );
  NOR2_X1 U566 ( .A1(G651), .A2(n584), .ZN(n798) );
  NOR2_X2 U567 ( .A1(n528), .A2(n527), .ZN(G160) );
  INV_X1 U568 ( .A(G2105), .ZN(n522) );
  NOR2_X1 U569 ( .A1(G2104), .A2(n522), .ZN(n886) );
  NAND2_X1 U570 ( .A1(G125), .A2(n886), .ZN(n518) );
  XNOR2_X1 U571 ( .A(n518), .B(KEYINPUT66), .ZN(n521) );
  INV_X1 U572 ( .A(G2104), .ZN(n523) );
  NAND2_X1 U573 ( .A1(G101), .A2(n890), .ZN(n519) );
  XOR2_X1 U574 ( .A(KEYINPUT23), .B(n519), .Z(n520) );
  NAND2_X1 U575 ( .A1(n521), .A2(n520), .ZN(n528) );
  NOR2_X4 U576 ( .A1(n523), .A2(n522), .ZN(n885) );
  NAND2_X1 U577 ( .A1(G113), .A2(n885), .ZN(n526) );
  XOR2_X2 U578 ( .A(KEYINPUT17), .B(n524), .Z(n893) );
  NAND2_X1 U579 ( .A1(G137), .A2(n893), .ZN(n525) );
  NAND2_X1 U580 ( .A1(n526), .A2(n525), .ZN(n527) );
  NAND2_X1 U581 ( .A1(G138), .A2(n893), .ZN(n530) );
  NAND2_X1 U582 ( .A1(G126), .A2(n886), .ZN(n529) );
  AND2_X1 U583 ( .A1(n530), .A2(n529), .ZN(n535) );
  NAND2_X1 U584 ( .A1(G114), .A2(n885), .ZN(n531) );
  XNOR2_X1 U585 ( .A(KEYINPUT91), .B(n531), .ZN(n533) );
  AND2_X1 U586 ( .A1(n890), .A2(G102), .ZN(n532) );
  NOR2_X1 U587 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U588 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U589 ( .A(KEYINPUT92), .B(n536), .Z(G164) );
  XOR2_X1 U590 ( .A(KEYINPUT0), .B(G543), .Z(n584) );
  INV_X1 U591 ( .A(G651), .ZN(n537) );
  NAND2_X1 U592 ( .A1(G72), .A2(n801), .ZN(n541) );
  NOR2_X1 U593 ( .A1(G543), .A2(n537), .ZN(n539) );
  XNOR2_X1 U594 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n538) );
  XNOR2_X1 U595 ( .A(n539), .B(n538), .ZN(n797) );
  NAND2_X1 U596 ( .A1(G60), .A2(n797), .ZN(n540) );
  NAND2_X1 U597 ( .A1(n541), .A2(n540), .ZN(n545) );
  NOR2_X1 U598 ( .A1(G651), .A2(G543), .ZN(n802) );
  NAND2_X1 U599 ( .A1(G85), .A2(n802), .ZN(n543) );
  NAND2_X1 U600 ( .A1(G47), .A2(n798), .ZN(n542) );
  NAND2_X1 U601 ( .A1(n543), .A2(n542), .ZN(n544) );
  OR2_X1 U602 ( .A1(n545), .A2(n544), .ZN(G290) );
  NAND2_X1 U603 ( .A1(G89), .A2(n802), .ZN(n546) );
  XOR2_X1 U604 ( .A(KEYINPUT4), .B(n546), .Z(n547) );
  XNOR2_X1 U605 ( .A(n547), .B(KEYINPUT77), .ZN(n549) );
  NAND2_X1 U606 ( .A1(G76), .A2(n801), .ZN(n548) );
  NAND2_X1 U607 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U608 ( .A(n550), .B(KEYINPUT5), .ZN(n555) );
  NAND2_X1 U609 ( .A1(G63), .A2(n797), .ZN(n552) );
  NAND2_X1 U610 ( .A1(G51), .A2(n798), .ZN(n551) );
  NAND2_X1 U611 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U612 ( .A(KEYINPUT6), .B(n553), .Z(n554) );
  NAND2_X1 U613 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U614 ( .A(n556), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U615 ( .A1(n798), .A2(G52), .ZN(n558) );
  NAND2_X1 U616 ( .A1(n797), .A2(G64), .ZN(n557) );
  NAND2_X1 U617 ( .A1(n558), .A2(n557), .ZN(n563) );
  NAND2_X1 U618 ( .A1(G77), .A2(n801), .ZN(n560) );
  NAND2_X1 U619 ( .A1(G90), .A2(n802), .ZN(n559) );
  NAND2_X1 U620 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U621 ( .A(KEYINPUT9), .B(n561), .Z(n562) );
  NOR2_X1 U622 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U623 ( .A(KEYINPUT68), .B(n564), .ZN(G171) );
  XOR2_X1 U624 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U625 ( .A1(G88), .A2(n802), .ZN(n565) );
  XOR2_X1 U626 ( .A(KEYINPUT86), .B(n565), .Z(n570) );
  NAND2_X1 U627 ( .A1(G62), .A2(n797), .ZN(n567) );
  NAND2_X1 U628 ( .A1(G50), .A2(n798), .ZN(n566) );
  NAND2_X1 U629 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U630 ( .A(KEYINPUT85), .B(n568), .Z(n569) );
  NOR2_X1 U631 ( .A1(n570), .A2(n569), .ZN(n572) );
  NAND2_X1 U632 ( .A1(n801), .A2(G75), .ZN(n571) );
  NAND2_X1 U633 ( .A1(n572), .A2(n571), .ZN(G303) );
  INV_X1 U634 ( .A(G303), .ZN(G166) );
  NAND2_X1 U635 ( .A1(n797), .A2(G61), .ZN(n573) );
  XNOR2_X1 U636 ( .A(KEYINPUT81), .B(n573), .ZN(n580) );
  XOR2_X1 U637 ( .A(KEYINPUT83), .B(KEYINPUT2), .Z(n575) );
  NAND2_X1 U638 ( .A1(G73), .A2(n801), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U640 ( .A(n576), .B(KEYINPUT82), .ZN(n578) );
  NAND2_X1 U641 ( .A1(n802), .A2(G86), .ZN(n577) );
  NAND2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U643 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U644 ( .A(n581), .B(KEYINPUT84), .ZN(n583) );
  NAND2_X1 U645 ( .A1(G48), .A2(n798), .ZN(n582) );
  NAND2_X1 U646 ( .A1(n583), .A2(n582), .ZN(G305) );
  NAND2_X1 U647 ( .A1(G87), .A2(n584), .ZN(n585) );
  XNOR2_X1 U648 ( .A(n585), .B(KEYINPUT80), .ZN(n590) );
  NAND2_X1 U649 ( .A1(G49), .A2(n798), .ZN(n587) );
  NAND2_X1 U650 ( .A1(G74), .A2(G651), .ZN(n586) );
  NAND2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U652 ( .A1(n797), .A2(n588), .ZN(n589) );
  NAND2_X1 U653 ( .A1(n590), .A2(n589), .ZN(G288) );
  NOR2_X1 U654 ( .A1(G1384), .A2(G164), .ZN(n635) );
  NAND2_X1 U655 ( .A1(G160), .A2(G40), .ZN(n629) );
  NOR2_X1 U656 ( .A1(n635), .A2(n629), .ZN(n627) );
  XNOR2_X1 U657 ( .A(G2067), .B(KEYINPUT37), .ZN(n591) );
  XNOR2_X1 U658 ( .A(n591), .B(KEYINPUT93), .ZN(n601) );
  NAND2_X1 U659 ( .A1(G116), .A2(n885), .ZN(n593) );
  NAND2_X1 U660 ( .A1(G128), .A2(n886), .ZN(n592) );
  NAND2_X1 U661 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U662 ( .A(n594), .B(KEYINPUT35), .ZN(n599) );
  NAND2_X1 U663 ( .A1(G140), .A2(n893), .ZN(n596) );
  NAND2_X1 U664 ( .A1(G104), .A2(n890), .ZN(n595) );
  NAND2_X1 U665 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U666 ( .A(KEYINPUT34), .B(n597), .Z(n598) );
  NAND2_X1 U667 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U668 ( .A(n600), .B(KEYINPUT36), .ZN(n905) );
  NAND2_X1 U669 ( .A1(n601), .A2(n905), .ZN(n997) );
  NAND2_X1 U670 ( .A1(n627), .A2(n997), .ZN(n625) );
  NOR2_X1 U671 ( .A1(n601), .A2(n905), .ZN(n1005) );
  NAND2_X1 U672 ( .A1(G141), .A2(n893), .ZN(n603) );
  NAND2_X1 U673 ( .A1(G129), .A2(n886), .ZN(n602) );
  NAND2_X1 U674 ( .A1(n603), .A2(n602), .ZN(n606) );
  NAND2_X1 U675 ( .A1(n890), .A2(G105), .ZN(n604) );
  XOR2_X1 U676 ( .A(KEYINPUT38), .B(n604), .Z(n605) );
  NOR2_X1 U677 ( .A1(n606), .A2(n605), .ZN(n608) );
  NAND2_X1 U678 ( .A1(n885), .A2(G117), .ZN(n607) );
  NAND2_X1 U679 ( .A1(n608), .A2(n607), .ZN(n897) );
  NOR2_X1 U680 ( .A1(G1996), .A2(n897), .ZN(n1009) );
  NOR2_X1 U681 ( .A1(G1986), .A2(G290), .ZN(n615) );
  NAND2_X1 U682 ( .A1(G107), .A2(n885), .ZN(n610) );
  NAND2_X1 U683 ( .A1(G119), .A2(n886), .ZN(n609) );
  NAND2_X1 U684 ( .A1(n610), .A2(n609), .ZN(n614) );
  NAND2_X1 U685 ( .A1(G131), .A2(n893), .ZN(n612) );
  NAND2_X1 U686 ( .A1(G95), .A2(n890), .ZN(n611) );
  NAND2_X1 U687 ( .A1(n612), .A2(n611), .ZN(n613) );
  OR2_X1 U688 ( .A1(n614), .A2(n613), .ZN(n882) );
  NOR2_X1 U689 ( .A1(G1991), .A2(n882), .ZN(n995) );
  NOR2_X1 U690 ( .A1(n615), .A2(n995), .ZN(n619) );
  NAND2_X1 U691 ( .A1(G1991), .A2(n882), .ZN(n617) );
  NAND2_X1 U692 ( .A1(G1996), .A2(n897), .ZN(n616) );
  NAND2_X1 U693 ( .A1(n617), .A2(n616), .ZN(n1004) );
  NAND2_X1 U694 ( .A1(n627), .A2(n1004), .ZN(n618) );
  XOR2_X1 U695 ( .A(KEYINPUT94), .B(n618), .Z(n752) );
  NOR2_X1 U696 ( .A1(n619), .A2(n752), .ZN(n620) );
  NOR2_X1 U697 ( .A1(n1009), .A2(n620), .ZN(n621) );
  XNOR2_X1 U698 ( .A(n621), .B(KEYINPUT39), .ZN(n622) );
  XNOR2_X1 U699 ( .A(n622), .B(KEYINPUT104), .ZN(n623) );
  NOR2_X1 U700 ( .A1(n1005), .A2(n623), .ZN(n624) );
  NOR2_X1 U701 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U702 ( .A(KEYINPUT105), .B(n626), .ZN(n733) );
  XOR2_X1 U703 ( .A(G1986), .B(G290), .Z(n934) );
  NAND2_X1 U704 ( .A1(n997), .A2(n934), .ZN(n628) );
  NAND2_X1 U705 ( .A1(n628), .A2(n627), .ZN(n754) );
  INV_X1 U706 ( .A(n754), .ZN(n731) );
  INV_X1 U707 ( .A(n629), .ZN(n634) );
  NAND2_X2 U708 ( .A1(n635), .A2(n634), .ZN(n703) );
  NOR2_X1 U709 ( .A1(G2084), .A2(n703), .ZN(n714) );
  NOR2_X1 U710 ( .A1(n717), .A2(n714), .ZN(n630) );
  NAND2_X1 U711 ( .A1(n630), .A2(G8), .ZN(n631) );
  XNOR2_X1 U712 ( .A(n631), .B(KEYINPUT30), .ZN(n632) );
  NOR2_X1 U713 ( .A1(n632), .A2(G168), .ZN(n633) );
  XNOR2_X1 U714 ( .A(n633), .B(KEYINPUT99), .ZN(n640) );
  XOR2_X1 U715 ( .A(G2078), .B(KEYINPUT25), .Z(n975) );
  NOR2_X1 U716 ( .A1(n975), .A2(n703), .ZN(n637) );
  AND2_X1 U717 ( .A1(n635), .A2(n634), .ZN(n666) );
  NOR2_X1 U718 ( .A1(n666), .A2(G1961), .ZN(n636) );
  NOR2_X1 U719 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U720 ( .A(KEYINPUT95), .B(n638), .ZN(n698) );
  OR2_X1 U721 ( .A1(n698), .A2(G171), .ZN(n639) );
  NAND2_X1 U722 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U723 ( .A(n641), .B(KEYINPUT31), .ZN(n702) );
  NAND2_X1 U724 ( .A1(G65), .A2(n797), .ZN(n643) );
  NAND2_X1 U725 ( .A1(G53), .A2(n798), .ZN(n642) );
  NAND2_X1 U726 ( .A1(n643), .A2(n642), .ZN(n647) );
  NAND2_X1 U727 ( .A1(G78), .A2(n801), .ZN(n645) );
  NAND2_X1 U728 ( .A1(G91), .A2(n802), .ZN(n644) );
  NAND2_X1 U729 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U730 ( .A1(n647), .A2(n646), .ZN(n927) );
  NAND2_X1 U731 ( .A1(G1956), .A2(n703), .ZN(n648) );
  XNOR2_X1 U732 ( .A(KEYINPUT97), .B(n648), .ZN(n652) );
  NAND2_X1 U733 ( .A1(n666), .A2(G2072), .ZN(n650) );
  XOR2_X1 U734 ( .A(KEYINPUT96), .B(KEYINPUT27), .Z(n649) );
  XOR2_X1 U735 ( .A(n650), .B(n649), .Z(n651) );
  NOR2_X1 U736 ( .A1(n652), .A2(n651), .ZN(n691) );
  NOR2_X1 U737 ( .A1(n927), .A2(n691), .ZN(n654) );
  XOR2_X1 U738 ( .A(KEYINPUT28), .B(KEYINPUT98), .Z(n653) );
  XNOR2_X1 U739 ( .A(n654), .B(n653), .ZN(n695) );
  NAND2_X1 U740 ( .A1(G79), .A2(n801), .ZN(n656) );
  NAND2_X1 U741 ( .A1(G54), .A2(n798), .ZN(n655) );
  NAND2_X1 U742 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U743 ( .A(KEYINPUT74), .B(n657), .ZN(n661) );
  NAND2_X1 U744 ( .A1(G92), .A2(n802), .ZN(n659) );
  NAND2_X1 U745 ( .A1(G66), .A2(n797), .ZN(n658) );
  NAND2_X1 U746 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U747 ( .A1(n661), .A2(n660), .ZN(n663) );
  XNOR2_X1 U748 ( .A(KEYINPUT75), .B(KEYINPUT15), .ZN(n662) );
  XNOR2_X1 U749 ( .A(n663), .B(n662), .ZN(n919) );
  AND2_X1 U750 ( .A1(n666), .A2(G2067), .ZN(n665) );
  INV_X1 U751 ( .A(G1348), .ZN(n951) );
  NOR2_X1 U752 ( .A1(n666), .A2(n951), .ZN(n664) );
  NOR2_X1 U753 ( .A1(n665), .A2(n664), .ZN(n688) );
  NAND2_X1 U754 ( .A1(n919), .A2(n688), .ZN(n687) );
  NAND2_X1 U755 ( .A1(n666), .A2(G1996), .ZN(n668) );
  INV_X1 U756 ( .A(KEYINPUT26), .ZN(n667) );
  XNOR2_X1 U757 ( .A(n668), .B(n667), .ZN(n684) );
  NAND2_X1 U758 ( .A1(n703), .A2(G1341), .ZN(n682) );
  NAND2_X1 U759 ( .A1(n797), .A2(G56), .ZN(n669) );
  XNOR2_X1 U760 ( .A(n669), .B(KEYINPUT14), .ZN(n677) );
  NAND2_X1 U761 ( .A1(G68), .A2(n801), .ZN(n673) );
  XOR2_X1 U762 ( .A(KEYINPUT71), .B(KEYINPUT12), .Z(n671) );
  NAND2_X1 U763 ( .A1(G81), .A2(n802), .ZN(n670) );
  XNOR2_X1 U764 ( .A(n671), .B(n670), .ZN(n672) );
  NAND2_X1 U765 ( .A1(n673), .A2(n672), .ZN(n675) );
  NAND2_X1 U766 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U767 ( .A(n678), .B(KEYINPUT73), .ZN(n680) );
  NAND2_X1 U768 ( .A1(G43), .A2(n798), .ZN(n679) );
  NAND2_X1 U769 ( .A1(n680), .A2(n679), .ZN(n922) );
  INV_X1 U770 ( .A(n922), .ZN(n681) );
  NAND2_X1 U771 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U772 ( .A(KEYINPUT65), .B(n685), .ZN(n686) );
  NAND2_X1 U773 ( .A1(n687), .A2(n686), .ZN(n690) );
  OR2_X1 U774 ( .A1(n919), .A2(n688), .ZN(n689) );
  NAND2_X1 U775 ( .A1(n690), .A2(n689), .ZN(n693) );
  NAND2_X1 U776 ( .A1(n927), .A2(n691), .ZN(n692) );
  NAND2_X1 U777 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U778 ( .A1(n695), .A2(n694), .ZN(n697) );
  NAND2_X1 U779 ( .A1(n698), .A2(G171), .ZN(n699) );
  NAND2_X1 U780 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U781 ( .A1(n702), .A2(n701), .ZN(n715) );
  NAND2_X1 U782 ( .A1(n715), .A2(G286), .ZN(n710) );
  NOR2_X1 U783 ( .A1(G1971), .A2(n749), .ZN(n705) );
  NOR2_X1 U784 ( .A1(G2090), .A2(n703), .ZN(n704) );
  NOR2_X1 U785 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U786 ( .A(KEYINPUT100), .B(n706), .Z(n707) );
  NOR2_X1 U787 ( .A1(G166), .A2(n707), .ZN(n708) );
  XNOR2_X1 U788 ( .A(n708), .B(KEYINPUT101), .ZN(n709) );
  NAND2_X1 U789 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U790 ( .A(n711), .B(KEYINPUT102), .ZN(n712) );
  NAND2_X1 U791 ( .A1(n712), .A2(G8), .ZN(n713) );
  XNOR2_X1 U792 ( .A(n713), .B(KEYINPUT32), .ZN(n721) );
  NAND2_X1 U793 ( .A1(G8), .A2(n714), .ZN(n719) );
  INV_X1 U794 ( .A(n715), .ZN(n716) );
  NOR2_X1 U795 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U796 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U797 ( .A1(n721), .A2(n720), .ZN(n735) );
  NOR2_X1 U798 ( .A1(G2090), .A2(G303), .ZN(n722) );
  NAND2_X1 U799 ( .A1(G8), .A2(n722), .ZN(n723) );
  NAND2_X1 U800 ( .A1(n735), .A2(n723), .ZN(n724) );
  AND2_X1 U801 ( .A1(n724), .A2(n749), .ZN(n728) );
  NOR2_X1 U802 ( .A1(G1981), .A2(G305), .ZN(n725) );
  XOR2_X1 U803 ( .A(n725), .B(KEYINPUT24), .Z(n726) );
  NOR2_X1 U804 ( .A1(n749), .A2(n726), .ZN(n727) );
  NOR2_X1 U805 ( .A1(n728), .A2(n727), .ZN(n729) );
  NOR2_X1 U806 ( .A1(G1976), .A2(G288), .ZN(n745) );
  NOR2_X1 U807 ( .A1(G1971), .A2(G303), .ZN(n734) );
  NOR2_X1 U808 ( .A1(n745), .A2(n734), .ZN(n920) );
  NAND2_X1 U809 ( .A1(n735), .A2(n920), .ZN(n736) );
  NAND2_X1 U810 ( .A1(G1976), .A2(G288), .ZN(n928) );
  NAND2_X1 U811 ( .A1(n736), .A2(n928), .ZN(n737) );
  NOR2_X1 U812 ( .A1(n737), .A2(n749), .ZN(n739) );
  XNOR2_X1 U813 ( .A(n739), .B(n738), .ZN(n741) );
  INV_X1 U814 ( .A(KEYINPUT103), .ZN(n744) );
  NOR2_X1 U815 ( .A1(n749), .A2(n744), .ZN(n740) );
  NOR2_X1 U816 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U817 ( .A1(KEYINPUT33), .A2(n742), .ZN(n751) );
  NAND2_X1 U818 ( .A1(n745), .A2(KEYINPUT33), .ZN(n743) );
  NAND2_X1 U819 ( .A1(n744), .A2(n743), .ZN(n747) );
  NAND2_X1 U820 ( .A1(n745), .A2(KEYINPUT103), .ZN(n746) );
  NAND2_X1 U821 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U822 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U823 ( .A1(n751), .A2(n750), .ZN(n757) );
  XOR2_X1 U824 ( .A(G1981), .B(G305), .Z(n916) );
  INV_X1 U825 ( .A(n752), .ZN(n753) );
  AND2_X1 U826 ( .A1(n916), .A2(n753), .ZN(n755) );
  AND2_X1 U827 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U828 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U829 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U830 ( .A(n760), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U831 ( .A(G2438), .B(G2454), .Z(n762) );
  XNOR2_X1 U832 ( .A(G2435), .B(G2430), .ZN(n761) );
  XNOR2_X1 U833 ( .A(n762), .B(n761), .ZN(n763) );
  XOR2_X1 U834 ( .A(n763), .B(G2427), .Z(n765) );
  XNOR2_X1 U835 ( .A(G1348), .B(G1341), .ZN(n764) );
  XNOR2_X1 U836 ( .A(n765), .B(n764), .ZN(n769) );
  XOR2_X1 U837 ( .A(G2443), .B(G2446), .Z(n767) );
  XNOR2_X1 U838 ( .A(KEYINPUT106), .B(G2451), .ZN(n766) );
  XNOR2_X1 U839 ( .A(n767), .B(n766), .ZN(n768) );
  XOR2_X1 U840 ( .A(n769), .B(n768), .Z(n770) );
  AND2_X1 U841 ( .A1(G14), .A2(n770), .ZN(G401) );
  AND2_X1 U842 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U843 ( .A1(G111), .A2(n885), .ZN(n772) );
  NAND2_X1 U844 ( .A1(G135), .A2(n893), .ZN(n771) );
  NAND2_X1 U845 ( .A1(n772), .A2(n771), .ZN(n775) );
  NAND2_X1 U846 ( .A1(n886), .A2(G123), .ZN(n773) );
  XOR2_X1 U847 ( .A(KEYINPUT18), .B(n773), .Z(n774) );
  NOR2_X1 U848 ( .A1(n775), .A2(n774), .ZN(n777) );
  NAND2_X1 U849 ( .A1(n890), .A2(G99), .ZN(n776) );
  NAND2_X1 U850 ( .A1(n777), .A2(n776), .ZN(n992) );
  XNOR2_X1 U851 ( .A(G2096), .B(n992), .ZN(n778) );
  OR2_X1 U852 ( .A1(G2100), .A2(n778), .ZN(G156) );
  INV_X1 U853 ( .A(G82), .ZN(G220) );
  INV_X1 U854 ( .A(G57), .ZN(G237) );
  NAND2_X1 U855 ( .A1(G7), .A2(G661), .ZN(n779) );
  XNOR2_X1 U856 ( .A(n779), .B(KEYINPUT10), .ZN(n780) );
  XNOR2_X1 U857 ( .A(KEYINPUT70), .B(n780), .ZN(G223) );
  INV_X1 U858 ( .A(G223), .ZN(n835) );
  NAND2_X1 U859 ( .A1(n835), .A2(G567), .ZN(n781) );
  XOR2_X1 U860 ( .A(KEYINPUT11), .B(n781), .Z(G234) );
  INV_X1 U861 ( .A(G860), .ZN(n788) );
  OR2_X1 U862 ( .A1(n922), .A2(n788), .ZN(G153) );
  INV_X1 U863 ( .A(G171), .ZN(G301) );
  OR2_X1 U864 ( .A1(n919), .A2(G868), .ZN(n782) );
  XNOR2_X1 U865 ( .A(n782), .B(KEYINPUT76), .ZN(n784) );
  NAND2_X1 U866 ( .A1(G868), .A2(G301), .ZN(n783) );
  NAND2_X1 U867 ( .A1(n784), .A2(n783), .ZN(G284) );
  INV_X1 U868 ( .A(n927), .ZN(G299) );
  INV_X1 U869 ( .A(G868), .ZN(n785) );
  NOR2_X1 U870 ( .A1(G286), .A2(n785), .ZN(n787) );
  NOR2_X1 U871 ( .A1(G868), .A2(G299), .ZN(n786) );
  NOR2_X1 U872 ( .A1(n787), .A2(n786), .ZN(G297) );
  NAND2_X1 U873 ( .A1(G559), .A2(n788), .ZN(n789) );
  XNOR2_X1 U874 ( .A(KEYINPUT78), .B(n789), .ZN(n790) );
  NAND2_X1 U875 ( .A1(n790), .A2(n919), .ZN(n791) );
  XNOR2_X1 U876 ( .A(KEYINPUT16), .B(n791), .ZN(G148) );
  NAND2_X1 U877 ( .A1(n919), .A2(G868), .ZN(n792) );
  XOR2_X1 U878 ( .A(KEYINPUT79), .B(n792), .Z(n793) );
  NOR2_X1 U879 ( .A1(G559), .A2(n793), .ZN(n795) );
  NOR2_X1 U880 ( .A1(G868), .A2(n922), .ZN(n794) );
  NOR2_X1 U881 ( .A1(n795), .A2(n794), .ZN(G282) );
  NAND2_X1 U882 ( .A1(n919), .A2(G559), .ZN(n817) );
  XNOR2_X1 U883 ( .A(n922), .B(n817), .ZN(n796) );
  NOR2_X1 U884 ( .A1(n796), .A2(G860), .ZN(n807) );
  NAND2_X1 U885 ( .A1(G67), .A2(n797), .ZN(n800) );
  NAND2_X1 U886 ( .A1(G55), .A2(n798), .ZN(n799) );
  NAND2_X1 U887 ( .A1(n800), .A2(n799), .ZN(n806) );
  NAND2_X1 U888 ( .A1(G80), .A2(n801), .ZN(n804) );
  NAND2_X1 U889 ( .A1(G93), .A2(n802), .ZN(n803) );
  NAND2_X1 U890 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U891 ( .A1(n806), .A2(n805), .ZN(n809) );
  XNOR2_X1 U892 ( .A(n807), .B(n809), .ZN(G145) );
  NOR2_X1 U893 ( .A1(n809), .A2(G868), .ZN(n808) );
  XNOR2_X1 U894 ( .A(KEYINPUT89), .B(n808), .ZN(n821) );
  XNOR2_X1 U895 ( .A(n922), .B(G305), .ZN(n816) );
  XNOR2_X1 U896 ( .A(n809), .B(KEYINPUT19), .ZN(n810) );
  XNOR2_X1 U897 ( .A(n810), .B(KEYINPUT87), .ZN(n813) );
  XNOR2_X1 U898 ( .A(n927), .B(G303), .ZN(n811) );
  XNOR2_X1 U899 ( .A(n811), .B(G290), .ZN(n812) );
  XNOR2_X1 U900 ( .A(n813), .B(n812), .ZN(n814) );
  XNOR2_X1 U901 ( .A(n814), .B(G288), .ZN(n815) );
  XNOR2_X1 U902 ( .A(n816), .B(n815), .ZN(n841) );
  XNOR2_X1 U903 ( .A(n841), .B(n817), .ZN(n818) );
  NAND2_X1 U904 ( .A1(n818), .A2(G868), .ZN(n819) );
  XNOR2_X1 U905 ( .A(KEYINPUT88), .B(n819), .ZN(n820) );
  NAND2_X1 U906 ( .A1(n821), .A2(n820), .ZN(G295) );
  NAND2_X1 U907 ( .A1(G2078), .A2(G2084), .ZN(n822) );
  XOR2_X1 U908 ( .A(KEYINPUT20), .B(n822), .Z(n823) );
  NAND2_X1 U909 ( .A1(G2090), .A2(n823), .ZN(n824) );
  XNOR2_X1 U910 ( .A(KEYINPUT21), .B(n824), .ZN(n825) );
  NAND2_X1 U911 ( .A1(n825), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U912 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U913 ( .A(KEYINPUT69), .B(G132), .ZN(G219) );
  NAND2_X1 U914 ( .A1(G108), .A2(G120), .ZN(n826) );
  NOR2_X1 U915 ( .A1(G237), .A2(n826), .ZN(n827) );
  NAND2_X1 U916 ( .A1(G69), .A2(n827), .ZN(n839) );
  NAND2_X1 U917 ( .A1(n839), .A2(G567), .ZN(n833) );
  NOR2_X1 U918 ( .A1(G220), .A2(G219), .ZN(n828) );
  XNOR2_X1 U919 ( .A(KEYINPUT22), .B(n828), .ZN(n829) );
  NAND2_X1 U920 ( .A1(n829), .A2(G96), .ZN(n830) );
  NOR2_X1 U921 ( .A1(G218), .A2(n830), .ZN(n831) );
  XOR2_X1 U922 ( .A(KEYINPUT90), .B(n831), .Z(n840) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n840), .ZN(n832) );
  NAND2_X1 U924 ( .A1(n833), .A2(n832), .ZN(n915) );
  NAND2_X1 U925 ( .A1(G661), .A2(G483), .ZN(n834) );
  NOR2_X1 U926 ( .A1(n915), .A2(n834), .ZN(n838) );
  NAND2_X1 U927 ( .A1(n838), .A2(G36), .ZN(G176) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n835), .ZN(G217) );
  AND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n836) );
  NAND2_X1 U930 ( .A1(G661), .A2(n836), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U932 ( .A1(n838), .A2(n837), .ZN(G188) );
  XNOR2_X1 U933 ( .A(G120), .B(KEYINPUT107), .ZN(G236) );
  NOR2_X1 U934 ( .A1(n840), .A2(n839), .ZN(G325) );
  XOR2_X1 U935 ( .A(KEYINPUT108), .B(G325), .Z(G261) );
  INV_X1 U937 ( .A(G108), .ZN(G238) );
  INV_X1 U938 ( .A(G96), .ZN(G221) );
  XNOR2_X1 U939 ( .A(n841), .B(KEYINPUT116), .ZN(n843) );
  XNOR2_X1 U940 ( .A(n919), .B(G286), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(n844) );
  XNOR2_X1 U942 ( .A(G301), .B(n844), .ZN(n845) );
  NOR2_X1 U943 ( .A1(G37), .A2(n845), .ZN(G397) );
  XOR2_X1 U944 ( .A(G2100), .B(G2096), .Z(n847) );
  XNOR2_X1 U945 ( .A(KEYINPUT42), .B(G2678), .ZN(n846) );
  XNOR2_X1 U946 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U947 ( .A(KEYINPUT43), .B(G2090), .Z(n849) );
  XNOR2_X1 U948 ( .A(G2067), .B(G2072), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U950 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U951 ( .A(G2078), .B(G2084), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(G227) );
  XOR2_X1 U953 ( .A(G1986), .B(G1956), .Z(n855) );
  XNOR2_X1 U954 ( .A(G1966), .B(G1961), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U956 ( .A(G1976), .B(G1971), .Z(n857) );
  XNOR2_X1 U957 ( .A(G1991), .B(G1996), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U959 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U960 ( .A(G2474), .B(KEYINPUT41), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n861), .B(n860), .ZN(n863) );
  XOR2_X1 U962 ( .A(G1981), .B(KEYINPUT109), .Z(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(G229) );
  NAND2_X1 U964 ( .A1(n890), .A2(G100), .ZN(n870) );
  NAND2_X1 U965 ( .A1(G112), .A2(n885), .ZN(n865) );
  NAND2_X1 U966 ( .A1(G136), .A2(n893), .ZN(n864) );
  NAND2_X1 U967 ( .A1(n865), .A2(n864), .ZN(n868) );
  NAND2_X1 U968 ( .A1(n886), .A2(G124), .ZN(n866) );
  XOR2_X1 U969 ( .A(KEYINPUT44), .B(n866), .Z(n867) );
  NOR2_X1 U970 ( .A1(n868), .A2(n867), .ZN(n869) );
  NAND2_X1 U971 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U972 ( .A(KEYINPUT110), .B(n871), .Z(G162) );
  NAND2_X1 U973 ( .A1(G106), .A2(n890), .ZN(n874) );
  NAND2_X1 U974 ( .A1(n893), .A2(G142), .ZN(n872) );
  XOR2_X1 U975 ( .A(KEYINPUT111), .B(n872), .Z(n873) );
  NAND2_X1 U976 ( .A1(n874), .A2(n873), .ZN(n877) );
  XNOR2_X1 U977 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n875) );
  XNOR2_X1 U978 ( .A(n875), .B(KEYINPUT45), .ZN(n876) );
  XNOR2_X1 U979 ( .A(n877), .B(n876), .ZN(n881) );
  NAND2_X1 U980 ( .A1(G118), .A2(n885), .ZN(n879) );
  NAND2_X1 U981 ( .A1(G130), .A2(n886), .ZN(n878) );
  NAND2_X1 U982 ( .A1(n879), .A2(n878), .ZN(n880) );
  NOR2_X1 U983 ( .A1(n881), .A2(n880), .ZN(n902) );
  XNOR2_X1 U984 ( .A(KEYINPUT48), .B(KEYINPUT115), .ZN(n884) );
  XNOR2_X1 U985 ( .A(n882), .B(KEYINPUT46), .ZN(n883) );
  XNOR2_X1 U986 ( .A(n884), .B(n883), .ZN(n900) );
  NAND2_X1 U987 ( .A1(G115), .A2(n885), .ZN(n888) );
  NAND2_X1 U988 ( .A1(G127), .A2(n886), .ZN(n887) );
  NAND2_X1 U989 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U990 ( .A(n889), .B(KEYINPUT47), .ZN(n892) );
  NAND2_X1 U991 ( .A1(G103), .A2(n890), .ZN(n891) );
  NAND2_X1 U992 ( .A1(n892), .A2(n891), .ZN(n896) );
  NAND2_X1 U993 ( .A1(n893), .A2(G139), .ZN(n894) );
  XOR2_X1 U994 ( .A(KEYINPUT114), .B(n894), .Z(n895) );
  NOR2_X1 U995 ( .A1(n896), .A2(n895), .ZN(n1000) );
  XNOR2_X1 U996 ( .A(n1000), .B(n897), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n898), .B(G164), .ZN(n899) );
  XNOR2_X1 U998 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U999 ( .A(n902), .B(n901), .ZN(n907) );
  XNOR2_X1 U1000 ( .A(G160), .B(n992), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n903), .B(G162), .ZN(n904) );
  XOR2_X1 U1002 ( .A(n905), .B(n904), .Z(n906) );
  XNOR2_X1 U1003 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n908), .ZN(G395) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(KEYINPUT49), .B(n909), .ZN(n910) );
  NOR2_X1 U1007 ( .A1(G397), .A2(n910), .ZN(n914) );
  NOR2_X1 U1008 ( .A1(G401), .A2(n915), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(KEYINPUT117), .B(n911), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(G395), .A2(n912), .ZN(n913) );
  NAND2_X1 U1011 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(n915), .ZN(G319) );
  INV_X1 U1014 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1015 ( .A(G16), .B(KEYINPUT56), .Z(n939) );
  XNOR2_X1 U1016 ( .A(G1966), .B(G168), .ZN(n917) );
  NAND2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(n918) );
  XNOR2_X1 U1018 ( .A(n918), .B(KEYINPUT57), .ZN(n926) );
  XNOR2_X1 U1019 ( .A(n919), .B(G1348), .ZN(n921) );
  NAND2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n924) );
  XNOR2_X1 U1021 ( .A(G1341), .B(n922), .ZN(n923) );
  NOR2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n937) );
  XNOR2_X1 U1024 ( .A(n927), .B(G1956), .ZN(n929) );
  NAND2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n933) );
  XNOR2_X1 U1026 ( .A(G171), .B(G1961), .ZN(n931) );
  NAND2_X1 U1027 ( .A1(G1971), .A2(G303), .ZN(n930) );
  NAND2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n935) );
  NAND2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1032 ( .A1(n939), .A2(n938), .ZN(n967) );
  XOR2_X1 U1033 ( .A(G1986), .B(G24), .Z(n942) );
  XOR2_X1 U1034 ( .A(G22), .B(KEYINPUT126), .Z(n940) );
  XNOR2_X1 U1035 ( .A(n940), .B(G1971), .ZN(n941) );
  NAND2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n945) );
  XOR2_X1 U1037 ( .A(KEYINPUT127), .B(G1976), .Z(n943) );
  XNOR2_X1 U1038 ( .A(G23), .B(n943), .ZN(n944) );
  NOR2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(KEYINPUT58), .B(n946), .ZN(n950) );
  XNOR2_X1 U1041 ( .A(G1966), .B(G21), .ZN(n948) );
  XNOR2_X1 U1042 ( .A(G5), .B(G1961), .ZN(n947) );
  NOR2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n961) );
  XNOR2_X1 U1045 ( .A(KEYINPUT59), .B(G4), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(n952), .B(n951), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(G20), .B(G1956), .ZN(n953) );
  NOR2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n958) );
  XNOR2_X1 U1049 ( .A(G1341), .B(G19), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(G1981), .B(G6), .ZN(n955) );
  NOR2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1053 ( .A(KEYINPUT60), .B(n959), .ZN(n960) );
  NOR2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1055 ( .A(n962), .B(KEYINPUT61), .ZN(n964) );
  XNOR2_X1 U1056 ( .A(G16), .B(KEYINPUT125), .ZN(n963) );
  NAND2_X1 U1057 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1058 ( .A1(G11), .A2(n965), .ZN(n966) );
  NOR2_X1 U1059 ( .A1(n967), .A2(n966), .ZN(n991) );
  XOR2_X1 U1060 ( .A(G29), .B(KEYINPUT124), .Z(n989) );
  XOR2_X1 U1061 ( .A(G2084), .B(G34), .Z(n968) );
  XNOR2_X1 U1062 ( .A(KEYINPUT54), .B(n968), .ZN(n985) );
  XNOR2_X1 U1063 ( .A(G2090), .B(G35), .ZN(n983) );
  XNOR2_X1 U1064 ( .A(G1991), .B(G25), .ZN(n973) );
  XNOR2_X1 U1065 ( .A(G2067), .B(G26), .ZN(n970) );
  XNOR2_X1 U1066 ( .A(G2072), .B(G33), .ZN(n969) );
  NOR2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1068 ( .A(KEYINPUT121), .B(n971), .ZN(n972) );
  NOR2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1070 ( .A1(G28), .A2(n974), .ZN(n980) );
  XNOR2_X1 U1071 ( .A(G1996), .B(G32), .ZN(n977) );
  XNOR2_X1 U1072 ( .A(n975), .B(G27), .ZN(n976) );
  NOR2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1074 ( .A(KEYINPUT122), .B(n978), .Z(n979) );
  NOR2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1076 ( .A(KEYINPUT53), .B(n981), .ZN(n982) );
  NOR2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(n986), .B(KEYINPUT123), .ZN(n987) );
  XNOR2_X1 U1080 ( .A(n987), .B(KEYINPUT55), .ZN(n988) );
  NAND2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n1021) );
  INV_X1 U1083 ( .A(G29), .ZN(n1019) );
  XNOR2_X1 U1084 ( .A(G160), .B(G2084), .ZN(n993) );
  NAND2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(n996), .B(KEYINPUT118), .ZN(n998) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1089 ( .A(KEYINPUT119), .B(n999), .ZN(n1015) );
  XOR2_X1 U1090 ( .A(G2072), .B(n1000), .Z(n1002) );
  XOR2_X1 U1091 ( .A(G164), .B(G2078), .Z(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(KEYINPUT50), .B(n1003), .ZN(n1007) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1013) );
  XOR2_X1 U1096 ( .A(G2090), .B(KEYINPUT120), .Z(n1008) );
  XNOR2_X1 U1097 ( .A(G162), .B(n1008), .ZN(n1010) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(KEYINPUT51), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(KEYINPUT52), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1103 ( .A1(KEYINPUT55), .A2(n1017), .ZN(n1018) );
  NOR2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1105 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1106 ( .A(KEYINPUT62), .B(n1022), .ZN(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

