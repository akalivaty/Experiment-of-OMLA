//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT0), .A2(G128), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  AND3_X1   g010(.A1(new_n192), .A2(KEYINPUT64), .A3(G146), .ZN(new_n197));
  AOI21_X1  g011(.A(KEYINPUT64), .B1(new_n192), .B2(G146), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n191), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(KEYINPUT0), .B(G128), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n196), .B1(new_n202), .B2(KEYINPUT65), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n199), .A2(new_n204), .A3(new_n201), .ZN(new_n205));
  INV_X1    g019(.A(G104), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT3), .B1(new_n206), .B2(G107), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n208));
  INV_X1    g022(.A(G107), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(G104), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n206), .A2(G107), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n207), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT4), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n213), .A3(G101), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(G101), .ZN(new_n215));
  INV_X1    g029(.A(G101), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n207), .A2(new_n210), .A3(new_n216), .A4(new_n211), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n215), .A2(KEYINPUT4), .A3(new_n217), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n203), .A2(new_n205), .A3(new_n214), .A4(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n206), .A2(G107), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n209), .A2(G104), .ZN(new_n221));
  OAI21_X1  g035(.A(G101), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n217), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G128), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(new_n191), .A3(new_n193), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT64), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n227), .B1(new_n190), .B2(G143), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n192), .A2(KEYINPUT64), .A3(G146), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n228), .A2(new_n229), .B1(G143), .B2(new_n190), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n224), .B1(new_n191), .B2(KEYINPUT1), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n226), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n223), .A2(new_n232), .A3(KEYINPUT10), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT1), .B1(new_n192), .B2(G146), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n234), .A2(G128), .B1(new_n191), .B2(new_n193), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n225), .A2(new_n191), .A3(new_n193), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n217), .B(new_n222), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT10), .ZN(new_n238));
  AOI21_X1  g052(.A(KEYINPUT79), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n237), .A2(KEYINPUT79), .A3(new_n238), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n219), .B(new_n233), .C1(new_n239), .C2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G137), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(KEYINPUT11), .A3(G134), .ZN(new_n243));
  OR2_X1    g057(.A1(KEYINPUT66), .A2(G134), .ZN(new_n244));
  NAND2_X1  g058(.A1(KEYINPUT66), .A2(G134), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n243), .B1(new_n246), .B2(new_n242), .ZN(new_n247));
  AOI21_X1  g061(.A(G137), .B1(new_n244), .B2(new_n245), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT67), .B1(new_n248), .B2(KEYINPUT11), .ZN(new_n249));
  AND2_X1   g063(.A1(KEYINPUT66), .A2(G134), .ZN(new_n250));
  NOR2_X1   g064(.A1(KEYINPUT66), .A2(G134), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n242), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT67), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT11), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n252), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n247), .B1(new_n249), .B2(new_n255), .ZN(new_n256));
  AND2_X1   g070(.A1(KEYINPUT68), .A2(G131), .ZN(new_n257));
  NOR2_X1   g071(.A1(KEYINPUT68), .A2(G131), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n261));
  INV_X1    g075(.A(new_n243), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n250), .A2(new_n251), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n262), .B1(new_n263), .B2(G137), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n252), .A2(new_n253), .A3(new_n254), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n253), .B1(new_n252), .B2(new_n254), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n261), .B(new_n264), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G131), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n256), .A2(new_n261), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n260), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(KEYINPUT80), .B1(new_n241), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT68), .B(G131), .ZN(new_n272));
  AOI211_X1 g086(.A(new_n272), .B(new_n247), .C1(new_n249), .C2(new_n255), .ZN(new_n273));
  INV_X1    g087(.A(G131), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n274), .B1(new_n256), .B2(new_n261), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT69), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n273), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n233), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n218), .A2(new_n214), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT65), .B1(new_n230), .B2(new_n200), .ZN(new_n281));
  INV_X1    g095(.A(new_n196), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n205), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n279), .B1(new_n280), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT80), .ZN(new_n286));
  INV_X1    g100(.A(new_n239), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n237), .A2(KEYINPUT79), .A3(new_n238), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n278), .A2(new_n285), .A3(new_n286), .A4(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n271), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n277), .A2(G131), .A3(new_n267), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n285), .A2(new_n289), .B1(new_n292), .B2(new_n260), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(G110), .B(G140), .ZN(new_n296));
  INV_X1    g110(.A(G953), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n297), .A2(G227), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n296), .B(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n295), .A2(KEYINPUT81), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT81), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n293), .B1(new_n271), .B2(new_n290), .ZN(new_n302));
  INV_X1    g116(.A(new_n299), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n299), .B1(new_n271), .B2(new_n290), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n237), .B1(new_n223), .B2(new_n232), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n270), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT12), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n270), .A2(KEYINPUT12), .A3(new_n306), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n305), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n300), .A2(new_n304), .A3(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G469), .ZN(new_n314));
  INV_X1    g128(.A(G902), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n311), .A2(new_n291), .ZN(new_n317));
  AOI22_X1  g131(.A1(new_n317), .A2(new_n299), .B1(new_n294), .B2(new_n305), .ZN(new_n318));
  OAI21_X1  g132(.A(G469), .B1(new_n318), .B2(G902), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n189), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(G113), .B(G122), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n321), .B(new_n206), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT86), .ZN(new_n323));
  INV_X1    g137(.A(G237), .ZN(new_n324));
  AND4_X1   g138(.A1(G143), .A2(new_n324), .A3(new_n297), .A4(G214), .ZN(new_n325));
  NOR2_X1   g139(.A1(G237), .A2(G953), .ZN(new_n326));
  AOI21_X1  g140(.A(G143), .B1(new_n326), .B2(G214), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n325), .A2(new_n327), .A3(new_n272), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n324), .A2(new_n297), .A3(G214), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n192), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n326), .A2(G143), .A3(G214), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n259), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n323), .B1(new_n328), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G140), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G125), .ZN(new_n335));
  INV_X1    g149(.A(G125), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G140), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n335), .A2(new_n337), .A3(KEYINPUT16), .ZN(new_n338));
  OR3_X1    g152(.A1(new_n336), .A2(KEYINPUT16), .A3(G140), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n339), .A3(G146), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n272), .B1(new_n325), .B2(new_n327), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n330), .A2(new_n259), .A3(new_n331), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(KEYINPUT86), .A3(new_n342), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n335), .A2(new_n337), .A3(KEYINPUT19), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT19), .B1(new_n335), .B2(new_n337), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n190), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n333), .A2(new_n340), .A3(new_n343), .A4(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(G125), .B(G140), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n348), .B(new_n190), .ZN(new_n349));
  NAND2_X1  g163(.A1(KEYINPUT18), .A2(G131), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n330), .A2(new_n331), .A3(new_n350), .ZN(new_n351));
  OAI211_X1 g165(.A(KEYINPUT18), .B(G131), .C1(new_n325), .C2(new_n327), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n349), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n322), .B1(new_n347), .B2(new_n353), .ZN(new_n354));
  NOR3_X1   g168(.A1(new_n328), .A2(new_n332), .A3(KEYINPUT17), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n338), .A2(new_n339), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n190), .ZN(new_n357));
  OAI211_X1 g171(.A(KEYINPUT17), .B(new_n272), .C1(new_n325), .C2(new_n327), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n340), .A3(new_n358), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n322), .B(new_n353), .C1(new_n355), .C2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n354), .A2(new_n361), .ZN(new_n362));
  NOR4_X1   g176(.A1(new_n362), .A2(KEYINPUT20), .A3(G475), .A4(G902), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT87), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n364), .B1(new_n354), .B2(new_n361), .ZN(new_n365));
  AND3_X1   g179(.A1(new_n349), .A2(new_n351), .A3(new_n352), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n346), .A2(new_n340), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT86), .B1(new_n341), .B2(new_n342), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n366), .B1(new_n369), .B2(new_n343), .ZN(new_n370));
  OAI211_X1 g184(.A(KEYINPUT87), .B(new_n360), .C1(new_n370), .C2(new_n322), .ZN(new_n371));
  NOR2_X1   g185(.A1(G475), .A2(G902), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n365), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n363), .B1(KEYINPUT20), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G475), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n353), .B1(new_n355), .B2(new_n359), .ZN(new_n376));
  XOR2_X1   g190(.A(new_n376), .B(new_n322), .Z(new_n377));
  AOI21_X1  g191(.A(new_n375), .B1(new_n377), .B2(new_n315), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(G116), .B(G122), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n380), .B(new_n209), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n192), .A2(G128), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n224), .A2(G143), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n263), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT13), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n192), .A2(KEYINPUT13), .A3(G128), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n387), .A3(new_n383), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT88), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n388), .A2(new_n389), .A3(G134), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n389), .B1(new_n388), .B2(G134), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n381), .B(new_n384), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G116), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(KEYINPUT14), .A3(G122), .ZN(new_n394));
  INV_X1    g208(.A(new_n380), .ZN(new_n395));
  OAI211_X1 g209(.A(G107), .B(new_n394), .C1(new_n395), .C2(KEYINPUT14), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n382), .A2(new_n383), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n246), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n384), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n380), .A2(new_n209), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n396), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT89), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT89), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n396), .A2(new_n399), .A3(new_n403), .A4(new_n400), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n392), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G217), .ZN(new_n406));
  NOR3_X1   g220(.A1(new_n187), .A2(new_n406), .A3(G953), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n392), .A2(new_n402), .A3(new_n404), .A4(new_n407), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n315), .ZN(new_n412));
  INV_X1    g226(.A(G478), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(KEYINPUT15), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n411), .B(new_n315), .C1(KEYINPUT15), .C2(new_n413), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n379), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G952), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n418), .A2(KEYINPUT90), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n418), .A2(KEYINPUT90), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n297), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n421), .B1(G234), .B2(G237), .ZN(new_n422));
  XOR2_X1   g236(.A(KEYINPUT21), .B(G898), .Z(new_n423));
  XNOR2_X1  g237(.A(new_n423), .B(KEYINPUT92), .ZN(new_n424));
  NAND2_X1  g238(.A1(G234), .A2(G237), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(G902), .A3(G953), .ZN(new_n426));
  XOR2_X1   g240(.A(new_n426), .B(KEYINPUT91), .Z(new_n427));
  AOI21_X1  g241(.A(new_n422), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(G214), .B1(G237), .B2(G902), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n283), .A2(G125), .ZN(new_n431));
  OR2_X1    g245(.A1(new_n232), .A2(G125), .ZN(new_n432));
  INV_X1    g246(.A(G224), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n433), .A2(G953), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n431), .A2(new_n432), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n435), .B1(new_n431), .B2(new_n432), .ZN(new_n437));
  OR2_X1    g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(G110), .B(G122), .ZN(new_n439));
  OAI21_X1  g253(.A(KEYINPUT71), .B1(new_n393), .B2(G119), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT71), .ZN(new_n441));
  INV_X1    g255(.A(G119), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n441), .A2(new_n442), .A3(G116), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n393), .A2(G119), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n440), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT2), .ZN(new_n446));
  INV_X1    g260(.A(G113), .ZN(new_n447));
  OAI21_X1  g261(.A(KEYINPUT70), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT70), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(KEYINPUT2), .A3(G113), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(KEYINPUT2), .A2(G113), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n445), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI22_X1  g267(.A1(new_n448), .A2(new_n450), .B1(new_n446), .B2(new_n447), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n440), .A2(new_n443), .A3(new_n444), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(new_n218), .A3(new_n214), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n440), .A2(new_n443), .A3(KEYINPUT5), .A4(new_n444), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n393), .A2(G119), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT5), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n447), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n223), .A2(new_n456), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n439), .B1(new_n458), .B2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT83), .B(KEYINPUT6), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n458), .A2(new_n464), .ZN(new_n468));
  INV_X1    g282(.A(new_n439), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(KEYINPUT82), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n458), .A2(new_n439), .A3(new_n464), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(KEYINPUT6), .A3(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n465), .A2(KEYINPUT82), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n438), .B(new_n467), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n454), .A2(new_n455), .B1(new_n459), .B2(new_n462), .ZN(new_n475));
  OR3_X1    g289(.A1(new_n475), .A2(KEYINPUT85), .A3(new_n223), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT84), .ZN(new_n477));
  OR2_X1    g291(.A1(new_n462), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n462), .A2(new_n477), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n478), .A2(new_n459), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(new_n223), .A3(new_n456), .ZN(new_n481));
  OAI21_X1  g295(.A(KEYINPUT85), .B1(new_n475), .B2(new_n223), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n476), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n439), .B(KEYINPUT8), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n436), .A2(KEYINPUT7), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI22_X1  g299(.A1(new_n431), .A2(new_n432), .B1(KEYINPUT7), .B2(new_n435), .ZN(new_n486));
  INV_X1    g300(.A(new_n468), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n486), .B1(new_n487), .B2(new_n439), .ZN(new_n488));
  AOI21_X1  g302(.A(G902), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(G210), .B1(G237), .B2(G902), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n474), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n490), .B1(new_n474), .B2(new_n489), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n429), .B(new_n430), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n417), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n320), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(KEYINPUT93), .ZN(new_n496));
  NOR2_X1   g310(.A1(G472), .A2(G902), .ZN(new_n497));
  XOR2_X1   g311(.A(new_n497), .B(KEYINPUT74), .Z(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n499), .A2(KEYINPUT32), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n283), .B1(new_n292), .B2(new_n260), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n242), .A2(G134), .ZN(new_n502));
  OAI21_X1  g316(.A(G131), .B1(new_n248), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n232), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n273), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n457), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT72), .ZN(new_n507));
  INV_X1    g321(.A(new_n457), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n508), .B1(new_n273), .B2(new_n504), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n507), .B1(new_n501), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n509), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n511), .B(KEYINPUT72), .C1(new_n278), .C2(new_n283), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n506), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT28), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n501), .A2(new_n509), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n515), .A2(KEYINPUT28), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n326), .A2(G210), .ZN(new_n519));
  XOR2_X1   g333(.A(new_n519), .B(KEYINPUT27), .Z(new_n520));
  XNOR2_X1  g334(.A(KEYINPUT26), .B(G101), .ZN(new_n521));
  XOR2_X1   g335(.A(new_n520), .B(new_n521), .Z(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n510), .A2(new_n512), .A3(new_n522), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT30), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n270), .A2(new_n284), .ZN(new_n527));
  INV_X1    g341(.A(new_n505), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AOI211_X1 g343(.A(KEYINPUT30), .B(new_n505), .C1(new_n270), .C2(new_n284), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n457), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n525), .A2(new_n531), .A3(KEYINPUT31), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT31), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT30), .B1(new_n501), .B2(new_n505), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n527), .A2(new_n526), .A3(new_n528), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n508), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n510), .A2(new_n512), .A3(new_n522), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n533), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n532), .A2(new_n538), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n524), .A2(KEYINPUT73), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(KEYINPUT73), .B1(new_n524), .B2(new_n539), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n500), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n514), .A2(KEYINPUT75), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT75), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n513), .A2(new_n544), .A3(KEYINPUT28), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT29), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n523), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n543), .A2(new_n517), .A3(new_n545), .A4(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n518), .A2(new_n523), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n510), .A2(new_n512), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n536), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n546), .B1(new_n551), .B2(new_n522), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n548), .B(new_n315), .C1(new_n549), .C2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(G472), .ZN(new_n554));
  AOI21_X1  g368(.A(KEYINPUT31), .B1(new_n525), .B2(new_n531), .ZN(new_n555));
  NOR3_X1   g369(.A1(new_n536), .A2(new_n537), .A3(new_n533), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n516), .B1(new_n513), .B2(KEYINPUT28), .ZN(new_n557));
  OAI22_X1  g371(.A1(new_n555), .A2(new_n556), .B1(new_n557), .B2(new_n522), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT73), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n524), .A2(KEYINPUT73), .A3(new_n539), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n498), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n542), .B(new_n554), .C1(new_n562), .C2(KEYINPUT32), .ZN(new_n563));
  OAI21_X1  g377(.A(KEYINPUT23), .B1(new_n224), .B2(G119), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT76), .B1(new_n442), .B2(G128), .ZN(new_n565));
  XOR2_X1   g379(.A(new_n564), .B(new_n565), .Z(new_n566));
  XNOR2_X1  g380(.A(G119), .B(G128), .ZN(new_n567));
  XOR2_X1   g381(.A(KEYINPUT24), .B(G110), .Z(new_n568));
  OAI22_X1  g382(.A1(new_n566), .A2(G110), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n348), .A2(new_n190), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(new_n570), .A3(new_n340), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n566), .A2(G110), .B1(new_n567), .B2(new_n568), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n357), .A2(new_n340), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n297), .A2(G221), .A3(G234), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(KEYINPUT77), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT22), .B(G137), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n571), .A2(new_n574), .A3(new_n579), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT25), .ZN(new_n583));
  AOI21_X1  g397(.A(G902), .B1(new_n583), .B2(KEYINPUT78), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n581), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n583), .A2(KEYINPUT78), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n406), .B1(G234), .B2(new_n315), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n590), .B1(new_n585), .B2(new_n587), .ZN(new_n591));
  OR2_X1    g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n581), .A2(new_n582), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n590), .A2(G902), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n496), .A2(new_n563), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(G101), .ZN(G3));
  OAI21_X1  g413(.A(new_n315), .B1(new_n540), .B2(new_n541), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n562), .B1(G472), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n316), .A2(new_n319), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n188), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(new_n596), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g419(.A(new_n605), .B(KEYINPUT94), .Z(new_n606));
  NOR2_X1   g420(.A1(new_n413), .A2(G902), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n408), .A2(KEYINPUT95), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n610), .B1(new_n405), .B2(KEYINPUT96), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n410), .A2(KEYINPUT96), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n405), .A2(KEYINPUT96), .A3(new_n610), .ZN(new_n614));
  OAI21_X1  g428(.A(KEYINPUT33), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OR2_X1    g429(.A1(new_n411), .A2(KEYINPUT33), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n608), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(G478), .B1(new_n411), .B2(new_n315), .ZN(new_n618));
  OAI22_X1  g432(.A1(new_n374), .A2(new_n378), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n493), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n606), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT34), .B(G104), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G6));
  OAI21_X1  g438(.A(new_n430), .B1(new_n491), .B2(new_n492), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n373), .A2(KEYINPUT20), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT20), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n365), .A2(new_n371), .A3(new_n628), .A4(new_n372), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n378), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT97), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n428), .B1(new_n415), .B2(new_n416), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n630), .A2(new_n632), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(KEYINPUT97), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n626), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n606), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT98), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT35), .B(G107), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  INV_X1    g454(.A(new_n594), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n575), .A2(KEYINPUT99), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT99), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n571), .A2(new_n643), .A3(new_n574), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n645), .B1(KEYINPUT36), .B2(new_n580), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n580), .A2(KEYINPUT36), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n642), .A2(new_n647), .A3(new_n644), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n641), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(KEYINPUT100), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  OAI22_X1  g465(.A1(new_n649), .A2(KEYINPUT100), .B1(new_n589), .B2(new_n591), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n496), .A2(new_n601), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT37), .B(G110), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G12));
  INV_X1    g471(.A(new_n563), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n603), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n654), .A2(new_n626), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n415), .A2(new_n416), .ZN(new_n661));
  INV_X1    g475(.A(G900), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n422), .B1(new_n427), .B2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n630), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n659), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G128), .ZN(G30));
  XOR2_X1   g482(.A(new_n663), .B(KEYINPUT39), .Z(new_n669));
  NAND2_X1  g483(.A1(new_n320), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n670), .B(KEYINPUT102), .Z(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  OR2_X1    g486(.A1(new_n672), .A2(KEYINPUT40), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(KEYINPUT40), .ZN(new_n674));
  AOI21_X1  g488(.A(KEYINPUT101), .B1(new_n513), .B2(new_n523), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n513), .A2(KEYINPUT101), .A3(new_n523), .ZN(new_n676));
  AOI211_X1 g490(.A(new_n675), .B(new_n676), .C1(new_n531), .C2(new_n525), .ZN(new_n677));
  OAI21_X1  g491(.A(G472), .B1(new_n677), .B2(G902), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n542), .B(new_n678), .C1(new_n562), .C2(KEYINPUT32), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n661), .B1(new_n374), .B2(new_n378), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n492), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n474), .A2(new_n489), .A3(new_n490), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT38), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n686), .A2(new_n430), .A3(new_n653), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n673), .A2(new_n674), .A3(new_n682), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G143), .ZN(G45));
  NOR2_X1   g503(.A1(new_n619), .A2(new_n663), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n660), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n659), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G146), .ZN(G48));
  NOR2_X1   g508(.A1(new_n658), .A2(new_n596), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n313), .A2(new_n315), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(G469), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n316), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n698), .A2(new_n621), .A3(new_n189), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(KEYINPUT41), .B(G113), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT103), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n700), .B(new_n702), .ZN(G15));
  NOR3_X1   g517(.A1(new_n698), .A2(new_n636), .A3(new_n189), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n695), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G116), .ZN(G18));
  AND3_X1   g520(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n314), .B1(new_n313), .B2(new_n315), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n709), .A2(KEYINPUT104), .A3(new_n188), .A4(new_n626), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n697), .A2(new_n188), .A3(new_n316), .A4(new_n626), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT104), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n653), .A2(new_n417), .A3(new_n428), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n714), .A2(new_n563), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  NAND3_X1  g531(.A1(new_n543), .A2(new_n517), .A3(new_n545), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n523), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n498), .B1(new_n719), .B2(new_n539), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n720), .B1(new_n600), .B2(G472), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n698), .A2(new_n189), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n625), .A2(new_n681), .A3(new_n428), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n721), .A2(new_n597), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G122), .ZN(G24));
  NAND4_X1  g539(.A1(new_n714), .A2(new_n654), .A3(new_n690), .A4(new_n721), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G125), .ZN(G27));
  INV_X1    g541(.A(new_n430), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n685), .A2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n603), .A2(new_n691), .A3(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n563), .A2(new_n597), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT42), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n563), .A2(KEYINPUT42), .A3(new_n597), .A4(new_n731), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G131), .ZN(G33));
  XNOR2_X1  g551(.A(new_n665), .B(KEYINPUT105), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n603), .A2(new_n738), .A3(new_n730), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n542), .A2(new_n554), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n560), .A2(new_n561), .ZN(new_n741));
  AOI21_X1  g555(.A(KEYINPUT32), .B1(new_n741), .B2(new_n499), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n597), .B(new_n739), .C1(new_n740), .C2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G134), .ZN(G36));
  OR2_X1    g558(.A1(new_n318), .A2(KEYINPUT45), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n318), .A2(KEYINPUT45), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(G469), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(G469), .A2(G902), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT46), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n707), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(new_n750), .B2(new_n749), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n188), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n669), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(KEYINPUT106), .ZN(new_n756));
  INV_X1    g570(.A(new_n601), .ZN(new_n757));
  OR2_X1    g571(.A1(new_n617), .A2(new_n618), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n379), .ZN(new_n759));
  XOR2_X1   g573(.A(new_n759), .B(KEYINPUT43), .Z(new_n760));
  NAND3_X1  g574(.A1(new_n757), .A2(new_n654), .A3(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT44), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n730), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n763), .B1(new_n762), .B2(new_n761), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n756), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(new_n242), .ZN(G39));
  NAND2_X1  g580(.A1(new_n754), .A2(KEYINPUT47), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT47), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n753), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  NOR4_X1   g584(.A1(new_n563), .A2(new_n597), .A3(new_n691), .A4(new_n730), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT107), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n770), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G140), .ZN(G42));
  INV_X1    g590(.A(new_n721), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n760), .A2(new_n422), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n777), .A2(new_n778), .A3(new_n596), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n779), .A2(new_n729), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n767), .A2(KEYINPUT116), .A3(new_n769), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n781), .B1(new_n188), .B2(new_n698), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT116), .B1(new_n767), .B2(new_n769), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n780), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  XOR2_X1   g598(.A(new_n784), .B(KEYINPUT117), .Z(new_n785));
  NAND2_X1  g599(.A1(new_n722), .A2(new_n729), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n778), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n787), .A2(new_n654), .A3(new_n721), .ZN(new_n788));
  XOR2_X1   g602(.A(new_n788), .B(KEYINPUT119), .Z(new_n789));
  NAND4_X1  g603(.A1(new_n722), .A2(new_n422), .A3(new_n597), .A4(new_n729), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT120), .ZN(new_n791));
  OR3_X1    g605(.A1(new_n790), .A2(new_n679), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n791), .B1(new_n790), .B2(new_n679), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n758), .A2(new_n378), .A3(new_n374), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NOR4_X1   g609(.A1(new_n686), .A2(new_n698), .A3(new_n189), .A4(new_n430), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT118), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n797), .A2(new_n779), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n798), .A2(KEYINPUT50), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n798), .A2(KEYINPUT50), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n789), .B(new_n795), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT121), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT51), .B1(new_n785), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n695), .A2(new_n787), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT48), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n421), .B1(new_n779), .B2(new_n714), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n792), .A2(new_n793), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n698), .A2(new_n188), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n780), .B1(new_n770), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT51), .ZN(new_n811));
  OAI221_X1 g625(.A(new_n807), .B1(new_n619), .B2(new_n808), .C1(new_n801), .C2(new_n811), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n803), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT112), .ZN(new_n814));
  XOR2_X1   g628(.A(new_n663), .B(KEYINPUT111), .Z(new_n815));
  NAND2_X1  g629(.A1(new_n653), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n814), .B1(new_n603), .B2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n320), .A2(new_n653), .A3(KEYINPUT112), .A4(new_n815), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n681), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n819), .A2(new_n626), .A3(new_n679), .A4(new_n820), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n563), .B(new_n320), .C1(new_n666), .C2(new_n692), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n821), .A2(new_n726), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT113), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n825), .B(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n417), .B1(new_n758), .B2(new_n379), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(new_n493), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n601), .A2(new_n604), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n598), .A2(new_n655), .A3(new_n832), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n563), .B(new_n597), .C1(new_n699), .C2(new_n704), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n834), .A2(new_n716), .A3(new_n724), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT109), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT109), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n834), .A2(new_n716), .A3(new_n724), .A4(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n833), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n721), .A2(new_n654), .A3(new_n731), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n630), .A2(new_n664), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n653), .A2(new_n661), .A3(new_n841), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n842), .A2(new_n320), .A3(new_n729), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n563), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n743), .A2(new_n840), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT110), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT110), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n743), .A2(new_n840), .A3(new_n844), .A4(new_n847), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n846), .A2(new_n736), .A3(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n828), .A2(new_n829), .A3(new_n839), .A4(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT52), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n823), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n821), .A2(new_n726), .A3(new_n822), .A4(KEYINPUT52), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n839), .A2(new_n849), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT53), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n850), .A2(KEYINPUT54), .A3(new_n856), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n833), .A2(new_n835), .A3(new_n829), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n849), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n827), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT115), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n855), .A2(new_n862), .A3(new_n829), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n862), .B1(new_n855), .B2(new_n829), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n857), .B1(new_n865), .B2(KEYINPUT54), .ZN(new_n866));
  OAI22_X1  g680(.A1(new_n813), .A2(new_n866), .B1(G952), .B2(G953), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n698), .A2(KEYINPUT49), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n698), .A2(KEYINPUT49), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n597), .A2(new_n188), .A3(new_n430), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n686), .A2(new_n870), .A3(new_n759), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n680), .A2(new_n868), .A3(new_n869), .A4(new_n871), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n872), .B(KEYINPUT108), .Z(new_n873));
  NAND2_X1  g687(.A1(new_n867), .A2(new_n873), .ZN(G75));
  NAND2_X1  g688(.A1(new_n855), .A2(new_n829), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT115), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n855), .A2(new_n862), .A3(new_n829), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n860), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT123), .B1(new_n878), .B2(new_n315), .ZN(new_n879));
  INV_X1    g693(.A(new_n490), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT123), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n865), .A2(new_n881), .A3(G902), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n467), .B1(new_n472), .B2(new_n473), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(new_n438), .ZN(new_n885));
  XOR2_X1   g699(.A(KEYINPUT122), .B(KEYINPUT55), .Z(new_n886));
  XNOR2_X1  g700(.A(new_n885), .B(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n887), .A2(KEYINPUT56), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n297), .A2(G952), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n865), .A2(G210), .A3(G902), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT56), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n890), .B1(new_n893), .B2(new_n887), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n889), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(KEYINPUT124), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT124), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n889), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n896), .A2(new_n898), .ZN(G51));
  XNOR2_X1  g713(.A(new_n865), .B(KEYINPUT54), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n748), .B(KEYINPUT57), .Z(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n313), .ZN(new_n903));
  INV_X1    g717(.A(new_n747), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n879), .A2(new_n904), .A3(new_n882), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n890), .B1(new_n903), .B2(new_n905), .ZN(G54));
  AND2_X1   g720(.A1(new_n365), .A2(new_n371), .ZN(new_n907));
  AND2_X1   g721(.A1(KEYINPUT58), .A2(G475), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n879), .A2(new_n907), .A3(new_n882), .A4(new_n908), .ZN(new_n909));
  OR2_X1    g723(.A1(new_n909), .A2(KEYINPUT125), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(KEYINPUT125), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n879), .A2(new_n882), .A3(new_n908), .ZN(new_n912));
  INV_X1    g726(.A(new_n907), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n890), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n910), .A2(new_n911), .A3(new_n914), .ZN(G60));
  NAND2_X1  g729(.A1(new_n615), .A2(new_n616), .ZN(new_n916));
  XNOR2_X1  g730(.A(KEYINPUT126), .B(KEYINPUT59), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n413), .A2(new_n315), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n917), .B(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n916), .B1(new_n866), .B2(new_n919), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n916), .A2(new_n919), .ZN(new_n921));
  AOI211_X1 g735(.A(new_n890), .B(new_n920), .C1(new_n900), .C2(new_n921), .ZN(G63));
  NAND2_X1  g736(.A1(G217), .A2(G902), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT60), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n878), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n646), .A2(new_n648), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n890), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n927), .B(new_n928), .C1(new_n593), .C2(new_n925), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT61), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(G66));
  OAI21_X1  g745(.A(G953), .B1(new_n424), .B2(new_n433), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n932), .B1(new_n839), .B2(G953), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n884), .B1(G898), .B2(new_n297), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(G69));
  NAND3_X1  g749(.A1(new_n695), .A2(new_n626), .A3(new_n820), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n756), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n726), .A2(new_n822), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n775), .B1(new_n756), .B2(new_n764), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n939), .A2(new_n941), .A3(new_n736), .A4(new_n743), .ZN(new_n942));
  OR2_X1    g756(.A1(new_n942), .A2(G953), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n943), .B1(new_n662), .B2(new_n297), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n534), .A2(new_n535), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n344), .A2(new_n345), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(G227), .A2(G900), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(G953), .ZN(new_n950));
  INV_X1    g764(.A(new_n688), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n951), .A2(new_n938), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT62), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n830), .A2(new_n730), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n695), .A2(new_n671), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n941), .A2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n953), .A2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n947), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n958), .A2(new_n297), .A3(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n948), .A2(new_n950), .A3(new_n960), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n944), .A2(G953), .A3(new_n949), .A4(new_n947), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n961), .A2(new_n962), .ZN(G72));
  NAND2_X1  g777(.A1(G472), .A2(G902), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT63), .Z(new_n965));
  INV_X1    g779(.A(new_n839), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n965), .B1(new_n958), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n551), .A2(new_n523), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n536), .A2(new_n550), .A3(new_n522), .ZN(new_n970));
  INV_X1    g784(.A(new_n965), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n968), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n850), .A2(new_n856), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n965), .B1(new_n942), .B2(new_n966), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n890), .B1(new_n974), .B2(new_n970), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n969), .A2(new_n973), .A3(new_n975), .ZN(G57));
endmodule


