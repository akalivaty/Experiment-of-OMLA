//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT2), .B(G113), .Z(new_n188));
  XNOR2_X1  g002(.A(G116), .B(G119), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT2), .B(G113), .ZN(new_n191));
  INV_X1    g005(.A(G116), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G119), .ZN(new_n193));
  INV_X1    g007(.A(G119), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(G116), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n191), .B1(new_n193), .B2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n190), .A2(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(new_n197), .B(KEYINPUT68), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n201), .A2(new_n203), .A3(KEYINPUT0), .A4(G128), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(G143), .B(G146), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n207), .A2(KEYINPUT65), .A3(KEYINPUT0), .A4(G128), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n210), .B1(new_n200), .B2(G143), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n202), .A2(KEYINPUT64), .A3(G146), .ZN(new_n212));
  AOI22_X1  g026(.A1(new_n211), .A2(new_n212), .B1(G143), .B2(new_n200), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT0), .B(G128), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G137), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(G134), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(KEYINPUT11), .A3(G134), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT67), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n217), .A2(KEYINPUT67), .A3(KEYINPUT11), .A4(G134), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n218), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G131), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT11), .ZN(new_n225));
  INV_X1    g039(.A(G134), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(G137), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI211_X1 g043(.A(KEYINPUT66), .B(new_n225), .C1(new_n226), .C2(G137), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  AND3_X1   g045(.A1(new_n223), .A2(new_n224), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n224), .B1(new_n223), .B2(new_n231), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n216), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n223), .A2(new_n224), .A3(new_n231), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT1), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n207), .A2(new_n236), .A3(G128), .ZN(new_n237));
  INV_X1    g051(.A(G128), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n238), .B1(new_n201), .B2(KEYINPUT1), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n237), .B1(new_n213), .B2(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n226), .A2(G137), .ZN(new_n241));
  OAI21_X1  g055(.A(G131), .B1(new_n241), .B2(new_n218), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n235), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n234), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n199), .B1(new_n244), .B2(KEYINPUT69), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n234), .A2(new_n246), .A3(new_n243), .ZN(new_n247));
  AOI21_X1  g061(.A(KEYINPUT28), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n244), .A2(new_n199), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n234), .A2(new_n198), .A3(new_n243), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n248), .B1(KEYINPUT28), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G237), .ZN(new_n253));
  INV_X1    g067(.A(G953), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n254), .A3(G210), .ZN(new_n255));
  INV_X1    g069(.A(G101), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n258));
  XOR2_X1   g072(.A(new_n257), .B(new_n258), .Z(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT29), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(G902), .B1(new_n252), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n244), .A2(KEYINPUT69), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(new_n198), .A3(new_n247), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT28), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n250), .ZN(new_n268));
  AOI22_X1  g082(.A1(new_n234), .A2(new_n243), .B1(new_n196), .B2(new_n190), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT28), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n267), .A2(new_n259), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT30), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n206), .B(new_n208), .C1(new_n213), .C2(new_n214), .ZN(new_n273));
  INV_X1    g087(.A(new_n218), .ZN(new_n274));
  AOI21_X1  g088(.A(KEYINPUT67), .B1(new_n241), .B2(KEYINPUT11), .ZN(new_n275));
  INV_X1    g089(.A(new_n222), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n230), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n217), .A2(G134), .ZN(new_n279));
  AOI21_X1  g093(.A(KEYINPUT66), .B1(new_n279), .B2(new_n225), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(G131), .B1(new_n277), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n273), .B1(new_n282), .B2(new_n235), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n235), .A2(new_n240), .A3(new_n242), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n272), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n234), .A2(KEYINPUT30), .A3(new_n243), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(new_n286), .A3(new_n197), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n250), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n260), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n271), .A2(new_n261), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n187), .B1(new_n263), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G902), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n187), .A2(new_n293), .A3(KEYINPUT71), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT71), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n295), .B1(G472), .B2(G902), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n287), .A2(new_n259), .A3(new_n250), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT31), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT31), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n287), .A2(new_n301), .A3(new_n259), .A4(new_n250), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n259), .B1(new_n267), .B2(new_n270), .ZN(new_n304));
  OAI21_X1  g118(.A(KEYINPUT70), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n269), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n266), .B1(new_n306), .B2(new_n250), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n260), .B1(new_n248), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT70), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n308), .A2(new_n309), .A3(new_n300), .A4(new_n302), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n298), .B1(new_n305), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(KEYINPUT72), .B1(new_n311), .B2(KEYINPUT32), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT32), .ZN(new_n313));
  AOI211_X1 g127(.A(new_n313), .B(new_n298), .C1(new_n305), .C2(new_n310), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n305), .A2(new_n310), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n297), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n317), .A2(KEYINPUT72), .A3(new_n313), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n292), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  XOR2_X1   g133(.A(KEYINPUT24), .B(G110), .Z(new_n320));
  XNOR2_X1  g134(.A(new_n320), .B(KEYINPUT74), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n238), .A2(G119), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT73), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n194), .A2(G128), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT73), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n324), .B1(new_n322), .B2(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n322), .B(KEYINPUT23), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n325), .ZN(new_n329));
  OAI22_X1  g143(.A1(new_n321), .A2(new_n327), .B1(new_n329), .B2(G110), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI221_X1 g146(.A(KEYINPUT77), .B1(new_n329), .B2(G110), .C1(new_n321), .C2(new_n327), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT16), .ZN(new_n334));
  INV_X1    g148(.A(G125), .ZN(new_n335));
  OAI21_X1  g149(.A(G140), .B1(new_n335), .B2(KEYINPUT75), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT75), .ZN(new_n337));
  INV_X1    g151(.A(G140), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(new_n338), .A3(G125), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n334), .B1(new_n336), .B2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(KEYINPUT16), .B1(new_n338), .B2(G125), .ZN(new_n341));
  OAI21_X1  g155(.A(G146), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n338), .A2(G125), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n335), .A2(G140), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n344), .A3(new_n200), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n332), .A2(new_n333), .A3(new_n342), .A4(new_n345), .ZN(new_n346));
  AOI22_X1  g160(.A1(new_n321), .A2(new_n327), .B1(new_n329), .B2(G110), .ZN(new_n347));
  INV_X1    g161(.A(new_n342), .ZN(new_n348));
  NOR3_X1   g162(.A1(new_n340), .A2(G146), .A3(new_n341), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT76), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT76), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n347), .B(new_n352), .C1(new_n348), .C2(new_n349), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n346), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT22), .B(G137), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n254), .A2(G221), .A3(G234), .ZN(new_n356));
  XOR2_X1   g170(.A(new_n355), .B(new_n356), .Z(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n346), .A2(new_n351), .A3(new_n353), .A4(new_n357), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n293), .A3(new_n360), .ZN(new_n361));
  AND2_X1   g175(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G217), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n364), .B1(G234), .B2(new_n293), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT78), .B(KEYINPUT25), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n363), .B(new_n365), .C1(new_n361), .C2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT79), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n359), .A2(new_n360), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n365), .A2(G902), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n367), .A2(new_n368), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n368), .B1(new_n367), .B2(new_n371), .ZN(new_n373));
  OR2_X1    g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(G210), .B1(G237), .B2(G902), .ZN(new_n375));
  OR2_X1    g189(.A1(new_n240), .A2(G125), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n273), .A2(G125), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT86), .ZN(new_n379));
  OR2_X1    g193(.A1(new_n379), .A2(KEYINPUT7), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n254), .A2(G224), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(KEYINPUT7), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n378), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT87), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT7), .A4(new_n381), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT87), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n378), .A2(new_n387), .A3(new_n383), .ZN(new_n388));
  XOR2_X1   g202(.A(G110), .B(G122), .Z(new_n389));
  XOR2_X1   g203(.A(new_n389), .B(KEYINPUT8), .Z(new_n390));
  INV_X1    g204(.A(G104), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G107), .ZN(new_n392));
  INV_X1    g206(.A(G107), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G104), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n256), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n393), .A2(KEYINPUT3), .A3(G104), .ZN(new_n396));
  AOI21_X1  g210(.A(KEYINPUT3), .B1(new_n393), .B2(G104), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n256), .B(new_n392), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT80), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n393), .A2(G104), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT3), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n401), .B1(new_n391), .B2(G107), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n393), .A2(KEYINPUT3), .A3(G104), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n400), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT80), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(new_n405), .A3(new_n256), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n395), .B1(new_n399), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n189), .A2(KEYINPUT5), .ZN(new_n408));
  INV_X1    g222(.A(G113), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT5), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n409), .B1(new_n193), .B2(new_n410), .ZN(new_n411));
  AOI22_X1  g225(.A1(new_n408), .A2(new_n411), .B1(new_n188), .B2(new_n189), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n407), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n395), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n402), .A2(new_n403), .ZN(new_n415));
  AND4_X1   g229(.A1(new_n405), .A2(new_n415), .A3(new_n256), .A4(new_n392), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n405), .B1(new_n404), .B2(new_n256), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n414), .B(new_n412), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n390), .B1(new_n413), .B2(new_n419), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n385), .A2(new_n386), .A3(new_n388), .A4(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n389), .ZN(new_n422));
  OAI21_X1  g236(.A(KEYINPUT4), .B1(new_n404), .B2(new_n256), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n423), .B1(new_n406), .B2(new_n399), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n415), .A2(new_n392), .ZN(new_n425));
  XOR2_X1   g239(.A(KEYINPUT81), .B(KEYINPUT4), .Z(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(G101), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n197), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n418), .B(new_n422), .C1(new_n424), .C2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT84), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n425), .A2(G101), .ZN(new_n431));
  OAI211_X1 g245(.A(KEYINPUT4), .B(new_n431), .C1(new_n416), .C2(new_n417), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n427), .A2(new_n197), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT84), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n434), .A2(new_n435), .A3(new_n422), .A4(new_n418), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n430), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n293), .B1(new_n421), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n418), .B1(new_n424), .B2(new_n428), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT6), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(KEYINPUT83), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n440), .A2(new_n389), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n442), .B1(new_n440), .B2(new_n389), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n430), .A2(new_n436), .A3(KEYINPUT6), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n378), .B(new_n381), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(KEYINPUT85), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT85), .ZN(new_n451));
  AOI211_X1 g265(.A(new_n451), .B(new_n448), .C1(new_n445), .C2(new_n446), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n375), .B(new_n439), .C1(new_n450), .C2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(KEYINPUT88), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n430), .A2(KEYINPUT6), .A3(new_n436), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n432), .A2(new_n433), .B1(new_n407), .B2(new_n412), .ZN(new_n456));
  OAI22_X1  g270(.A1(new_n456), .A2(new_n422), .B1(KEYINPUT83), .B2(new_n441), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n440), .A2(new_n389), .A3(new_n442), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n449), .B1(new_n455), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n451), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n447), .A2(KEYINPUT85), .A3(new_n449), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n375), .B1(new_n463), .B2(new_n439), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n454), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(G214), .B1(G237), .B2(G902), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n438), .B1(new_n461), .B2(new_n462), .ZN(new_n468));
  NOR3_X1   g282(.A1(new_n468), .A2(KEYINPUT88), .A3(new_n375), .ZN(new_n469));
  NOR3_X1   g283(.A1(new_n465), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT93), .ZN(new_n471));
  OR3_X1    g285(.A1(new_n348), .A2(new_n471), .A3(new_n349), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n471), .B1(new_n348), .B2(new_n349), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n253), .A2(new_n254), .A3(G214), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(G143), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n475), .A2(new_n224), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT17), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n474), .B(new_n202), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G131), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n475), .A2(new_n224), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT17), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n472), .A2(new_n473), .A3(new_n477), .A4(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT18), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n475), .B1(new_n484), .B2(new_n224), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n336), .A2(new_n339), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(G146), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n345), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n485), .B(new_n488), .C1(new_n484), .C2(new_n479), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT89), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n476), .A2(KEYINPUT18), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n492), .A2(new_n488), .A3(new_n485), .A4(KEYINPUT89), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(G113), .B(G122), .ZN(new_n495));
  XNOR2_X1  g309(.A(KEYINPUT92), .B(G104), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n495), .B(new_n496), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n483), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n497), .B1(new_n483), .B2(new_n494), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n293), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(G475), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT20), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n486), .A2(KEYINPUT19), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT19), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n343), .A2(new_n344), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n503), .A2(new_n200), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT91), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n508), .A2(new_n348), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n479), .A2(new_n480), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT90), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n479), .A2(new_n480), .A3(KEYINPUT90), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n506), .A2(new_n507), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n509), .A2(new_n512), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n497), .B1(new_n494), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n483), .A2(new_n494), .A3(new_n497), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(G475), .A2(G902), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n502), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n502), .B(new_n520), .C1(new_n498), .C2(new_n516), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n501), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT94), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n520), .B1(new_n498), .B2(new_n516), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT20), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n522), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT94), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n528), .A2(new_n529), .A3(new_n501), .ZN(new_n530));
  XNOR2_X1  g344(.A(G116), .B(G122), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n531), .B(new_n393), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n238), .A2(G143), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT13), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n226), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n202), .A2(G128), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n533), .ZN(new_n537));
  OR2_X1    g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n535), .A2(new_n537), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n532), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  OR2_X1    g354(.A1(new_n192), .A2(G122), .ZN(new_n541));
  AND2_X1   g355(.A1(KEYINPUT14), .A2(G107), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n532), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n537), .B(G134), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n531), .A2(new_n542), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n540), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT9), .B(G234), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n549), .A2(new_n364), .A3(G953), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n540), .B(new_n550), .C1(new_n544), .C2(new_n547), .ZN(new_n553));
  AOI21_X1  g367(.A(G902), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(G478), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n555), .A2(KEYINPUT15), .ZN(new_n556));
  XOR2_X1   g370(.A(new_n554), .B(new_n556), .Z(new_n557));
  INV_X1    g371(.A(G952), .ZN(new_n558));
  AOI211_X1 g372(.A(G953), .B(new_n558), .C1(G234), .C2(G237), .ZN(new_n559));
  XOR2_X1   g373(.A(KEYINPUT21), .B(G898), .Z(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  AOI211_X1 g375(.A(new_n293), .B(new_n254), .C1(G234), .C2(G237), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n559), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n557), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n525), .A2(new_n530), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(G469), .A2(G902), .ZN(new_n566));
  INV_X1    g380(.A(G469), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n237), .B1(new_n239), .B2(new_n207), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n407), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT10), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n232), .A2(new_n233), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n432), .A2(new_n216), .A3(new_n427), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n407), .A2(KEYINPUT10), .A3(new_n240), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n571), .A2(new_n572), .A3(new_n573), .A4(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(G110), .B(G140), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n254), .A2(G227), .ZN(new_n577));
  XOR2_X1   g391(.A(new_n576), .B(new_n577), .Z(new_n578));
  NAND2_X1  g392(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n569), .B1(new_n240), .B2(new_n407), .ZN(new_n580));
  INV_X1    g394(.A(new_n572), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(KEYINPUT12), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n580), .A2(new_n581), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT12), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n579), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n571), .A2(new_n574), .A3(new_n573), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n581), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n578), .B1(new_n588), .B2(new_n575), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n567), .B(new_n293), .C1(new_n586), .C2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n585), .A2(new_n582), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n575), .ZN(new_n592));
  INV_X1    g406(.A(new_n578), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT82), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n579), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n575), .A2(KEYINPUT82), .A3(new_n578), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(new_n597), .A3(new_n588), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n566), .B(new_n590), .C1(new_n599), .C2(new_n567), .ZN(new_n600));
  INV_X1    g414(.A(G221), .ZN(new_n601));
  INV_X1    g415(.A(new_n549), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n601), .B1(new_n602), .B2(new_n293), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n565), .A2(new_n605), .ZN(new_n606));
  AND4_X1   g420(.A1(new_n319), .A2(new_n374), .A3(new_n470), .A4(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(new_n256), .ZN(G3));
  INV_X1    g422(.A(KEYINPUT95), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n609), .B1(new_n468), .B2(new_n375), .ZN(new_n610));
  INV_X1    g424(.A(new_n375), .ZN(new_n611));
  AOI211_X1 g425(.A(new_n611), .B(new_n438), .C1(new_n461), .C2(new_n462), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n466), .B1(new_n453), .B2(new_n609), .ZN(new_n614));
  OAI21_X1  g428(.A(KEYINPUT96), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n467), .B1(new_n612), .B2(KEYINPUT95), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT96), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n616), .B(new_n617), .C1(new_n612), .C2(new_n610), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n372), .A2(new_n373), .ZN(new_n620));
  OR3_X1    g434(.A1(new_n554), .A2(KEYINPUT98), .A3(G478), .ZN(new_n621));
  OAI21_X1  g435(.A(KEYINPUT98), .B1(new_n554), .B2(G478), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT97), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n548), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(KEYINPUT33), .ZN(new_n626));
  INV_X1    g440(.A(new_n552), .ZN(new_n627));
  INV_X1    g441(.A(new_n553), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n552), .A2(new_n625), .A3(KEYINPUT33), .A4(new_n553), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n629), .A2(G478), .A3(new_n293), .A4(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n623), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(KEYINPUT99), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT99), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n623), .A2(new_n631), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n528), .A2(new_n529), .A3(new_n501), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n529), .B1(new_n528), .B2(new_n501), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NOR4_X1   g453(.A1(new_n619), .A2(new_n620), .A3(new_n563), .A4(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(G902), .B1(new_n305), .B2(new_n310), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n641), .A2(new_n187), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n642), .A2(new_n605), .A3(new_n311), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT100), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT34), .B(G104), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G6));
  NAND2_X1  g461(.A1(new_n643), .A2(new_n374), .ZN(new_n648));
  INV_X1    g462(.A(new_n524), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n557), .ZN(new_n650));
  NOR4_X1   g464(.A1(new_n619), .A2(new_n648), .A3(new_n563), .A4(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT35), .B(G107), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  OR2_X1    g467(.A1(new_n358), .A2(KEYINPUT36), .ZN(new_n654));
  XOR2_X1   g468(.A(new_n354), .B(new_n654), .Z(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n370), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n367), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n642), .A2(new_n658), .A3(new_n311), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n470), .A2(new_n659), .A3(new_n606), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT37), .B(G110), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G12));
  INV_X1    g476(.A(KEYINPUT101), .ZN(new_n663));
  INV_X1    g477(.A(new_n605), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n319), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(G900), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n559), .B1(new_n562), .B2(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n650), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n615), .A2(new_n618), .A3(new_n657), .A4(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n663), .B1(new_n665), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n317), .A2(new_n313), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n311), .A2(KEYINPUT32), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n671), .A2(KEYINPUT72), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n312), .A2(new_n314), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n605), .B1(new_n675), .B2(new_n292), .ZN(new_n676));
  AND4_X1   g490(.A1(new_n618), .A2(new_n615), .A3(new_n657), .A4(new_n668), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n676), .A2(new_n677), .A3(KEYINPUT101), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n670), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G128), .ZN(G30));
  XNOR2_X1  g494(.A(new_n667), .B(KEYINPUT39), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n605), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n682), .A2(KEYINPUT40), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n682), .A2(KEYINPUT40), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n525), .A2(new_n530), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n685), .A2(new_n557), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n466), .A3(new_n658), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n683), .A2(new_n684), .A3(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n288), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n689), .A2(new_n260), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n293), .B1(new_n251), .B2(new_n259), .ZN(new_n691));
  OAI21_X1  g505(.A(G472), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n675), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n463), .A2(new_n439), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n611), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n695), .A2(KEYINPUT88), .A3(new_n453), .ZN(new_n696));
  INV_X1    g510(.A(new_n469), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(KEYINPUT38), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n688), .A2(new_n693), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G143), .ZN(G45));
  INV_X1    g516(.A(new_n667), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n685), .A2(new_n636), .A3(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n705), .A2(new_n615), .A3(new_n618), .A4(new_n657), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n665), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(new_n200), .ZN(G48));
  AOI21_X1  g522(.A(new_n291), .B1(new_n673), .B2(new_n674), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n586), .A2(new_n589), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n293), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(G469), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n590), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n603), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n709), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n640), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT41), .B(G113), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G15));
  INV_X1    g533(.A(new_n563), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n649), .A2(new_n720), .A3(new_n557), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n619), .A2(new_n715), .A3(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n709), .A2(new_n620), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G116), .ZN(G18));
  NOR3_X1   g539(.A1(new_n619), .A2(new_n565), .A3(new_n658), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n716), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G119), .ZN(G21));
  NAND3_X1  g542(.A1(new_n615), .A2(new_n618), .A3(new_n686), .ZN(new_n729));
  INV_X1    g543(.A(new_n641), .ZN(new_n730));
  XNOR2_X1  g544(.A(KEYINPUT103), .B(G472), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n300), .B(new_n302), .C1(new_n252), .C2(new_n259), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n297), .B(KEYINPUT102), .ZN(new_n733));
  AOI22_X1  g547(.A1(new_n730), .A2(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n367), .A2(new_n371), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n734), .A2(new_n714), .A3(new_n735), .A4(new_n720), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n729), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  NAND2_X1  g552(.A1(new_n732), .A2(new_n733), .ZN(new_n739));
  INV_X1    g553(.A(new_n731), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n657), .B(new_n739), .C1(new_n641), .C2(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n704), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n742), .A2(new_n618), .A3(new_n615), .A4(new_n714), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G125), .ZN(G27));
  AOI21_X1  g558(.A(new_n467), .B1(new_n696), .B2(new_n697), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n709), .A2(new_n620), .A3(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT104), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n747), .A2(new_n748), .A3(new_n664), .A4(new_n705), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n319), .A2(new_n745), .A3(new_n374), .A4(new_n664), .ZN(new_n750));
  OAI21_X1  g564(.A(KEYINPUT104), .B1(new_n750), .B2(new_n704), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT42), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n749), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT105), .ZN(new_n754));
  AOI211_X1 g568(.A(new_n291), .B(new_n314), .C1(new_n671), .C2(new_n754), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n755), .B1(new_n754), .B2(new_n671), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n756), .A2(new_n735), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n746), .A2(new_n704), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n757), .A2(KEYINPUT42), .A3(new_n664), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n753), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G131), .ZN(G33));
  NAND4_X1  g575(.A1(new_n723), .A2(new_n664), .A3(new_n668), .A4(new_n745), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G134), .ZN(G36));
  INV_X1    g577(.A(new_n599), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n764), .A2(KEYINPUT45), .ZN(new_n765));
  OAI21_X1  g579(.A(G469), .B1(new_n764), .B2(KEYINPUT45), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n767), .A2(KEYINPUT46), .A3(new_n566), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT46), .B1(new_n767), .B2(new_n566), .ZN(new_n769));
  INV_X1    g583(.A(new_n590), .ZN(new_n770));
  OR3_X1    g584(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n604), .ZN(new_n772));
  OR3_X1    g586(.A1(new_n772), .A2(KEYINPUT106), .A3(new_n681), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT106), .B1(new_n772), .B2(new_n681), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n637), .A2(new_n638), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT107), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n636), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT43), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n776), .B(new_n636), .C1(KEYINPUT107), .C2(KEYINPUT43), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n782), .B(new_n657), .C1(new_n311), .C2(new_n642), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT44), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n746), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n775), .B(new_n785), .C1(new_n784), .C2(new_n783), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G137), .ZN(G39));
  INV_X1    g601(.A(KEYINPUT47), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n771), .A2(new_n788), .A3(new_n604), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n788), .B1(new_n771), .B2(new_n604), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR4_X1   g606(.A1(new_n319), .A2(new_n746), .A3(new_n374), .A4(new_n704), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT108), .ZN(new_n795));
  XOR2_X1   g609(.A(KEYINPUT109), .B(G140), .Z(new_n796));
  XNOR2_X1  g610(.A(new_n795), .B(new_n796), .ZN(G42));
  NAND3_X1  g611(.A1(new_n735), .A2(new_n466), .A3(new_n604), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n798), .B1(KEYINPUT49), .B2(new_n713), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n799), .B1(KEYINPUT49), .B2(new_n713), .ZN(new_n800));
  OR4_X1    g614(.A1(new_n693), .A2(new_n700), .A3(new_n778), .A4(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT51), .ZN(new_n802));
  OAI22_X1  g616(.A1(new_n790), .A2(new_n791), .B1(new_n604), .B2(new_n713), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n782), .A2(new_n559), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n734), .A2(new_n735), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n806), .A2(new_n807), .A3(new_n746), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(new_n803), .B2(new_n804), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n802), .B1(new_n805), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n700), .A2(new_n466), .ZN(new_n812));
  INV_X1    g626(.A(new_n806), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n807), .A2(new_n715), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n812), .A2(new_n813), .A3(KEYINPUT50), .A4(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT116), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n815), .A2(new_n816), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT114), .ZN(new_n819));
  INV_X1    g633(.A(new_n812), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n813), .A2(new_n814), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  XOR2_X1   g636(.A(KEYINPUT115), .B(KEYINPUT50), .Z(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n820), .A2(new_n821), .A3(new_n819), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n817), .B(new_n818), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n745), .A2(new_n714), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n806), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(new_n741), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n374), .A2(new_n559), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n693), .A2(new_n827), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n685), .A2(new_n636), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n831), .A2(KEYINPUT117), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT117), .B1(new_n831), .B2(new_n832), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n829), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n811), .A2(new_n826), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n803), .A2(new_n808), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n826), .A2(new_n837), .A3(new_n835), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(new_n802), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n831), .A2(new_n685), .A3(new_n636), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n558), .A2(G953), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n840), .B(new_n841), .C1(new_n821), .C2(new_n619), .ZN(new_n842));
  INV_X1    g656(.A(new_n757), .ZN(new_n843));
  OR3_X1    g657(.A1(new_n843), .A2(new_n828), .A3(KEYINPUT48), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT48), .B1(new_n843), .B2(new_n828), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n842), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n836), .A2(new_n839), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n743), .B1(new_n665), .B2(new_n706), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n848), .B1(new_n670), .B2(new_n678), .ZN(new_n849));
  INV_X1    g663(.A(new_n729), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n605), .A2(new_n657), .A3(new_n667), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n850), .A2(new_n693), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT52), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n848), .ZN(new_n854));
  AND4_X1   g668(.A1(KEYINPUT52), .A2(new_n679), .A3(new_n854), .A4(new_n852), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n640), .A2(new_n716), .B1(new_n722), .B2(new_n723), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n525), .A2(new_n530), .A3(new_n557), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n563), .B1(new_n639), .B2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n643), .A2(new_n859), .A3(new_n470), .A4(new_n374), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n860), .B(new_n660), .C1(new_n729), .C2(new_n736), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n861), .A2(new_n607), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n857), .A2(new_n862), .A3(new_n727), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n524), .A2(new_n557), .A3(new_n667), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n864), .B(new_n466), .C1(new_n465), .C2(new_n469), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT110), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n658), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n698), .A2(KEYINPUT110), .A3(new_n466), .A4(new_n864), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n867), .A2(new_n319), .A3(new_n664), .A4(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n741), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n705), .A2(new_n745), .A3(new_n664), .A4(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n668), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n869), .B(new_n871), .C1(new_n750), .C2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT111), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n762), .A2(KEYINPUT111), .A3(new_n871), .A4(new_n869), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n760), .A2(new_n863), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT53), .B1(new_n856), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n679), .A2(new_n854), .A3(new_n852), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT52), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n849), .A2(KEYINPUT52), .A3(new_n852), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n857), .A2(new_n862), .A3(new_n727), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n885), .B1(new_n875), .B2(new_n876), .ZN(new_n886));
  XOR2_X1   g700(.A(KEYINPUT112), .B(KEYINPUT53), .Z(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n884), .A2(new_n886), .A3(new_n760), .A4(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n879), .A2(KEYINPUT54), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n888), .B1(new_n856), .B2(new_n878), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n884), .A2(new_n886), .A3(KEYINPUT53), .A4(new_n760), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(KEYINPUT113), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT113), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n890), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n847), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(G952), .A2(G953), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n801), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT119), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT119), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n903), .B(new_n801), .C1(new_n899), .C2(new_n900), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n902), .A2(new_n904), .ZN(G75));
  NOR2_X1   g719(.A1(new_n254), .A2(G952), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n891), .A2(new_n893), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(G902), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT56), .B1(new_n910), .B2(G210), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n447), .B(KEYINPUT120), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT55), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(new_n448), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n907), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n909), .B(KEYINPUT121), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n611), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT56), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n914), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n915), .B1(new_n917), .B2(new_n919), .ZN(G51));
  INV_X1    g734(.A(new_n767), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n566), .B(KEYINPUT57), .Z(new_n922));
  INV_X1    g736(.A(new_n894), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n892), .B1(new_n891), .B2(new_n893), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n710), .ZN(new_n926));
  AOI22_X1  g740(.A1(new_n921), .A2(new_n916), .B1(new_n926), .B2(KEYINPUT122), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n926), .A2(KEYINPUT122), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n906), .B1(new_n927), .B2(new_n928), .ZN(G54));
  NOR2_X1   g743(.A1(new_n909), .A2(KEYINPUT121), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT121), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n931), .B1(new_n908), .B2(G902), .ZN(new_n932));
  OAI211_X1 g746(.A(KEYINPUT58), .B(G475), .C1(new_n930), .C2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n933), .A2(new_n518), .A3(new_n517), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n916), .A2(KEYINPUT58), .A3(G475), .A4(new_n519), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n934), .A2(new_n935), .A3(new_n907), .ZN(G60));
  NOR2_X1   g750(.A1(new_n923), .A2(new_n924), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n629), .A2(new_n630), .ZN(new_n938));
  NAND2_X1  g752(.A1(G478), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT59), .Z(new_n940));
  NOR3_X1   g754(.A1(new_n937), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n940), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n896), .A2(new_n898), .A3(new_n942), .ZN(new_n943));
  AOI211_X1 g757(.A(new_n906), .B(new_n941), .C1(new_n938), .C2(new_n943), .ZN(G63));
  NAND2_X1  g758(.A1(G217), .A2(G902), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT60), .Z(new_n946));
  NAND3_X1  g760(.A1(new_n908), .A2(new_n655), .A3(new_n946), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n908), .A2(new_n946), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n907), .B(new_n947), .C1(new_n948), .C2(new_n369), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n949), .B1(KEYINPUT123), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(KEYINPUT123), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT124), .Z(new_n953));
  XNOR2_X1  g767(.A(new_n951), .B(new_n953), .ZN(G66));
  INV_X1    g768(.A(G224), .ZN(new_n955));
  OAI21_X1  g769(.A(G953), .B1(new_n561), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n956), .B1(new_n863), .B2(G953), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT125), .Z(new_n958));
  INV_X1    g772(.A(G898), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n912), .B1(new_n959), .B2(G953), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n958), .B(new_n960), .ZN(G69));
  NAND2_X1  g775(.A1(new_n285), .A2(new_n286), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT126), .Z(new_n963));
  NAND2_X1  g777(.A1(new_n503), .A2(new_n505), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n963), .B(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n795), .A2(new_n786), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT127), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT62), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n849), .B(new_n701), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n968), .A2(new_n969), .ZN(new_n971));
  OR2_X1    g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n970), .A2(new_n971), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n682), .B1(new_n639), .B2(new_n858), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n747), .A2(new_n974), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n967), .A2(new_n972), .A3(new_n973), .A4(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n966), .B1(new_n976), .B2(new_n254), .ZN(new_n977));
  INV_X1    g791(.A(new_n762), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n843), .A2(new_n729), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n978), .B1(new_n775), .B2(new_n979), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n795), .A2(new_n786), .A3(new_n980), .A4(new_n849), .ZN(new_n981));
  INV_X1    g795(.A(new_n760), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n254), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n254), .A2(G900), .ZN(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n965), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n254), .B1(G227), .B2(G900), .ZN(new_n987));
  OR3_X1    g801(.A1(new_n977), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n987), .B1(new_n977), .B2(new_n986), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(G72));
  NAND2_X1  g804(.A1(G472), .A2(G902), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT63), .Z(new_n992));
  OAI21_X1  g806(.A(new_n992), .B1(new_n976), .B2(new_n885), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n906), .B1(new_n993), .B2(new_n690), .ZN(new_n994));
  INV_X1    g808(.A(new_n992), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n995), .B1(new_n289), .B2(new_n299), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n879), .A2(new_n889), .A3(new_n996), .ZN(new_n997));
  NOR3_X1   g811(.A1(new_n981), .A2(new_n982), .A3(new_n885), .ZN(new_n998));
  OAI211_X1 g812(.A(new_n260), .B(new_n689), .C1(new_n998), .C2(new_n995), .ZN(new_n999));
  AND3_X1   g813(.A1(new_n994), .A2(new_n997), .A3(new_n999), .ZN(G57));
endmodule


