//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 0 0 0 1 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 1 1 1 0 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G250), .ZN(new_n205));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(G13), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  INV_X1    g0011(.A(G264), .ZN(new_n212));
  AOI211_X1 g0012(.A(new_n205), .B(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT64), .B(G244), .ZN(new_n215));
  AOI22_X1  g0015(.A1(new_n215), .A2(G77), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G50), .ZN(new_n217));
  INV_X1    g0017(.A(G226), .ZN(new_n218));
  INV_X1    g0018(.A(G107), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n212), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n221), .A2(new_n205), .ZN(new_n222));
  INV_X1    g0022(.A(G58), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G68), .ZN(new_n226));
  INV_X1    g0026(.A(G238), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NOR4_X1   g0028(.A1(new_n220), .A2(new_n222), .A3(new_n225), .A4(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G97), .A2(G257), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n208), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT1), .Z(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n233), .A2(new_n207), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n202), .A2(G50), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  AOI211_X1 g0036(.A(new_n214), .B(new_n232), .C1(new_n234), .C2(new_n236), .ZN(G361));
  XOR2_X1   g0037(.A(G250), .B(G257), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT66), .B(G264), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n242));
  XNOR2_X1  g0042(.A(G238), .B(G244), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G226), .B(G232), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n241), .B(new_n246), .ZN(G358));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT67), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G68), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n251), .B(new_n254), .Z(G351));
  AOI21_X1  g0055(.A(new_n207), .B1(new_n201), .B2(new_n217), .ZN(new_n256));
  XOR2_X1   g0056(.A(new_n256), .B(KEYINPUT70), .Z(new_n257));
  NAND2_X1  g0057(.A1(new_n207), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT69), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XOR2_X1   g0060(.A(KEYINPUT8), .B(G58), .Z(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n260), .A2(new_n261), .B1(G150), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n265), .A2(new_n233), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n206), .A2(G20), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(new_n209), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n217), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n266), .A2(G50), .A3(new_n269), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n268), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  AND2_X1   g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(G1698), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G222), .ZN(new_n278));
  INV_X1    g0078(.A(G77), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT3), .ZN(new_n280));
  INV_X1    g0080(.A(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G1698), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT68), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n284), .A2(KEYINPUT68), .A3(G1698), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G223), .ZN(new_n290));
  OAI221_X1 g0090(.A(new_n278), .B1(new_n279), .B2(new_n284), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n233), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G41), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n297));
  INV_X1    g0097(.A(G274), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n294), .A2(new_n297), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n296), .B(new_n300), .C1(new_n218), .C2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G179), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n303), .A2(KEYINPUT71), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(KEYINPUT71), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n273), .B1(new_n302), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n301), .A2(new_n218), .ZN(new_n309));
  AOI211_X1 g0109(.A(new_n309), .B(new_n299), .C1(new_n291), .C2(new_n295), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n310), .A2(G169), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT9), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n273), .A2(new_n313), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n268), .A2(KEYINPUT9), .A3(new_n271), .A4(new_n272), .ZN(new_n315));
  INV_X1    g0115(.A(G200), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n314), .B(new_n315), .C1(new_n310), .C2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G190), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n302), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(KEYINPUT10), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n314), .A2(new_n315), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n302), .A2(G200), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT10), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n310), .A2(G190), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n321), .A2(new_n322), .A3(new_n323), .A4(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n312), .B1(new_n320), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G1698), .ZN(new_n327));
  OAI211_X1 g0127(.A(G226), .B(new_n327), .C1(new_n274), .C2(new_n275), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT74), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n284), .A2(KEYINPUT74), .A3(G226), .A4(new_n327), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n284), .A2(G232), .A3(G1698), .ZN(new_n332));
  NAND2_X1  g0132(.A1(G33), .A2(G97), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n330), .A2(new_n331), .A3(new_n332), .A4(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT75), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n328), .A2(new_n329), .B1(G33), .B2(G97), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT75), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n336), .A2(new_n337), .A3(new_n331), .A4(new_n332), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n335), .A2(new_n295), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT13), .ZN(new_n340));
  INV_X1    g0140(.A(new_n301), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT76), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT76), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n227), .B1(new_n301), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n299), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n339), .A2(new_n340), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n340), .B1(new_n339), .B2(new_n345), .ZN(new_n347));
  OAI21_X1  g0147(.A(G169), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT14), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n339), .A2(new_n345), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT13), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n339), .A2(new_n340), .A3(new_n345), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(G179), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT14), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n354), .B(G169), .C1(new_n346), .C2(new_n347), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n349), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n270), .ZN(new_n357));
  NOR3_X1   g0157(.A1(new_n357), .A2(KEYINPUT12), .A3(G68), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT12), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n359), .B1(new_n270), .B2(new_n226), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n266), .A2(new_n269), .ZN(new_n361));
  OAI22_X1  g0161(.A1(new_n358), .A2(new_n360), .B1(new_n226), .B2(new_n361), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n260), .A2(G77), .B1(G20), .B2(new_n226), .ZN(new_n363));
  INV_X1    g0163(.A(new_n262), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n363), .B1(new_n217), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n267), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT11), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT11), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n365), .A2(new_n368), .A3(new_n267), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n362), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n356), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(G200), .B1(new_n346), .B2(new_n347), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n351), .A2(G190), .A3(new_n352), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(new_n374), .A3(new_n370), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT77), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT77), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n373), .A2(new_n374), .A3(new_n377), .A4(new_n370), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n326), .A2(new_n372), .A3(new_n376), .A4(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n357), .A2(G77), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n261), .A2(new_n262), .B1(G20), .B2(G77), .ZN(new_n381));
  XNOR2_X1  g0181(.A(KEYINPUT15), .B(G87), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT73), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n382), .B(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n381), .B1(new_n385), .B2(new_n258), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n380), .B1(new_n386), .B2(new_n267), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(new_n279), .B2(new_n361), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n277), .A2(G232), .ZN(new_n389));
  XNOR2_X1  g0189(.A(KEYINPUT72), .B(G107), .ZN(new_n390));
  OAI221_X1 g0190(.A(new_n389), .B1(new_n284), .B2(new_n390), .C1(new_n289), .C2(new_n227), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n295), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n341), .A2(new_n215), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n392), .A2(new_n300), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n388), .B1(new_n394), .B2(G200), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n392), .A2(G190), .A3(new_n300), .A4(new_n393), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT16), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n282), .A2(new_n207), .A3(new_n283), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT7), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n282), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n283), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n226), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n223), .A2(new_n226), .ZN(new_n405));
  OAI21_X1  g0205(.A(G20), .B1(new_n405), .B2(new_n201), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n262), .A2(G159), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n399), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT7), .B1(new_n276), .B2(new_n207), .ZN(new_n410));
  INV_X1    g0210(.A(new_n403), .ZN(new_n411));
  OAI21_X1  g0211(.A(G68), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n408), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(KEYINPUT16), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n409), .A2(new_n414), .A3(new_n267), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT78), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT78), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n409), .A2(new_n414), .A3(new_n417), .A4(new_n267), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n300), .B1(new_n301), .B2(new_n224), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n290), .A2(new_n327), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n218), .A2(G1698), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n421), .B(new_n422), .C1(new_n274), .C2(new_n275), .ZN(new_n423));
  NAND2_X1  g0223(.A1(G33), .A2(G87), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n294), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n316), .B1(new_n420), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT79), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n423), .A2(new_n424), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n427), .B1(new_n428), .B2(new_n295), .ZN(new_n429));
  AOI211_X1 g0229(.A(KEYINPUT79), .B(new_n294), .C1(new_n423), .C2(new_n424), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n318), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n426), .B1(new_n431), .B2(new_n420), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n261), .A2(new_n270), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n433), .B1(new_n261), .B2(new_n361), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  AND4_X1   g0235(.A1(KEYINPUT17), .A2(new_n419), .A3(new_n432), .A4(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n434), .B1(new_n416), .B2(new_n418), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT17), .B1(new_n437), .B2(new_n432), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n419), .A2(new_n435), .ZN(new_n440));
  INV_X1    g0240(.A(new_n420), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n306), .B(new_n441), .C1(new_n429), .C2(new_n430), .ZN(new_n442));
  INV_X1    g0242(.A(G169), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n420), .B2(new_n425), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n442), .A2(KEYINPUT80), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT80), .B1(new_n442), .B2(new_n444), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n440), .A2(KEYINPUT18), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT18), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n442), .A2(new_n444), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT80), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n442), .A2(KEYINPUT80), .A3(new_n444), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n449), .B1(new_n437), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n448), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n392), .A2(new_n300), .A3(new_n306), .A4(new_n393), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n457), .A2(new_n388), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n394), .A2(new_n443), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n439), .A2(new_n456), .A3(new_n460), .ZN(new_n461));
  NOR3_X1   g0261(.A1(new_n379), .A2(new_n398), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT21), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n284), .A2(G257), .A3(new_n327), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n276), .A2(G303), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n465), .B(new_n466), .C1(new_n285), .C2(new_n212), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n295), .ZN(new_n468));
  XNOR2_X1  g0268(.A(KEYINPUT5), .B(G41), .ZN(new_n469));
  INV_X1    g0269(.A(G45), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(G1), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n469), .A2(G274), .A3(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n469), .A2(new_n471), .B1(new_n292), .B2(new_n293), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G270), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n468), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G169), .ZN(new_n476));
  OR2_X1    g0276(.A1(KEYINPUT84), .A2(G116), .ZN(new_n477));
  NAND2_X1  g0277(.A1(KEYINPUT84), .A2(G116), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n270), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n206), .A2(G33), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n357), .A2(new_n266), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(G116), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n266), .B1(G20), .B2(new_n479), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G283), .ZN(new_n486));
  INV_X1    g0286(.A(G97), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n486), .B(new_n207), .C1(G33), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT20), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n485), .A2(KEYINPUT20), .A3(new_n488), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n484), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n464), .B1(new_n476), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n491), .A2(new_n492), .ZN(new_n495));
  INV_X1    g0295(.A(new_n484), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n497), .A2(KEYINPUT21), .A3(G169), .A4(new_n475), .ZN(new_n498));
  AND2_X1   g0298(.A1(new_n468), .A2(new_n474), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n497), .A2(G179), .A3(new_n472), .A4(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n494), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n475), .A2(G200), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n503), .B(new_n493), .C1(new_n318), .C2(new_n475), .ZN(new_n504));
  AND2_X1   g0304(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(G41), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G41), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n471), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n294), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n472), .B1(new_n512), .B2(new_n211), .ZN(new_n513));
  OAI211_X1 g0313(.A(G244), .B(new_n327), .C1(new_n274), .C2(new_n275), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT4), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n284), .A2(KEYINPUT4), .A3(G244), .A4(new_n327), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n284), .A2(G250), .A3(G1698), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n516), .A2(new_n517), .A3(new_n486), .A4(new_n518), .ZN(new_n519));
  AOI211_X1 g0319(.A(new_n306), .B(new_n513), .C1(new_n295), .C2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n516), .A2(new_n517), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n518), .A2(new_n486), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n295), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n513), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n443), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n357), .A2(G97), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n482), .A2(new_n487), .ZN(new_n528));
  INV_X1    g0328(.A(new_n390), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n410), .B2(new_n411), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n487), .A2(new_n219), .A3(KEYINPUT6), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT6), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G97), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n219), .A2(KEYINPUT81), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT81), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G107), .ZN(new_n536));
  AND4_X1   g0336(.A1(new_n531), .A2(new_n533), .A3(new_n534), .A4(new_n536), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n531), .A2(new_n533), .B1(new_n534), .B2(new_n536), .ZN(new_n538));
  OAI21_X1  g0338(.A(G20), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n262), .A2(G77), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n530), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AOI211_X1 g0341(.A(new_n527), .B(new_n528), .C1(new_n541), .C2(new_n267), .ZN(new_n542));
  OAI21_X1  g0342(.A(KEYINPUT83), .B1(new_n526), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n523), .A2(new_n307), .A3(new_n524), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n513), .B1(new_n519), .B2(new_n295), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n544), .B1(new_n443), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n541), .A2(new_n267), .ZN(new_n547));
  INV_X1    g0347(.A(new_n527), .ZN(new_n548));
  INV_X1    g0348(.A(new_n528), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT83), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n546), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n543), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n482), .A2(new_n221), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n384), .A2(new_n357), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n284), .A2(new_n207), .A3(G68), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n258), .A2(new_n487), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n557), .A2(KEYINPUT19), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(G87), .A2(G97), .ZN(new_n560));
  AOI21_X1  g0360(.A(KEYINPUT85), .B1(new_n390), .B2(new_n560), .ZN(new_n561));
  AND2_X1   g0361(.A1(KEYINPUT72), .A2(G107), .ZN(new_n562));
  NOR2_X1   g0362(.A1(KEYINPUT72), .A2(G107), .ZN(new_n563));
  OAI211_X1 g0363(.A(KEYINPUT85), .B(new_n560), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n567), .A2(new_n207), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n556), .B(new_n559), .C1(new_n566), .C2(new_n568), .ZN(new_n569));
  AOI211_X1 g0369(.A(new_n554), .B(new_n555), .C1(new_n569), .C2(new_n267), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n227), .A2(new_n327), .ZN(new_n571));
  INV_X1    g0371(.A(G244), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(G1698), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n571), .B(new_n573), .C1(new_n274), .C2(new_n275), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n477), .A2(G33), .A3(new_n478), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n294), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n471), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n577), .A2(new_n298), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n294), .A2(new_n577), .A3(G250), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n579), .A2(new_n318), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n580), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n576), .A2(new_n582), .A3(new_n578), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n581), .B1(new_n583), .B2(G200), .ZN(new_n584));
  INV_X1    g0384(.A(new_n482), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n384), .ZN(new_n586));
  INV_X1    g0386(.A(new_n555), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n567), .A2(new_n207), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n561), .B2(new_n565), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n589), .A2(new_n556), .A3(new_n559), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n586), .B(new_n587), .C1(new_n590), .C2(new_n266), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n583), .A2(new_n307), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(new_n443), .B2(new_n583), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n570), .A2(new_n584), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n545), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n595), .A2(KEYINPUT82), .A3(G200), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT82), .ZN(new_n597));
  AOI21_X1  g0397(.A(G190), .B1(new_n597), .B2(G200), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n596), .B(new_n542), .C1(new_n595), .C2(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n482), .A2(new_n219), .ZN(new_n600));
  NOR3_X1   g0400(.A1(new_n207), .A2(KEYINPUT23), .A3(G107), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT23), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n575), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n601), .B1(new_n603), .B2(new_n207), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n207), .B(G87), .C1(new_n274), .C2(new_n275), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT22), .ZN(new_n606));
  OR2_X1    g0406(.A1(new_n606), .A2(KEYINPUT86), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n284), .A2(new_n207), .A3(G87), .A4(new_n607), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n529), .A2(KEYINPUT23), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n604), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT24), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT24), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n604), .A2(new_n611), .A3(new_n615), .A4(new_n612), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n600), .B1(new_n617), .B2(new_n267), .ZN(new_n618));
  OAI211_X1 g0418(.A(G257), .B(G1698), .C1(new_n274), .C2(new_n275), .ZN(new_n619));
  OAI211_X1 g0419(.A(G250), .B(new_n327), .C1(new_n274), .C2(new_n275), .ZN(new_n620));
  NAND2_X1  g0420(.A1(G33), .A2(G294), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n295), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n473), .A2(G264), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(new_n472), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT87), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n622), .A2(new_n295), .B1(new_n473), .B2(G264), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n628), .A2(KEYINPUT87), .A3(new_n472), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n627), .A2(new_n318), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n625), .A2(new_n316), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n270), .A2(new_n219), .ZN(new_n633));
  XNOR2_X1  g0433(.A(new_n633), .B(KEYINPUT25), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n618), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n553), .A2(new_n594), .A3(new_n599), .A4(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n623), .A2(G179), .A3(new_n472), .A4(new_n624), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT88), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT88), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n628), .A2(new_n640), .A3(G179), .A4(new_n472), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n625), .A2(new_n626), .ZN(new_n643));
  AOI21_X1  g0443(.A(KEYINPUT87), .B1(new_n628), .B2(new_n472), .ZN(new_n644));
  OAI21_X1  g0444(.A(G169), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n618), .A2(new_n635), .B1(new_n642), .B2(new_n645), .ZN(new_n646));
  NOR4_X1   g0446(.A1(new_n463), .A2(new_n506), .A3(new_n637), .A4(new_n646), .ZN(G372));
  AOI211_X1 g0447(.A(new_n600), .B(new_n634), .C1(new_n617), .C2(new_n267), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n443), .B1(new_n627), .B2(new_n629), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n639), .A2(new_n641), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT89), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n648), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n617), .A2(new_n267), .ZN(new_n654));
  INV_X1    g0454(.A(new_n600), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(new_n655), .A3(new_n635), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n642), .A2(new_n645), .ZN(new_n657));
  AOI21_X1  g0457(.A(KEYINPUT89), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n637), .B1(new_n659), .B2(new_n502), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n594), .A2(new_n543), .A3(new_n552), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(KEYINPUT26), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n591), .A2(new_n593), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n526), .A2(new_n542), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n594), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n662), .A2(new_n663), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n462), .B1(new_n660), .B2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n312), .ZN(new_n669));
  INV_X1    g0469(.A(new_n460), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n371), .A2(new_n356), .B1(new_n670), .B2(new_n375), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n437), .A2(new_n432), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT17), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n437), .A2(KEYINPUT17), .A3(new_n432), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n456), .B1(new_n671), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n320), .A2(new_n325), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n668), .A2(new_n669), .A3(new_n679), .ZN(G369));
  XOR2_X1   g0480(.A(KEYINPUT90), .B(KEYINPUT27), .Z(new_n681));
  NOR3_X1   g0481(.A1(new_n209), .A2(G1), .A3(G20), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n682), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G213), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(G343), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(new_n493), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n501), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n506), .B2(new_n689), .ZN(new_n691));
  XNOR2_X1  g0491(.A(KEYINPUT91), .B(G330), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n656), .A2(new_n657), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n656), .A2(new_n687), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(new_n695), .A3(new_n636), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n696), .A2(KEYINPUT92), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(KEYINPUT92), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n694), .B2(new_n688), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n693), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n502), .A2(new_n687), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n697), .A2(new_n698), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT93), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n688), .B1(new_n653), .B2(new_n658), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n704), .B1(new_n703), .B2(new_n705), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n701), .B1(new_n706), .B2(new_n707), .ZN(G399));
  NAND2_X1  g0508(.A1(new_n566), .A2(new_n483), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n210), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n711), .A2(KEYINPUT94), .A3(new_n507), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT94), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n210), .B2(G41), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n710), .A2(G1), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n716), .B1(new_n235), .B2(new_n715), .ZN(new_n717));
  XOR2_X1   g0517(.A(KEYINPUT95), .B(KEYINPUT28), .Z(new_n718));
  XNOR2_X1  g0518(.A(new_n717), .B(new_n718), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n546), .A2(new_n551), .A3(new_n550), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n551), .B1(new_n546), .B2(new_n550), .ZN(new_n721));
  OAI211_X1 g0521(.A(new_n594), .B(new_n599), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n636), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n724), .A2(new_n505), .A3(new_n694), .A4(new_n688), .ZN(new_n725));
  INV_X1    g0525(.A(new_n638), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n499), .A2(new_n726), .A3(new_n583), .A4(new_n545), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT30), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n475), .A2(new_n595), .A3(new_n306), .A4(new_n625), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n729), .A2(new_n583), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n688), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n731), .A2(KEYINPUT31), .ZN(new_n732));
  XNOR2_X1  g0532(.A(KEYINPUT96), .B(KEYINPUT31), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n725), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n692), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n555), .B1(new_n569), .B2(new_n267), .ZN(new_n738));
  INV_X1    g0538(.A(new_n554), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n584), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n663), .A2(new_n740), .A3(new_n550), .A4(new_n546), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n663), .A2(KEYINPUT98), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT98), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n591), .A2(new_n593), .A3(new_n743), .ZN(new_n744));
  AOI22_X1  g0544(.A1(new_n741), .A2(KEYINPUT26), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n594), .A2(new_n543), .A3(new_n665), .A4(new_n552), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n636), .B1(new_n646), .B2(new_n501), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n745), .B(new_n746), .C1(new_n747), .C2(new_n722), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT99), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n748), .A2(new_n749), .A3(new_n688), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n749), .B1(new_n748), .B2(new_n688), .ZN(new_n751));
  OAI21_X1  g0551(.A(KEYINPUT29), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n688), .B1(new_n660), .B2(new_n667), .ZN(new_n753));
  XOR2_X1   g0553(.A(KEYINPUT97), .B(KEYINPUT29), .Z(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n737), .B1(new_n752), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n719), .B1(new_n756), .B2(G1), .ZN(G364));
  NOR2_X1   g0557(.A1(G13), .A2(G33), .ZN(new_n758));
  XOR2_X1   g0558(.A(new_n758), .B(KEYINPUT101), .Z(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(G20), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n233), .B1(G20), .B2(new_n443), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n711), .A2(new_n276), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n765), .B1(new_n251), .B2(G45), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n236), .A2(new_n470), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n766), .A2(new_n767), .B1(new_n483), .B2(new_n210), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n711), .A2(G355), .A3(new_n284), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n764), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n715), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n209), .A2(G20), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G45), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n773), .A2(KEYINPUT100), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(KEYINPUT100), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n774), .A2(G1), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n771), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n207), .A2(G190), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n779), .A2(new_n303), .A3(G200), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n780), .B(KEYINPUT102), .Z(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G179), .A2(G200), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n784), .B(KEYINPUT103), .Z(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n782), .A2(G283), .B1(new_n786), .B2(G329), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT104), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n207), .A2(new_n318), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G200), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(G179), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n207), .B1(new_n783), .B2(G190), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n791), .A2(G303), .B1(G294), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n307), .A2(G200), .A3(new_n779), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(KEYINPUT105), .B(KEYINPUT33), .ZN(new_n797));
  INV_X1    g0597(.A(G317), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n797), .B(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n284), .B1(new_n796), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n788), .A2(new_n794), .A3(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n307), .A2(new_n316), .A3(new_n789), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n801), .B1(G322), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(G311), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n307), .A2(new_n779), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(G200), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G326), .ZN(new_n809));
  INV_X1    g0609(.A(new_n790), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n307), .A2(new_n810), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n804), .B1(new_n805), .B2(new_n808), .C1(new_n809), .C2(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT106), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n284), .B1(new_n795), .B2(new_n226), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n808), .A2(new_n279), .B1(new_n811), .B2(new_n217), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n814), .B(new_n815), .C1(G58), .C2(new_n803), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n781), .A2(new_n219), .ZN(new_n817));
  INV_X1    g0617(.A(new_n784), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(G159), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT32), .ZN(new_n820));
  INV_X1    g0620(.A(new_n791), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(new_n221), .ZN(new_n822));
  NOR3_X1   g0622(.A1(new_n817), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n816), .B(new_n823), .C1(new_n487), .C2(new_n792), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n813), .A2(new_n824), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n770), .B(new_n778), .C1(new_n825), .C2(new_n762), .ZN(new_n826));
  INV_X1    g0626(.A(new_n761), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n826), .B1(new_n691), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n693), .A2(new_n777), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n692), .B2(new_n691), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n828), .A2(new_n830), .ZN(G396));
  AND4_X1   g0631(.A1(new_n388), .A2(new_n459), .A3(new_n457), .A4(new_n688), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n388), .A2(new_n687), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n397), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n832), .B1(new_n834), .B2(new_n460), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n753), .A2(new_n836), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n688), .B(new_n835), .C1(new_n660), .C2(new_n667), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n737), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT107), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n841), .B(new_n778), .C1(new_n737), .C2(new_n839), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n836), .A2(new_n759), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n276), .B1(new_n821), .B2(new_n219), .ZN(new_n844));
  INV_X1    g0644(.A(G294), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n808), .A2(new_n479), .B1(new_n845), .B2(new_n802), .ZN(new_n846));
  INV_X1    g0646(.A(new_n811), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n844), .B(new_n846), .C1(G303), .C2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(G283), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n785), .A2(new_n805), .B1(new_n849), .B2(new_n795), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(G97), .B2(new_n793), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n848), .B(new_n851), .C1(new_n221), .C2(new_n781), .ZN(new_n852));
  AOI22_X1  g0652(.A1(G159), .A2(new_n807), .B1(new_n803), .B2(G143), .ZN(new_n853));
  INV_X1    g0653(.A(G137), .ZN(new_n854));
  INV_X1    g0654(.A(G150), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n853), .B1(new_n854), .B2(new_n811), .C1(new_n855), .C2(new_n795), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT34), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n786), .A2(G132), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n782), .A2(G68), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n276), .B1(new_n791), .B2(G50), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n857), .A2(new_n858), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n792), .A2(new_n223), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n852), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n762), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n762), .A2(new_n758), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n279), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n843), .A2(new_n777), .A3(new_n864), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n842), .A2(new_n867), .ZN(G384));
  INV_X1    g0668(.A(new_n685), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n415), .A2(new_n435), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n448), .A2(new_n455), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n869), .B(new_n870), .C1(new_n871), .C2(new_n676), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n440), .A2(new_n869), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n437), .A2(new_n454), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT110), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n873), .B(new_n672), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  XOR2_X1   g0676(.A(KEYINPUT111), .B(KEYINPUT37), .Z(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n440), .A2(new_n447), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n878), .B1(new_n879), .B2(KEYINPUT110), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n870), .B1(new_n447), .B2(new_n869), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n881), .A2(new_n672), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT37), .ZN(new_n883));
  OAI22_X1  g0683(.A1(new_n876), .A2(new_n880), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n872), .A2(KEYINPUT38), .A3(new_n884), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n879), .A2(new_n873), .A3(new_n672), .ZN(new_n886));
  OAI22_X1  g0686(.A1(new_n886), .A2(new_n878), .B1(new_n876), .B2(new_n880), .ZN(new_n887));
  INV_X1    g0687(.A(new_n873), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n871), .B2(new_n676), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT38), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(KEYINPUT40), .B1(new_n885), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n376), .A2(new_n378), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n371), .B(new_n687), .C1(new_n892), .C2(new_n356), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n371), .A2(KEYINPUT109), .A3(new_n687), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT109), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(new_n370), .B2(new_n688), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n372), .A2(new_n375), .A3(new_n894), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  OR2_X1    g0698(.A1(new_n731), .A2(new_n733), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n731), .A2(KEYINPUT31), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n725), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n898), .A2(new_n835), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n891), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT40), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT38), .B1(new_n872), .B2(new_n884), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n885), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n904), .B1(new_n906), .B2(new_n902), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT114), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(KEYINPUT114), .B(new_n904), .C1(new_n906), .C2(new_n902), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n903), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n462), .A2(new_n901), .ZN(new_n912));
  XOR2_X1   g0712(.A(new_n911), .B(new_n912), .Z(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n692), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT39), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n885), .B2(new_n890), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n356), .A2(new_n371), .A3(new_n688), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT38), .ZN(new_n919));
  INV_X1    g0719(.A(new_n870), .ZN(new_n920));
  AOI211_X1 g0720(.A(new_n685), .B(new_n920), .C1(new_n439), .C2(new_n456), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n883), .B1(new_n881), .B2(new_n672), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n672), .B1(new_n437), .B2(new_n685), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n875), .B1(new_n440), .B2(new_n447), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n877), .B1(new_n874), .B2(new_n875), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n922), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n919), .B1(new_n921), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n872), .A2(new_n884), .A3(KEYINPUT38), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n928), .A2(KEYINPUT39), .A3(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n916), .A2(new_n918), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n456), .A2(new_n869), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n832), .B(KEYINPUT108), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n838), .A2(new_n933), .B1(new_n893), .B2(new_n897), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n928), .A2(new_n929), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT112), .ZN(new_n937));
  AND3_X1   g0737(.A1(new_n931), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n937), .B1(new_n931), .B2(new_n936), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n914), .B(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n679), .A2(new_n669), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n752), .A2(new_n462), .A3(new_n755), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT113), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n752), .A2(new_n462), .A3(KEYINPUT113), .A4(new_n755), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n942), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n941), .B(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n206), .B2(new_n772), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n537), .A2(new_n538), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n483), .B1(new_n950), .B2(KEYINPUT35), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n951), .B(new_n234), .C1(KEYINPUT35), .C2(new_n950), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT36), .ZN(new_n953));
  OAI21_X1  g0753(.A(G77), .B1(new_n223), .B2(new_n226), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n235), .A2(new_n954), .B1(G50), .B2(new_n226), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n955), .A2(G1), .A3(new_n209), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n949), .A2(new_n953), .A3(new_n956), .ZN(G367));
  INV_X1    g0757(.A(new_n241), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n763), .B1(new_n958), .B2(new_n765), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(new_n210), .B2(new_n384), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT46), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n821), .B2(new_n479), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n962), .B1(new_n845), .B2(new_n795), .C1(new_n808), .C2(new_n849), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n791), .A2(KEYINPUT46), .A3(G116), .ZN(new_n964));
  INV_X1    g0764(.A(G303), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n964), .B1(new_n487), .B2(new_n780), .C1(new_n802), .C2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n284), .B1(new_n793), .B2(new_n529), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n967), .B(new_n968), .C1(new_n798), .C2(new_n784), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n963), .B(new_n969), .C1(G311), .C2(new_n847), .ZN(new_n970));
  INV_X1    g0770(.A(new_n780), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(G77), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n847), .A2(G143), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n973), .B1(new_n855), .B2(new_n802), .C1(new_n808), .C2(new_n217), .ZN(new_n974));
  INV_X1    g0774(.A(G159), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n795), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n792), .A2(new_n226), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n284), .B1(new_n854), .B2(new_n784), .C1(new_n821), .C2(new_n223), .ZN(new_n978));
  NOR4_X1   g0778(.A1(new_n974), .A2(new_n976), .A3(new_n977), .A4(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n970), .B1(new_n972), .B2(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT47), .Z(new_n981));
  AOI211_X1 g0781(.A(new_n778), .B(new_n960), .C1(new_n981), .C2(new_n762), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n594), .B1(new_n570), .B2(new_n688), .ZN(new_n983));
  OR3_X1    g0783(.A1(new_n663), .A2(new_n570), .A3(new_n688), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n761), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n982), .A2(new_n987), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n553), .B(new_n599), .C1(new_n542), .C2(new_n688), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n664), .A2(new_n687), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n703), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(KEYINPUT42), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n993), .A2(KEYINPUT42), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n553), .B1(new_n992), .B2(new_n694), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n994), .A2(new_n995), .B1(new_n688), .B2(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n985), .B(KEYINPUT115), .Z(new_n998));
  INV_X1    g0798(.A(KEYINPUT43), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n997), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n999), .B2(new_n986), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n997), .A2(new_n1001), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n701), .A2(new_n992), .ZN(new_n1005));
  AND3_X1   g0805(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1005), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n991), .B1(new_n706), .B2(new_n707), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT45), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OAI211_X1 g0812(.A(KEYINPUT45), .B(new_n991), .C1(new_n706), .C2(new_n707), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n703), .A2(new_n705), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(KEYINPUT93), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1016), .A2(new_n1017), .A3(new_n992), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT44), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1016), .A2(KEYINPUT44), .A3(new_n1017), .A4(new_n992), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1014), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n701), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n703), .B1(new_n700), .B2(new_n702), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(new_n693), .Z(new_n1027));
  INV_X1    g0827(.A(new_n756), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1014), .A2(new_n1022), .A3(new_n701), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1025), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n756), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n715), .B(KEYINPUT41), .Z(new_n1033));
  AOI21_X1  g0833(.A(new_n776), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n988), .B1(new_n1009), .B2(new_n1034), .ZN(G387));
  AOI21_X1  g0835(.A(new_n709), .B1(G68), .B2(G77), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n261), .A2(new_n217), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT50), .Z(new_n1038));
  NAND3_X1  g0838(.A1(new_n1036), .A2(new_n470), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n765), .B1(new_n246), .B2(G45), .ZN(new_n1040));
  NOR3_X1   g0840(.A1(new_n710), .A2(new_n210), .A3(new_n276), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1039), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n210), .A2(new_n219), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n764), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n821), .A2(new_n279), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n385), .A2(new_n792), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(G159), .B2(new_n847), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n226), .B2(new_n808), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1045), .B(new_n1048), .C1(new_n261), .C2(new_n796), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n782), .A2(G97), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n803), .A2(G50), .B1(G150), .B2(new_n818), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1049), .A2(new_n284), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(G322), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n795), .A2(new_n805), .B1(new_n811), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G303), .B2(new_n807), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n798), .B2(new_n802), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT48), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(new_n849), .B2(new_n792), .C1(new_n845), .C2(new_n821), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT49), .Z(new_n1059));
  OAI221_X1 g0859(.A(new_n276), .B1(new_n784), .B2(new_n809), .C1(new_n479), .C2(new_n780), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1052), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1044), .B1(new_n1061), .B2(new_n762), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1062), .B(new_n777), .C1(new_n700), .C2(new_n827), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n776), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n771), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1063), .B1(new_n1064), .B2(new_n1027), .C1(new_n1066), .C2(new_n1029), .ZN(G393));
  NAND3_X1  g0867(.A1(new_n1025), .A2(KEYINPUT116), .A3(new_n1030), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1030), .A2(KEYINPUT116), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n771), .B(new_n1031), .C1(new_n1070), .C2(new_n1029), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n763), .B1(new_n487), .B2(new_n711), .C1(new_n254), .C2(new_n765), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n777), .B(new_n1072), .C1(new_n991), .C2(new_n827), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n791), .A2(G68), .B1(G143), .B2(new_n818), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT117), .Z(new_n1075));
  NAND2_X1  g0875(.A1(new_n793), .A2(G77), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n261), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1076), .B1(new_n808), .B2(new_n1077), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n1075), .A2(new_n1078), .A3(new_n276), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n796), .A2(G50), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n802), .A2(new_n975), .B1(new_n811), .B2(new_n855), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT51), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n1082), .A2(new_n1081), .B1(new_n782), .B2(G87), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1079), .A2(new_n1080), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n802), .A2(new_n805), .B1(new_n811), .B2(new_n798), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT52), .Z(new_n1087));
  OAI21_X1  g0887(.A(new_n276), .B1(new_n795), .B2(new_n965), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n818), .A2(G322), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1089), .B1(new_n479), .B2(new_n792), .C1(new_n821), .C2(new_n849), .ZN(new_n1090));
  OR4_X1    g0890(.A1(new_n817), .A2(new_n1087), .A3(new_n1088), .A4(new_n1090), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n808), .A2(new_n845), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1085), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1073), .B1(new_n762), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(new_n1070), .B2(new_n776), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1071), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT118), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1071), .A2(KEYINPUT118), .A3(new_n1095), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(G390));
  NAND2_X1  g0900(.A1(new_n916), .A2(new_n930), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n838), .A2(new_n933), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n898), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n917), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n748), .A2(new_n688), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(KEYINPUT99), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n748), .A2(new_n749), .A3(new_n688), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n836), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n933), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n898), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n890), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n918), .B1(new_n1111), .B2(new_n929), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1101), .A2(new_n1104), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n898), .A2(G330), .A3(new_n835), .A4(new_n901), .ZN(new_n1114));
  OAI21_X1  g0914(.A(KEYINPUT119), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n898), .A2(new_n692), .A3(new_n735), .A4(new_n835), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT119), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1114), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n916), .A2(new_n930), .B1(new_n1103), .B2(new_n917), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n917), .B1(new_n885), .B2(new_n890), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n835), .B1(new_n750), .B2(new_n751), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n933), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1121), .B1(new_n1123), .B2(new_n898), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1118), .B(new_n1119), .C1(new_n1120), .C2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1115), .A2(new_n1117), .A3(new_n1125), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n462), .A2(G330), .A3(new_n901), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n942), .B(new_n1127), .C1(new_n945), .C2(new_n946), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n735), .A2(new_n692), .A3(new_n835), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n893), .A2(new_n897), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n1114), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n1102), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n901), .A2(G330), .A3(new_n835), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n1130), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1135), .A2(new_n933), .A3(new_n1116), .A4(new_n1122), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(KEYINPUT120), .B1(new_n1128), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1127), .ZN(new_n1139));
  AND4_X1   g0939(.A1(KEYINPUT120), .A2(new_n1137), .A3(new_n947), .A4(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1126), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n947), .A2(new_n1139), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1137), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1144), .A2(new_n1117), .A3(new_n1125), .A4(new_n1115), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1141), .A2(new_n771), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1101), .A2(new_n759), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n865), .A2(new_n1077), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n1076), .B1(new_n390), .B2(new_n795), .C1(new_n808), .C2(new_n487), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n822), .B(new_n1150), .C1(G116), .C2(new_n803), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n284), .B1(new_n786), .B2(G294), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n847), .A2(G283), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1151), .A2(new_n859), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n795), .A2(new_n854), .B1(new_n975), .B2(new_n792), .ZN(new_n1155));
  XOR2_X1   g0955(.A(KEYINPUT54), .B(G143), .Z(new_n1156));
  AOI21_X1  g0956(.A(new_n1155), .B1(new_n807), .B2(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT121), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n971), .A2(G50), .ZN(new_n1159));
  INV_X1    g0959(.A(G132), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n802), .A2(new_n1160), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n276), .B(new_n1161), .C1(G125), .C2(new_n786), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n791), .A2(G150), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n847), .A2(G128), .B1(new_n1163), .B2(KEYINPUT53), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1158), .A2(new_n1159), .A3(new_n1162), .A4(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1163), .A2(KEYINPUT53), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1154), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n778), .B(new_n1149), .C1(new_n762), .C2(new_n1167), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n1115), .A2(new_n1117), .A3(new_n1125), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1168), .B1(new_n1169), .B2(new_n776), .ZN(new_n1170));
  AND2_X1   g0970(.A1(new_n1146), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(G378));
  NAND2_X1  g0972(.A1(new_n273), .A2(new_n869), .ZN(new_n1173));
  XOR2_X1   g0973(.A(new_n326), .B(new_n1173), .Z(new_n1174));
  XNOR2_X1  g0974(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1174), .B(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n759), .ZN(new_n1178));
  INV_X1    g0978(.A(G124), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n507), .B1(new_n784), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n791), .A2(new_n1156), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n808), .B2(new_n854), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n803), .A2(G128), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n847), .A2(G125), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(new_n1160), .C2(new_n795), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n1182), .B(new_n1185), .C1(G150), .C2(new_n793), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT59), .ZN(new_n1187));
  AOI211_X1 g0987(.A(G33), .B(new_n1180), .C1(new_n1186), .C2(new_n1187), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1188), .B1(new_n1187), .B2(new_n1186), .C1(new_n975), .C2(new_n780), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n284), .B1(new_n796), .B2(G97), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1190), .B(new_n507), .C1(new_n219), .C2(new_n802), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n808), .A2(new_n385), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n785), .A2(new_n849), .ZN(new_n1193));
  NOR4_X1   g0993(.A1(new_n1191), .A2(new_n977), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n780), .A2(new_n223), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1045), .A2(new_n1195), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1194), .B(new_n1196), .C1(new_n483), .C2(new_n811), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT58), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n217), .B1(new_n274), .B2(G41), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1189), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n762), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n865), .A2(new_n217), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1178), .A2(new_n777), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT122), .ZN(new_n1207));
  INV_X1    g1007(.A(G330), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1208), .B(new_n903), .C1(new_n909), .C2(new_n910), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1177), .B1(new_n938), .B2(new_n939), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n931), .A2(new_n936), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(KEYINPUT112), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n931), .A2(new_n936), .A3(new_n937), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1212), .A2(new_n1213), .A3(new_n1176), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n1209), .A2(new_n1210), .A3(new_n1214), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1210), .A2(new_n1214), .B1(G330), .B2(new_n911), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1207), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n911), .A2(G330), .ZN(new_n1218));
  NOR3_X1   g1018(.A1(new_n938), .A2(new_n939), .A3(new_n1177), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1176), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1218), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1209), .A2(new_n1210), .A3(new_n1214), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1221), .A2(KEYINPUT122), .A3(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1217), .A2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1206), .B1(new_n1224), .B2(new_n776), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT123), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1142), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1128), .A2(KEYINPUT123), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n1169), .B2(new_n1144), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n1217), .B2(new_n1223), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n771), .B1(new_n1231), .B2(KEYINPUT57), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT124), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1221), .A2(KEYINPUT57), .A3(new_n1222), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1233), .B1(new_n1234), .B2(new_n1230), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1145), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1236), .A2(new_n1237), .A3(KEYINPUT124), .A4(KEYINPUT57), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1235), .A2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1225), .B1(new_n1232), .B2(new_n1239), .ZN(G375));
  NAND2_X1  g1040(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1033), .B(new_n1241), .C1(new_n1138), .C2(new_n1140), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1130), .A2(new_n758), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n865), .A2(new_n226), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n276), .B1(new_n786), .B2(G128), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n792), .A2(new_n217), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n1247), .B(new_n1195), .C1(G159), .C2(new_n791), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1246), .B(new_n1248), .C1(new_n855), .C2(new_n808), .ZN(new_n1249));
  XOR2_X1   g1049(.A(new_n1249), .B(KEYINPUT127), .Z(new_n1250));
  NAND3_X1  g1050(.A1(new_n847), .A2(KEYINPUT126), .A3(G132), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n803), .A2(G137), .ZN(new_n1252));
  AOI21_X1  g1052(.A(KEYINPUT126), .B1(new_n847), .B2(G132), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(new_n796), .B2(new_n1156), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1250), .A2(new_n1251), .A3(new_n1252), .A4(new_n1254), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n802), .A2(new_n849), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n276), .B1(new_n781), .B2(new_n279), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1257), .B(KEYINPUT125), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n795), .A2(new_n479), .B1(new_n811), .B2(new_n845), .ZN(new_n1259));
  AOI211_X1 g1059(.A(new_n1259), .B(new_n1046), .C1(new_n529), .C2(new_n807), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n786), .A2(G303), .B1(G97), .B2(new_n791), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1258), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1255), .B1(new_n1256), .B2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1245), .B1(new_n762), .B2(new_n1263), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n1137), .A2(new_n776), .B1(new_n1264), .B2(new_n777), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1242), .A2(new_n1265), .ZN(G381));
  OAI211_X1 g1066(.A(new_n1171), .B(new_n1225), .C1(new_n1232), .C2(new_n1239), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(new_n1267), .A2(G384), .A3(G381), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n988), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1064), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1269), .B1(new_n1271), .B2(new_n1008), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1098), .A2(new_n1272), .A3(new_n1099), .ZN(new_n1273));
  NOR3_X1   g1073(.A1(new_n1273), .A2(G396), .A3(G393), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1268), .A2(new_n1274), .ZN(G407));
  OAI211_X1 g1075(.A(G407), .B(G213), .C1(G343), .C2(new_n1267), .ZN(G409));
  AND3_X1   g1076(.A1(new_n1221), .A2(KEYINPUT122), .A3(new_n1222), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT122), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1033), .B(new_n1236), .C1(new_n1277), .C2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1237), .A2(new_n776), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1279), .A2(new_n1171), .A3(new_n1205), .A4(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n686), .A2(G213), .ZN(new_n1282));
  AND2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1224), .A2(new_n776), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1205), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1236), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT57), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n715), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1235), .A2(new_n1238), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1285), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1283), .B1(new_n1290), .B2(new_n1171), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT60), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1241), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1144), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1142), .A2(new_n1143), .A3(KEYINPUT60), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1293), .A2(new_n1294), .A3(new_n771), .A4(new_n1295), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1296), .A2(G384), .A3(new_n1265), .ZN(new_n1297));
  AOI21_X1  g1097(.A(G384), .B1(new_n1296), .B2(new_n1265), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n686), .A2(G213), .A3(G2897), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1300), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1302), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1301), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(KEYINPUT61), .B1(new_n1291), .B2(new_n1305), .ZN(new_n1306));
  OAI211_X1 g1106(.A(new_n1283), .B(new_n1299), .C1(new_n1290), .C2(new_n1171), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(KEYINPUT62), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(G375), .A2(G378), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT62), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1309), .A2(new_n1310), .A3(new_n1283), .A4(new_n1299), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1306), .A2(new_n1308), .A3(new_n1311), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(G393), .B(G396), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1071), .A2(KEYINPUT118), .A3(new_n1095), .ZN(new_n1315));
  AOI21_X1  g1115(.A(KEYINPUT118), .B1(new_n1071), .B2(new_n1095), .ZN(new_n1316));
  NOR3_X1   g1116(.A1(new_n1315), .A2(new_n1316), .A3(G387), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1272), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1314), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(G387), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1320), .A2(new_n1273), .A3(new_n1313), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1319), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1312), .A2(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1304), .B1(new_n1309), .B2(new_n1283), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT63), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1307), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT61), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1320), .A2(new_n1273), .A3(new_n1313), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1313), .B1(new_n1320), .B2(new_n1273), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1309), .A2(KEYINPUT63), .A3(new_n1283), .A4(new_n1299), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1326), .A2(new_n1327), .A3(new_n1330), .A4(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1323), .A2(new_n1332), .ZN(G405));
  NAND3_X1  g1133(.A1(new_n1322), .A2(new_n1267), .A3(new_n1309), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1309), .A2(new_n1267), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1330), .A2(new_n1335), .ZN(new_n1336));
  AND3_X1   g1136(.A1(new_n1334), .A2(new_n1336), .A3(new_n1299), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1299), .B1(new_n1334), .B2(new_n1336), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1337), .A2(new_n1338), .ZN(G402));
endmodule


