

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U556 ( .A1(n787), .A2(n788), .ZN(n523) );
  NOR2_X2 U557 ( .A1(n733), .A2(n732), .ZN(n739) );
  NOR2_X1 U558 ( .A1(G164), .A2(G1384), .ZN(n731) );
  XNOR2_X1 U559 ( .A(n786), .B(KEYINPUT104), .ZN(n800) );
  NOR2_X1 U560 ( .A1(n777), .A2(G168), .ZN(n778) );
  AND2_X1 U561 ( .A1(n806), .A2(n805), .ZN(n807) );
  NAND2_X1 U562 ( .A1(G8), .A2(n771), .ZN(n817) );
  NOR2_X2 U563 ( .A1(G2105), .A2(G2104), .ZN(n550) );
  AND2_X1 U564 ( .A1(n821), .A2(n820), .ZN(n822) );
  AND2_X1 U565 ( .A1(G8), .A2(n783), .ZN(n524) );
  OR2_X1 U566 ( .A1(n818), .A2(n817), .ZN(n525) );
  AND2_X1 U567 ( .A1(n775), .A2(n774), .ZN(n526) );
  INV_X1 U568 ( .A(G8), .ZN(n773) );
  NOR2_X1 U569 ( .A1(n939), .A2(n742), .ZN(n745) );
  NOR2_X1 U570 ( .A1(G2084), .A2(n771), .ZN(n772) );
  NOR2_X1 U571 ( .A1(n524), .A2(n784), .ZN(n785) );
  NAND2_X1 U572 ( .A1(n523), .A2(n785), .ZN(n786) );
  INV_X1 U573 ( .A(n739), .ZN(n771) );
  AND2_X1 U574 ( .A1(n819), .A2(n525), .ZN(n820) );
  NOR2_X1 U575 ( .A1(G543), .A2(n535), .ZN(n527) );
  NOR2_X1 U576 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U577 ( .A(KEYINPUT77), .B(n543), .Z(G168) );
  INV_X1 U578 ( .A(G651), .ZN(n535) );
  XOR2_X1 U579 ( .A(KEYINPUT1), .B(n527), .Z(n669) );
  NAND2_X1 U580 ( .A1(n669), .A2(G63), .ZN(n528) );
  XNOR2_X1 U581 ( .A(n528), .B(KEYINPUT76), .ZN(n531) );
  XOR2_X1 U582 ( .A(KEYINPUT0), .B(G543), .Z(n534) );
  NOR2_X1 U583 ( .A1(G651), .A2(n534), .ZN(n529) );
  XOR2_X2 U584 ( .A(KEYINPUT65), .B(n529), .Z(n664) );
  NAND2_X1 U585 ( .A1(G51), .A2(n664), .ZN(n530) );
  NAND2_X1 U586 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U587 ( .A(KEYINPUT6), .B(n532), .ZN(n541) );
  NOR2_X1 U588 ( .A1(G651), .A2(G543), .ZN(n655) );
  NAND2_X1 U589 ( .A1(n655), .A2(G89), .ZN(n533) );
  XNOR2_X1 U590 ( .A(n533), .B(KEYINPUT4), .ZN(n538) );
  OR2_X1 U591 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X2 U592 ( .A(KEYINPUT69), .B(n536), .ZN(n658) );
  NAND2_X1 U593 ( .A1(G76), .A2(n658), .ZN(n537) );
  NAND2_X1 U594 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U595 ( .A(n539), .B(KEYINPUT5), .Z(n540) );
  NOR2_X1 U596 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U597 ( .A(KEYINPUT7), .B(n542), .Z(n543) );
  INV_X1 U598 ( .A(G2104), .ZN(n551) );
  NOR2_X4 U599 ( .A1(G2105), .A2(n551), .ZN(n892) );
  NAND2_X1 U600 ( .A1(G101), .A2(n892), .ZN(n544) );
  XNOR2_X1 U601 ( .A(n544), .B(KEYINPUT23), .ZN(n546) );
  INV_X1 U602 ( .A(KEYINPUT66), .ZN(n545) );
  XNOR2_X1 U603 ( .A(n546), .B(n545), .ZN(n549) );
  NAND2_X1 U604 ( .A1(G2104), .A2(G2105), .ZN(n547) );
  XNOR2_X2 U605 ( .A(n547), .B(KEYINPUT67), .ZN(n897) );
  NAND2_X1 U606 ( .A1(G113), .A2(n897), .ZN(n548) );
  NAND2_X1 U607 ( .A1(n549), .A2(n548), .ZN(n555) );
  XOR2_X2 U608 ( .A(KEYINPUT17), .B(n550), .Z(n891) );
  NAND2_X1 U609 ( .A1(G137), .A2(n891), .ZN(n553) );
  AND2_X1 U610 ( .A1(n551), .A2(G2105), .ZN(n896) );
  NAND2_X1 U611 ( .A1(G125), .A2(n896), .ZN(n552) );
  NAND2_X1 U612 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X2 U613 ( .A1(n555), .A2(n554), .ZN(G160) );
  NAND2_X1 U614 ( .A1(G138), .A2(n891), .ZN(n557) );
  NAND2_X1 U615 ( .A1(G102), .A2(n892), .ZN(n556) );
  NAND2_X1 U616 ( .A1(n557), .A2(n556), .ZN(n561) );
  NAND2_X1 U617 ( .A1(G126), .A2(n896), .ZN(n559) );
  NAND2_X1 U618 ( .A1(G114), .A2(n897), .ZN(n558) );
  NAND2_X1 U619 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U620 ( .A1(n561), .A2(n560), .ZN(G164) );
  XOR2_X1 U621 ( .A(G2443), .B(G2446), .Z(n563) );
  XNOR2_X1 U622 ( .A(G2427), .B(G2451), .ZN(n562) );
  XNOR2_X1 U623 ( .A(n563), .B(n562), .ZN(n569) );
  XOR2_X1 U624 ( .A(G2430), .B(G2454), .Z(n565) );
  XNOR2_X1 U625 ( .A(G1341), .B(G1348), .ZN(n564) );
  XNOR2_X1 U626 ( .A(n565), .B(n564), .ZN(n567) );
  XOR2_X1 U627 ( .A(G2435), .B(G2438), .Z(n566) );
  XNOR2_X1 U628 ( .A(n567), .B(n566), .ZN(n568) );
  XOR2_X1 U629 ( .A(n569), .B(n568), .Z(n570) );
  AND2_X1 U630 ( .A1(G14), .A2(n570), .ZN(G401) );
  AND2_X1 U631 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U632 ( .A(G120), .ZN(G236) );
  INV_X1 U633 ( .A(G108), .ZN(G238) );
  INV_X1 U634 ( .A(G132), .ZN(G219) );
  INV_X1 U635 ( .A(G82), .ZN(G220) );
  NAND2_X1 U636 ( .A1(G7), .A2(G661), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(KEYINPUT72), .ZN(n572) );
  XOR2_X1 U638 ( .A(KEYINPUT10), .B(n572), .Z(n842) );
  INV_X1 U639 ( .A(n842), .ZN(G223) );
  INV_X1 U640 ( .A(G567), .ZN(n697) );
  NOR2_X1 U641 ( .A1(G223), .A2(n697), .ZN(n573) );
  XNOR2_X1 U642 ( .A(n573), .B(KEYINPUT11), .ZN(G234) );
  NAND2_X1 U643 ( .A1(n655), .A2(G81), .ZN(n574) );
  XNOR2_X1 U644 ( .A(n574), .B(KEYINPUT12), .ZN(n576) );
  NAND2_X1 U645 ( .A1(G68), .A2(n658), .ZN(n575) );
  NAND2_X1 U646 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U647 ( .A(KEYINPUT13), .B(n577), .ZN(n583) );
  NAND2_X1 U648 ( .A1(G56), .A2(n669), .ZN(n578) );
  XOR2_X1 U649 ( .A(KEYINPUT14), .B(n578), .Z(n581) );
  NAND2_X1 U650 ( .A1(G43), .A2(n664), .ZN(n579) );
  XNOR2_X1 U651 ( .A(KEYINPUT73), .B(n579), .ZN(n580) );
  NAND2_X1 U652 ( .A1(n583), .A2(n582), .ZN(n939) );
  INV_X1 U653 ( .A(G860), .ZN(n614) );
  OR2_X1 U654 ( .A1(n939), .A2(n614), .ZN(G153) );
  NAND2_X1 U655 ( .A1(G64), .A2(n669), .ZN(n585) );
  NAND2_X1 U656 ( .A1(G52), .A2(n664), .ZN(n584) );
  NAND2_X1 U657 ( .A1(n585), .A2(n584), .ZN(n590) );
  NAND2_X1 U658 ( .A1(G77), .A2(n658), .ZN(n587) );
  NAND2_X1 U659 ( .A1(G90), .A2(n655), .ZN(n586) );
  NAND2_X1 U660 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U661 ( .A(KEYINPUT9), .B(n588), .Z(n589) );
  NOR2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U663 ( .A(KEYINPUT71), .B(n591), .ZN(G301) );
  NAND2_X1 U664 ( .A1(G301), .A2(G868), .ZN(n592) );
  XNOR2_X1 U665 ( .A(n592), .B(KEYINPUT74), .ZN(n602) );
  INV_X1 U666 ( .A(G868), .ZN(n683) );
  NAND2_X1 U667 ( .A1(n664), .A2(G54), .ZN(n599) );
  NAND2_X1 U668 ( .A1(G79), .A2(n658), .ZN(n594) );
  NAND2_X1 U669 ( .A1(G66), .A2(n669), .ZN(n593) );
  NAND2_X1 U670 ( .A1(n594), .A2(n593), .ZN(n597) );
  NAND2_X1 U671 ( .A1(G92), .A2(n655), .ZN(n595) );
  XNOR2_X1 U672 ( .A(KEYINPUT75), .B(n595), .ZN(n596) );
  NOR2_X1 U673 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U674 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U675 ( .A(KEYINPUT15), .B(n600), .ZN(n938) );
  INV_X1 U676 ( .A(n938), .ZN(n749) );
  NAND2_X1 U677 ( .A1(n683), .A2(n749), .ZN(n601) );
  NAND2_X1 U678 ( .A1(n602), .A2(n601), .ZN(G284) );
  XOR2_X1 U679 ( .A(G168), .B(KEYINPUT8), .Z(n603) );
  XNOR2_X1 U680 ( .A(KEYINPUT78), .B(n603), .ZN(G286) );
  NAND2_X1 U681 ( .A1(G65), .A2(n669), .ZN(n605) );
  NAND2_X1 U682 ( .A1(G53), .A2(n664), .ZN(n604) );
  NAND2_X1 U683 ( .A1(n605), .A2(n604), .ZN(n609) );
  NAND2_X1 U684 ( .A1(G78), .A2(n658), .ZN(n607) );
  NAND2_X1 U685 ( .A1(G91), .A2(n655), .ZN(n606) );
  NAND2_X1 U686 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U687 ( .A1(n609), .A2(n608), .ZN(n760) );
  INV_X1 U688 ( .A(n760), .ZN(G299) );
  XOR2_X1 U689 ( .A(KEYINPUT79), .B(n683), .Z(n610) );
  NOR2_X1 U690 ( .A1(G286), .A2(n610), .ZN(n613) );
  NOR2_X1 U691 ( .A1(G868), .A2(G299), .ZN(n611) );
  XNOR2_X1 U692 ( .A(n611), .B(KEYINPUT80), .ZN(n612) );
  NOR2_X1 U693 ( .A1(n613), .A2(n612), .ZN(G297) );
  NAND2_X1 U694 ( .A1(n614), .A2(G559), .ZN(n615) );
  NAND2_X1 U695 ( .A1(n615), .A2(n938), .ZN(n616) );
  XNOR2_X1 U696 ( .A(n616), .B(KEYINPUT81), .ZN(n617) );
  XOR2_X1 U697 ( .A(KEYINPUT16), .B(n617), .Z(G148) );
  NOR2_X1 U698 ( .A1(G868), .A2(n939), .ZN(n620) );
  NAND2_X1 U699 ( .A1(G868), .A2(n938), .ZN(n618) );
  NOR2_X1 U700 ( .A1(G559), .A2(n618), .ZN(n619) );
  NOR2_X1 U701 ( .A1(n620), .A2(n619), .ZN(G282) );
  XOR2_X1 U702 ( .A(KEYINPUT82), .B(KEYINPUT18), .Z(n622) );
  NAND2_X1 U703 ( .A1(G123), .A2(n896), .ZN(n621) );
  XNOR2_X1 U704 ( .A(n622), .B(n621), .ZN(n626) );
  NAND2_X1 U705 ( .A1(G135), .A2(n891), .ZN(n624) );
  NAND2_X1 U706 ( .A1(G111), .A2(n897), .ZN(n623) );
  NAND2_X1 U707 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U708 ( .A1(n626), .A2(n625), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n892), .A2(G99), .ZN(n627) );
  NAND2_X1 U710 ( .A1(n628), .A2(n627), .ZN(n999) );
  XOR2_X1 U711 ( .A(n999), .B(G2096), .Z(n630) );
  XNOR2_X1 U712 ( .A(G2100), .B(KEYINPUT83), .ZN(n629) );
  NAND2_X1 U713 ( .A1(n630), .A2(n629), .ZN(G156) );
  NAND2_X1 U714 ( .A1(n938), .A2(G559), .ZN(n680) );
  XNOR2_X1 U715 ( .A(n939), .B(n680), .ZN(n631) );
  NOR2_X1 U716 ( .A1(n631), .A2(G860), .ZN(n638) );
  NAND2_X1 U717 ( .A1(G80), .A2(n658), .ZN(n633) );
  NAND2_X1 U718 ( .A1(G93), .A2(n655), .ZN(n632) );
  NAND2_X1 U719 ( .A1(n633), .A2(n632), .ZN(n637) );
  NAND2_X1 U720 ( .A1(G67), .A2(n669), .ZN(n635) );
  NAND2_X1 U721 ( .A1(G55), .A2(n664), .ZN(n634) );
  NAND2_X1 U722 ( .A1(n635), .A2(n634), .ZN(n636) );
  OR2_X1 U723 ( .A1(n637), .A2(n636), .ZN(n682) );
  XOR2_X1 U724 ( .A(n638), .B(n682), .Z(G145) );
  NAND2_X1 U725 ( .A1(G47), .A2(n664), .ZN(n639) );
  XNOR2_X1 U726 ( .A(n639), .B(KEYINPUT70), .ZN(n641) );
  NAND2_X1 U727 ( .A1(n658), .A2(G72), .ZN(n640) );
  NAND2_X1 U728 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U729 ( .A1(G85), .A2(n655), .ZN(n642) );
  XOR2_X1 U730 ( .A(KEYINPUT68), .B(n642), .Z(n643) );
  NOR2_X1 U731 ( .A1(n644), .A2(n643), .ZN(n646) );
  NAND2_X1 U732 ( .A1(n669), .A2(G60), .ZN(n645) );
  NAND2_X1 U733 ( .A1(n646), .A2(n645), .ZN(G290) );
  NAND2_X1 U734 ( .A1(n658), .A2(G75), .ZN(n653) );
  NAND2_X1 U735 ( .A1(G88), .A2(n655), .ZN(n648) );
  NAND2_X1 U736 ( .A1(G62), .A2(n669), .ZN(n647) );
  NAND2_X1 U737 ( .A1(n648), .A2(n647), .ZN(n651) );
  NAND2_X1 U738 ( .A1(n664), .A2(G50), .ZN(n649) );
  XOR2_X1 U739 ( .A(KEYINPUT86), .B(n649), .Z(n650) );
  NOR2_X1 U740 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U741 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U742 ( .A(KEYINPUT87), .B(n654), .ZN(G166) );
  INV_X1 U743 ( .A(G166), .ZN(G303) );
  NAND2_X1 U744 ( .A1(G86), .A2(n655), .ZN(n657) );
  NAND2_X1 U745 ( .A1(G61), .A2(n669), .ZN(n656) );
  NAND2_X1 U746 ( .A1(n657), .A2(n656), .ZN(n661) );
  NAND2_X1 U747 ( .A1(n658), .A2(G73), .ZN(n659) );
  XOR2_X1 U748 ( .A(KEYINPUT2), .B(n659), .Z(n660) );
  NOR2_X1 U749 ( .A1(n661), .A2(n660), .ZN(n663) );
  NAND2_X1 U750 ( .A1(n664), .A2(G48), .ZN(n662) );
  NAND2_X1 U751 ( .A1(n663), .A2(n662), .ZN(G305) );
  NAND2_X1 U752 ( .A1(G49), .A2(n664), .ZN(n666) );
  NAND2_X1 U753 ( .A1(G74), .A2(G651), .ZN(n665) );
  NAND2_X1 U754 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U755 ( .A(KEYINPUT84), .B(n667), .ZN(n668) );
  NOR2_X1 U756 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U757 ( .A(KEYINPUT85), .B(n670), .Z(n672) );
  NAND2_X1 U758 ( .A1(n534), .A2(G87), .ZN(n671) );
  NAND2_X1 U759 ( .A1(n672), .A2(n671), .ZN(G288) );
  XOR2_X1 U760 ( .A(KEYINPUT19), .B(KEYINPUT88), .Z(n673) );
  XNOR2_X1 U761 ( .A(G305), .B(n673), .ZN(n674) );
  XOR2_X1 U762 ( .A(G303), .B(n674), .Z(n676) );
  XOR2_X1 U763 ( .A(n939), .B(G299), .Z(n675) );
  XNOR2_X1 U764 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U765 ( .A(n682), .B(n677), .ZN(n678) );
  XNOR2_X1 U766 ( .A(G290), .B(n678), .ZN(n679) );
  XNOR2_X1 U767 ( .A(n679), .B(G288), .ZN(n913) );
  XNOR2_X1 U768 ( .A(n680), .B(n913), .ZN(n681) );
  NAND2_X1 U769 ( .A1(n681), .A2(G868), .ZN(n685) );
  NAND2_X1 U770 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U771 ( .A1(n685), .A2(n684), .ZN(G295) );
  NAND2_X1 U772 ( .A1(G2078), .A2(G2084), .ZN(n686) );
  XOR2_X1 U773 ( .A(KEYINPUT20), .B(n686), .Z(n687) );
  NAND2_X1 U774 ( .A1(G2090), .A2(n687), .ZN(n688) );
  XNOR2_X1 U775 ( .A(KEYINPUT21), .B(n688), .ZN(n689) );
  NAND2_X1 U776 ( .A1(n689), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U777 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U778 ( .A1(G220), .A2(G219), .ZN(n690) );
  XOR2_X1 U779 ( .A(KEYINPUT22), .B(n690), .Z(n691) );
  NOR2_X1 U780 ( .A1(G218), .A2(n691), .ZN(n692) );
  NAND2_X1 U781 ( .A1(G96), .A2(n692), .ZN(n849) );
  NAND2_X1 U782 ( .A1(G2106), .A2(n849), .ZN(n693) );
  XNOR2_X1 U783 ( .A(n693), .B(KEYINPUT89), .ZN(n699) );
  NAND2_X1 U784 ( .A1(G69), .A2(G57), .ZN(n694) );
  NOR2_X1 U785 ( .A1(G236), .A2(n694), .ZN(n695) );
  XOR2_X1 U786 ( .A(KEYINPUT90), .B(n695), .Z(n696) );
  NOR2_X1 U787 ( .A1(G238), .A2(n696), .ZN(n848) );
  NOR2_X1 U788 ( .A1(n697), .A2(n848), .ZN(n698) );
  NOR2_X1 U789 ( .A1(n699), .A2(n698), .ZN(G319) );
  INV_X1 U790 ( .A(G319), .ZN(n701) );
  NAND2_X1 U791 ( .A1(G483), .A2(G661), .ZN(n700) );
  NOR2_X1 U792 ( .A1(n701), .A2(n700), .ZN(n847) );
  NAND2_X1 U793 ( .A1(n847), .A2(G36), .ZN(G176) );
  NAND2_X1 U794 ( .A1(G160), .A2(G40), .ZN(n733) );
  NOR2_X1 U795 ( .A1(n731), .A2(n733), .ZN(n837) );
  XNOR2_X1 U796 ( .A(G2067), .B(KEYINPUT37), .ZN(n835) );
  NAND2_X1 U797 ( .A1(G140), .A2(n891), .ZN(n703) );
  NAND2_X1 U798 ( .A1(G104), .A2(n892), .ZN(n702) );
  NAND2_X1 U799 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U800 ( .A(KEYINPUT34), .B(n704), .ZN(n710) );
  NAND2_X1 U801 ( .A1(G128), .A2(n896), .ZN(n706) );
  NAND2_X1 U802 ( .A1(G116), .A2(n897), .ZN(n705) );
  NAND2_X1 U803 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U804 ( .A(KEYINPUT91), .B(n707), .ZN(n708) );
  XNOR2_X1 U805 ( .A(KEYINPUT35), .B(n708), .ZN(n709) );
  NOR2_X1 U806 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U807 ( .A(KEYINPUT36), .B(n711), .ZN(n903) );
  NOR2_X1 U808 ( .A1(n835), .A2(n903), .ZN(n1006) );
  NAND2_X1 U809 ( .A1(n837), .A2(n1006), .ZN(n833) );
  NAND2_X1 U810 ( .A1(G129), .A2(n896), .ZN(n713) );
  NAND2_X1 U811 ( .A1(G117), .A2(n897), .ZN(n712) );
  NAND2_X1 U812 ( .A1(n713), .A2(n712), .ZN(n717) );
  NAND2_X1 U813 ( .A1(G105), .A2(n892), .ZN(n714) );
  XNOR2_X1 U814 ( .A(n714), .B(KEYINPUT38), .ZN(n715) );
  XNOR2_X1 U815 ( .A(n715), .B(KEYINPUT93), .ZN(n716) );
  NOR2_X1 U816 ( .A1(n717), .A2(n716), .ZN(n719) );
  NAND2_X1 U817 ( .A1(n891), .A2(G141), .ZN(n718) );
  NAND2_X1 U818 ( .A1(n719), .A2(n718), .ZN(n906) );
  NAND2_X1 U819 ( .A1(G1996), .A2(n906), .ZN(n720) );
  XOR2_X1 U820 ( .A(KEYINPUT94), .B(n720), .Z(n729) );
  NAND2_X1 U821 ( .A1(G119), .A2(n896), .ZN(n722) );
  NAND2_X1 U822 ( .A1(G107), .A2(n897), .ZN(n721) );
  NAND2_X1 U823 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U824 ( .A(KEYINPUT92), .B(n723), .ZN(n727) );
  NAND2_X1 U825 ( .A1(G131), .A2(n891), .ZN(n725) );
  NAND2_X1 U826 ( .A1(G95), .A2(n892), .ZN(n724) );
  NAND2_X1 U827 ( .A1(n725), .A2(n724), .ZN(n726) );
  OR2_X1 U828 ( .A1(n727), .A2(n726), .ZN(n887) );
  AND2_X1 U829 ( .A1(n887), .A2(G1991), .ZN(n728) );
  NOR2_X1 U830 ( .A1(n729), .A2(n728), .ZN(n1008) );
  INV_X1 U831 ( .A(n1008), .ZN(n730) );
  NAND2_X1 U832 ( .A1(n730), .A2(n837), .ZN(n827) );
  NAND2_X1 U833 ( .A1(n833), .A2(n827), .ZN(n823) );
  INV_X1 U834 ( .A(n731), .ZN(n732) );
  NOR2_X1 U835 ( .A1(G1976), .A2(G288), .ZN(n802) );
  NAND2_X1 U836 ( .A1(n802), .A2(KEYINPUT33), .ZN(n734) );
  NOR2_X1 U837 ( .A1(n817), .A2(n734), .ZN(n809) );
  NAND2_X1 U838 ( .A1(G2067), .A2(n739), .ZN(n735) );
  XOR2_X1 U839 ( .A(KEYINPUT99), .B(n735), .Z(n737) );
  NAND2_X1 U840 ( .A1(G1348), .A2(n771), .ZN(n736) );
  NAND2_X1 U841 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U842 ( .A(KEYINPUT100), .B(n738), .Z(n747) );
  NAND2_X1 U843 ( .A1(G1996), .A2(n739), .ZN(n741) );
  XNOR2_X1 U844 ( .A(KEYINPUT64), .B(KEYINPUT26), .ZN(n740) );
  XOR2_X1 U845 ( .A(n741), .B(n740), .Z(n742) );
  NAND2_X1 U846 ( .A1(G1341), .A2(n771), .ZN(n743) );
  XNOR2_X1 U847 ( .A(KEYINPUT98), .B(n743), .ZN(n744) );
  NAND2_X1 U848 ( .A1(n745), .A2(n744), .ZN(n750) );
  NOR2_X1 U849 ( .A1(n749), .A2(n750), .ZN(n746) );
  NOR2_X1 U850 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U851 ( .A(n748), .B(KEYINPUT101), .ZN(n752) );
  NAND2_X1 U852 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U853 ( .A1(n752), .A2(n751), .ZN(n758) );
  NAND2_X1 U854 ( .A1(G1956), .A2(n771), .ZN(n753) );
  XNOR2_X1 U855 ( .A(KEYINPUT97), .B(n753), .ZN(n756) );
  INV_X1 U856 ( .A(n771), .ZN(n766) );
  NAND2_X1 U857 ( .A1(n766), .A2(G2072), .ZN(n754) );
  XNOR2_X1 U858 ( .A(KEYINPUT27), .B(n754), .ZN(n755) );
  NOR2_X1 U859 ( .A1(n756), .A2(n755), .ZN(n759) );
  NAND2_X1 U860 ( .A1(n760), .A2(n759), .ZN(n757) );
  NAND2_X1 U861 ( .A1(n758), .A2(n757), .ZN(n763) );
  NOR2_X1 U862 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U863 ( .A(n761), .B(KEYINPUT28), .Z(n762) );
  NAND2_X1 U864 ( .A1(n763), .A2(n762), .ZN(n765) );
  XOR2_X1 U865 ( .A(KEYINPUT29), .B(KEYINPUT102), .Z(n764) );
  XNOR2_X1 U866 ( .A(n765), .B(n764), .ZN(n770) );
  XOR2_X1 U867 ( .A(KEYINPUT25), .B(G2078), .Z(n976) );
  NOR2_X1 U868 ( .A1(n976), .A2(n771), .ZN(n768) );
  NOR2_X1 U869 ( .A1(n766), .A2(G1961), .ZN(n767) );
  NOR2_X1 U870 ( .A1(n768), .A2(n767), .ZN(n779) );
  OR2_X1 U871 ( .A1(n779), .A2(G301), .ZN(n769) );
  NAND2_X1 U872 ( .A1(n770), .A2(n769), .ZN(n787) );
  INV_X1 U873 ( .A(KEYINPUT30), .ZN(n776) );
  XNOR2_X1 U874 ( .A(n772), .B(KEYINPUT96), .ZN(n783) );
  INV_X1 U875 ( .A(n783), .ZN(n775) );
  NOR2_X1 U876 ( .A1(G1966), .A2(n817), .ZN(n784) );
  NOR2_X1 U877 ( .A1(n784), .A2(n773), .ZN(n774) );
  XNOR2_X1 U878 ( .A(n776), .B(n526), .ZN(n777) );
  XNOR2_X1 U879 ( .A(n778), .B(KEYINPUT103), .ZN(n781) );
  NAND2_X1 U880 ( .A1(n779), .A2(G301), .ZN(n780) );
  NAND2_X1 U881 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U882 ( .A(n782), .B(KEYINPUT31), .ZN(n788) );
  NAND2_X1 U883 ( .A1(n788), .A2(n787), .ZN(n789) );
  NAND2_X1 U884 ( .A1(n789), .A2(G286), .ZN(n796) );
  NOR2_X1 U885 ( .A1(G1971), .A2(n817), .ZN(n790) );
  XNOR2_X1 U886 ( .A(KEYINPUT105), .B(n790), .ZN(n794) );
  NOR2_X1 U887 ( .A1(G2090), .A2(n771), .ZN(n791) );
  XNOR2_X1 U888 ( .A(KEYINPUT106), .B(n791), .ZN(n792) );
  NOR2_X1 U889 ( .A1(G166), .A2(n792), .ZN(n793) );
  NAND2_X1 U890 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U891 ( .A1(n796), .A2(n795), .ZN(n797) );
  NAND2_X1 U892 ( .A1(n797), .A2(G8), .ZN(n798) );
  XNOR2_X1 U893 ( .A(n798), .B(KEYINPUT32), .ZN(n799) );
  NAND2_X1 U894 ( .A1(n800), .A2(n799), .ZN(n811) );
  NOR2_X1 U895 ( .A1(G1971), .A2(G303), .ZN(n801) );
  NOR2_X1 U896 ( .A1(n802), .A2(n801), .ZN(n932) );
  NAND2_X1 U897 ( .A1(n811), .A2(n932), .ZN(n806) );
  INV_X1 U898 ( .A(n817), .ZN(n804) );
  NAND2_X1 U899 ( .A1(G288), .A2(G1976), .ZN(n803) );
  XOR2_X1 U900 ( .A(KEYINPUT107), .B(n803), .Z(n931) );
  AND2_X1 U901 ( .A1(n804), .A2(n931), .ZN(n805) );
  NOR2_X1 U902 ( .A1(KEYINPUT33), .A2(n807), .ZN(n808) );
  NOR2_X1 U903 ( .A1(n809), .A2(n808), .ZN(n810) );
  XOR2_X1 U904 ( .A(G1981), .B(G305), .Z(n924) );
  NAND2_X1 U905 ( .A1(n810), .A2(n924), .ZN(n821) );
  NOR2_X1 U906 ( .A1(G2090), .A2(G303), .ZN(n812) );
  NAND2_X1 U907 ( .A1(G8), .A2(n812), .ZN(n813) );
  NAND2_X1 U908 ( .A1(n811), .A2(n813), .ZN(n814) );
  NAND2_X1 U909 ( .A1(n814), .A2(n817), .ZN(n819) );
  NOR2_X1 U910 ( .A1(G1981), .A2(G305), .ZN(n815) );
  XNOR2_X1 U911 ( .A(n815), .B(KEYINPUT95), .ZN(n816) );
  XNOR2_X1 U912 ( .A(n816), .B(KEYINPUT24), .ZN(n818) );
  NOR2_X1 U913 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U914 ( .A(n824), .B(KEYINPUT108), .ZN(n826) );
  XNOR2_X1 U915 ( .A(G1986), .B(G290), .ZN(n944) );
  NAND2_X1 U916 ( .A1(n944), .A2(n837), .ZN(n825) );
  NAND2_X1 U917 ( .A1(n826), .A2(n825), .ZN(n840) );
  NOR2_X1 U918 ( .A1(G1996), .A2(n906), .ZN(n997) );
  INV_X1 U919 ( .A(n827), .ZN(n830) );
  NOR2_X1 U920 ( .A1(G1986), .A2(G290), .ZN(n828) );
  NOR2_X1 U921 ( .A1(G1991), .A2(n887), .ZN(n1002) );
  NOR2_X1 U922 ( .A1(n828), .A2(n1002), .ZN(n829) );
  NOR2_X1 U923 ( .A1(n830), .A2(n829), .ZN(n831) );
  NOR2_X1 U924 ( .A1(n997), .A2(n831), .ZN(n832) );
  XNOR2_X1 U925 ( .A(n832), .B(KEYINPUT39), .ZN(n834) );
  NAND2_X1 U926 ( .A1(n834), .A2(n833), .ZN(n836) );
  NAND2_X1 U927 ( .A1(n835), .A2(n903), .ZN(n1010) );
  NAND2_X1 U928 ( .A1(n836), .A2(n1010), .ZN(n838) );
  NAND2_X1 U929 ( .A1(n838), .A2(n837), .ZN(n839) );
  NAND2_X1 U930 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U931 ( .A(n841), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U932 ( .A1(G2106), .A2(n842), .ZN(G217) );
  NAND2_X1 U933 ( .A1(G15), .A2(G2), .ZN(n844) );
  INV_X1 U934 ( .A(G661), .ZN(n843) );
  NOR2_X1 U935 ( .A1(n844), .A2(n843), .ZN(n845) );
  XNOR2_X1 U936 ( .A(n845), .B(KEYINPUT109), .ZN(G259) );
  NAND2_X1 U937 ( .A1(G3), .A2(G1), .ZN(n846) );
  NAND2_X1 U938 ( .A1(n847), .A2(n846), .ZN(G188) );
  XOR2_X1 U939 ( .A(G69), .B(KEYINPUT110), .Z(G235) );
  INV_X1 U941 ( .A(G96), .ZN(G221) );
  INV_X1 U942 ( .A(G57), .ZN(G237) );
  INV_X1 U943 ( .A(n848), .ZN(n850) );
  NOR2_X1 U944 ( .A1(n850), .A2(n849), .ZN(G325) );
  INV_X1 U945 ( .A(G325), .ZN(G261) );
  XOR2_X1 U946 ( .A(KEYINPUT114), .B(G1956), .Z(n852) );
  XNOR2_X1 U947 ( .A(G1996), .B(G1991), .ZN(n851) );
  XNOR2_X1 U948 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U949 ( .A(n853), .B(KEYINPUT41), .Z(n855) );
  XNOR2_X1 U950 ( .A(G1986), .B(G1961), .ZN(n854) );
  XNOR2_X1 U951 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U952 ( .A(G1976), .B(G1981), .Z(n857) );
  XNOR2_X1 U953 ( .A(G1966), .B(G1971), .ZN(n856) );
  XNOR2_X1 U954 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U955 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U956 ( .A(G2474), .B(KEYINPUT115), .ZN(n860) );
  XNOR2_X1 U957 ( .A(n861), .B(n860), .ZN(G229) );
  XNOR2_X1 U958 ( .A(G2067), .B(G2078), .ZN(n862) );
  XNOR2_X1 U959 ( .A(n862), .B(KEYINPUT42), .ZN(n872) );
  XOR2_X1 U960 ( .A(KEYINPUT113), .B(G2678), .Z(n864) );
  XNOR2_X1 U961 ( .A(KEYINPUT112), .B(G2096), .ZN(n863) );
  XNOR2_X1 U962 ( .A(n864), .B(n863), .ZN(n868) );
  XOR2_X1 U963 ( .A(G2100), .B(G2090), .Z(n866) );
  XNOR2_X1 U964 ( .A(G2072), .B(G2084), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U966 ( .A(n868), .B(n867), .Z(n870) );
  XNOR2_X1 U967 ( .A(KEYINPUT43), .B(KEYINPUT111), .ZN(n869) );
  XNOR2_X1 U968 ( .A(n870), .B(n869), .ZN(n871) );
  XNOR2_X1 U969 ( .A(n872), .B(n871), .ZN(G227) );
  NAND2_X1 U970 ( .A1(n896), .A2(G124), .ZN(n873) );
  XNOR2_X1 U971 ( .A(n873), .B(KEYINPUT44), .ZN(n875) );
  NAND2_X1 U972 ( .A1(G112), .A2(n897), .ZN(n874) );
  NAND2_X1 U973 ( .A1(n875), .A2(n874), .ZN(n879) );
  NAND2_X1 U974 ( .A1(G136), .A2(n891), .ZN(n877) );
  NAND2_X1 U975 ( .A1(G100), .A2(n892), .ZN(n876) );
  NAND2_X1 U976 ( .A1(n877), .A2(n876), .ZN(n878) );
  NOR2_X1 U977 ( .A1(n879), .A2(n878), .ZN(G162) );
  NAND2_X1 U978 ( .A1(G130), .A2(n896), .ZN(n881) );
  NAND2_X1 U979 ( .A1(G118), .A2(n897), .ZN(n880) );
  NAND2_X1 U980 ( .A1(n881), .A2(n880), .ZN(n886) );
  NAND2_X1 U981 ( .A1(G142), .A2(n891), .ZN(n883) );
  NAND2_X1 U982 ( .A1(G106), .A2(n892), .ZN(n882) );
  NAND2_X1 U983 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U984 ( .A(KEYINPUT45), .B(n884), .Z(n885) );
  NOR2_X1 U985 ( .A1(n886), .A2(n885), .ZN(n890) );
  XNOR2_X1 U986 ( .A(G164), .B(n887), .ZN(n888) );
  XNOR2_X1 U987 ( .A(n888), .B(n999), .ZN(n889) );
  XNOR2_X1 U988 ( .A(n890), .B(n889), .ZN(n905) );
  NAND2_X1 U989 ( .A1(G139), .A2(n891), .ZN(n894) );
  NAND2_X1 U990 ( .A1(G103), .A2(n892), .ZN(n893) );
  NAND2_X1 U991 ( .A1(n894), .A2(n893), .ZN(n895) );
  XNOR2_X1 U992 ( .A(KEYINPUT116), .B(n895), .ZN(n902) );
  NAND2_X1 U993 ( .A1(G127), .A2(n896), .ZN(n899) );
  NAND2_X1 U994 ( .A1(G115), .A2(n897), .ZN(n898) );
  NAND2_X1 U995 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U996 ( .A(KEYINPUT47), .B(n900), .Z(n901) );
  NOR2_X1 U997 ( .A1(n902), .A2(n901), .ZN(n1012) );
  XNOR2_X1 U998 ( .A(n903), .B(n1012), .ZN(n904) );
  XNOR2_X1 U999 ( .A(n905), .B(n904), .ZN(n911) );
  XNOR2_X1 U1000 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n908) );
  XNOR2_X1 U1001 ( .A(n906), .B(G162), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1003 ( .A(G160), .B(n909), .Z(n910) );
  XNOR2_X1 U1004 ( .A(n911), .B(n910), .ZN(n912) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n912), .ZN(G395) );
  XOR2_X1 U1006 ( .A(KEYINPUT117), .B(n913), .Z(n915) );
  XOR2_X1 U1007 ( .A(G301), .B(n938), .Z(n914) );
  XNOR2_X1 U1008 ( .A(n915), .B(n914), .ZN(n916) );
  XOR2_X1 U1009 ( .A(n916), .B(G286), .Z(n917) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n917), .ZN(G397) );
  NOR2_X1 U1011 ( .A1(G229), .A2(G227), .ZN(n918) );
  XOR2_X1 U1012 ( .A(KEYINPUT49), .B(n918), .Z(n919) );
  NAND2_X1 U1013 ( .A1(G319), .A2(n919), .ZN(n920) );
  NOR2_X1 U1014 ( .A1(G401), .A2(n920), .ZN(n921) );
  XNOR2_X1 U1015 ( .A(KEYINPUT118), .B(n921), .ZN(n923) );
  NOR2_X1 U1016 ( .A1(G395), .A2(G397), .ZN(n922) );
  NAND2_X1 U1017 ( .A1(n923), .A2(n922), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(G301), .ZN(G171) );
  INV_X1 U1020 ( .A(G16), .ZN(n971) );
  XOR2_X1 U1021 ( .A(KEYINPUT56), .B(n971), .Z(n948) );
  XOR2_X1 U1022 ( .A(G301), .B(G1961), .Z(n928) );
  XNOR2_X1 U1023 ( .A(G1966), .B(G168), .ZN(n925) );
  NAND2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1025 ( .A(n926), .B(KEYINPUT57), .ZN(n927) );
  NAND2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n937) );
  XOR2_X1 U1027 ( .A(G299), .B(G1956), .Z(n930) );
  NAND2_X1 U1028 ( .A1(G1971), .A2(G303), .ZN(n929) );
  NAND2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n934) );
  NAND2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1032 ( .A(KEYINPUT124), .B(n935), .Z(n936) );
  NOR2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n946) );
  XNOR2_X1 U1034 ( .A(n938), .B(G1348), .ZN(n942) );
  XNOR2_X1 U1035 ( .A(KEYINPUT125), .B(n939), .ZN(n940) );
  XNOR2_X1 U1036 ( .A(G1341), .B(n940), .ZN(n941) );
  NAND2_X1 U1037 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1038 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1040 ( .A1(n948), .A2(n947), .ZN(n1027) );
  XNOR2_X1 U1041 ( .A(KEYINPUT60), .B(KEYINPUT126), .ZN(n958) );
  XOR2_X1 U1042 ( .A(G1348), .B(KEYINPUT59), .Z(n949) );
  XNOR2_X1 U1043 ( .A(G4), .B(n949), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(G6), .B(G1981), .ZN(n950) );
  NOR2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n955) );
  XNOR2_X1 U1046 ( .A(G1341), .B(G19), .ZN(n953) );
  XNOR2_X1 U1047 ( .A(G1956), .B(G20), .ZN(n952) );
  NOR2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(n956), .B(KEYINPUT127), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(n958), .B(n957), .ZN(n962) );
  XNOR2_X1 U1052 ( .A(G1966), .B(G21), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(G1961), .B(G5), .ZN(n959) );
  NOR2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n969) );
  XNOR2_X1 U1056 ( .A(G1971), .B(G22), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(G23), .B(G1976), .ZN(n963) );
  NOR2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n966) );
  XOR2_X1 U1059 ( .A(G1986), .B(G24), .Z(n965) );
  NAND2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1061 ( .A(KEYINPUT58), .B(n967), .ZN(n968) );
  NOR2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1063 ( .A(KEYINPUT61), .B(n970), .ZN(n972) );
  NAND2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1065 ( .A1(n973), .A2(G11), .ZN(n1025) );
  XOR2_X1 U1066 ( .A(G2090), .B(G35), .Z(n988) );
  XNOR2_X1 U1067 ( .A(G2067), .B(G26), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(G32), .B(G1996), .ZN(n974) );
  NOR2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n980) );
  XNOR2_X1 U1070 ( .A(n976), .B(G27), .ZN(n978) );
  XNOR2_X1 U1071 ( .A(G2072), .B(G33), .ZN(n977) );
  NOR2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n984) );
  XOR2_X1 U1074 ( .A(G1991), .B(G25), .Z(n981) );
  NAND2_X1 U1075 ( .A1(n981), .A2(G28), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(n982), .B(KEYINPUT120), .ZN(n983) );
  NOR2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1078 ( .A(n985), .B(KEYINPUT53), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(n986), .B(KEYINPUT121), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n991) );
  XNOR2_X1 U1081 ( .A(G34), .B(G2084), .ZN(n989) );
  XNOR2_X1 U1082 ( .A(KEYINPUT54), .B(n989), .ZN(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  INV_X1 U1084 ( .A(KEYINPUT55), .ZN(n1019) );
  XNOR2_X1 U1085 ( .A(n992), .B(n1019), .ZN(n993) );
  XNOR2_X1 U1086 ( .A(KEYINPUT122), .B(n993), .ZN(n994) );
  NOR2_X1 U1087 ( .A1(G29), .A2(n994), .ZN(n995) );
  XNOR2_X1 U1088 ( .A(n995), .B(KEYINPUT123), .ZN(n1023) );
  XOR2_X1 U1089 ( .A(G2090), .B(G162), .Z(n996) );
  NOR2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1091 ( .A(KEYINPUT51), .B(n998), .Z(n1004) );
  XNOR2_X1 U1092 ( .A(G160), .B(G2084), .ZN(n1000) );
  NAND2_X1 U1093 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(n1009), .B(KEYINPUT119), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1017) );
  XOR2_X1 U1100 ( .A(G2072), .B(n1012), .Z(n1014) );
  XOR2_X1 U1101 ( .A(G164), .B(G2078), .Z(n1013) );
  NOR2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1103 ( .A(KEYINPUT50), .B(n1015), .Z(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1105 ( .A(n1018), .B(KEYINPUT52), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1107 ( .A1(G29), .A2(n1021), .ZN(n1022) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1109 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1110 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1111 ( .A(KEYINPUT62), .B(n1028), .ZN(G150) );
  INV_X1 U1112 ( .A(G150), .ZN(G311) );
endmodule

