//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n777, new_n778,
    new_n779, new_n781, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n868, new_n869, new_n870,
    new_n872, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n986, new_n987;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT1), .ZN(new_n203));
  INV_X1    g002(.A(G113gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n204), .A2(G120gat), .ZN(new_n205));
  INV_X1    g004(.A(G120gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n206), .A2(G113gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n203), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  OR2_X1    g007(.A1(KEYINPUT69), .A2(G127gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(KEYINPUT69), .A2(G127gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(G134gat), .A3(new_n210), .ZN(new_n211));
  OR2_X1    g010(.A1(KEYINPUT68), .A2(G134gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(KEYINPUT68), .A2(G134gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n212), .A2(G127gat), .A3(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n208), .A2(new_n211), .A3(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G127gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n216), .A2(G134gat), .ZN(new_n217));
  INV_X1    g016(.A(G134gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(G127gat), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT70), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n206), .A2(G113gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n204), .A2(G120gat), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT1), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n218), .A2(G127gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n216), .A2(G134gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT70), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n220), .A2(new_n223), .A3(new_n227), .ZN(new_n228));
  AND2_X1   g027(.A1(new_n215), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G183gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT27), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT27), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G183gat), .ZN(new_n233));
  INV_X1    g032(.A(G190gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n231), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT28), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT66), .B1(new_n236), .B2(KEYINPUT28), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT28), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n240), .A2(new_n241), .A3(KEYINPUT65), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n238), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G169gat), .ZN(new_n245));
  INV_X1    g044(.A(G176gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(G169gat), .A2(G176gat), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n247), .B(KEYINPUT67), .C1(new_n249), .C2(KEYINPUT26), .ZN(new_n250));
  NOR2_X1   g049(.A1(G169gat), .A2(G176gat), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT26), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n254), .B1(new_n255), .B2(new_n251), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n250), .A2(new_n253), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(G183gat), .A2(G190gat), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n235), .A2(new_n237), .A3(new_n239), .A4(new_n242), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n244), .A2(new_n257), .A3(new_n258), .A4(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n230), .A2(new_n234), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n261), .A2(KEYINPUT24), .A3(new_n258), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT64), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT23), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n264), .B1(G169gat), .B2(G176gat), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT24), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(G183gat), .A3(G190gat), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n262), .A2(new_n263), .A3(new_n265), .A4(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n258), .A2(KEYINPUT24), .ZN(new_n269));
  NOR2_X1   g068(.A1(G183gat), .A2(G190gat), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n265), .A2(new_n267), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n249), .B1(KEYINPUT23), .B2(new_n251), .ZN(new_n274));
  AOI22_X1  g073(.A1(KEYINPUT25), .A2(new_n268), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n265), .B(new_n267), .C1(new_n269), .C2(new_n270), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n248), .B1(new_n247), .B2(new_n264), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT25), .ZN(new_n278));
  NOR4_X1   g077(.A1(new_n276), .A2(new_n277), .A3(new_n263), .A4(new_n278), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n229), .B(new_n260), .C1(new_n275), .C2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT25), .B1(new_n276), .B2(KEYINPUT64), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n274), .A2(new_n262), .A3(new_n265), .A4(new_n267), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n273), .A2(KEYINPUT64), .A3(KEYINPUT25), .A4(new_n274), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n229), .B1(new_n286), .B2(new_n260), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G227gat), .ZN(new_n289));
  INV_X1    g088(.A(G233gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n202), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n291), .ZN(new_n293));
  NOR4_X1   g092(.A1(new_n281), .A2(new_n287), .A3(KEYINPUT71), .A4(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT32), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT33), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n296), .B1(new_n292), .B2(new_n294), .ZN(new_n297));
  XOR2_X1   g096(.A(G15gat), .B(G43gat), .Z(new_n298));
  XNOR2_X1  g097(.A(G71gat), .B(G99gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n295), .A2(new_n297), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n300), .ZN(new_n302));
  OAI221_X1 g101(.A(KEYINPUT32), .B1(new_n296), .B2(new_n302), .C1(new_n292), .C2(new_n294), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT72), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT34), .ZN(new_n306));
  INV_X1    g105(.A(new_n287), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(new_n280), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n306), .B1(new_n308), .B2(new_n293), .ZN(new_n309));
  NOR3_X1   g108(.A1(new_n288), .A2(KEYINPUT34), .A3(new_n291), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n305), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n311), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n304), .A2(KEYINPUT72), .A3(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G78gat), .B(G106gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n315), .B(G22gat), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT2), .ZN(new_n319));
  INV_X1    g118(.A(G148gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n320), .A2(KEYINPUT76), .A3(G141gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n318), .ZN(new_n322));
  NOR2_X1   g121(.A1(G155gat), .A2(G162gat), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n319), .B(new_n321), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n320), .A2(G141gat), .ZN(new_n325));
  INV_X1    g124(.A(G141gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(G148gat), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT76), .ZN(new_n328));
  AND3_X1   g127(.A1(new_n325), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT77), .B1(new_n324), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n323), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n318), .B1(new_n331), .B2(KEYINPUT2), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n325), .A2(new_n327), .A3(new_n328), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n332), .A2(new_n333), .A3(new_n334), .A4(new_n321), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n325), .A2(new_n327), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT75), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT75), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n325), .A2(new_n327), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n338), .A2(new_n319), .A3(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n322), .A2(new_n323), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n336), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G197gat), .B(G204gat), .ZN(new_n345));
  INV_X1    g144(.A(G211gat), .ZN(new_n346));
  INV_X1    g145(.A(G218gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n345), .B1(KEYINPUT22), .B2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G211gat), .B(G218gat), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n350), .B(new_n345), .C1(KEYINPUT22), .C2(new_n348), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT29), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n344), .B1(KEYINPUT3), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT79), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT73), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n352), .A2(new_n357), .A3(new_n353), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n349), .A2(KEYINPUT73), .A3(new_n351), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT3), .ZN(new_n361));
  AND3_X1   g160(.A1(new_n336), .A2(new_n361), .A3(new_n343), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n360), .B1(new_n362), .B2(KEYINPUT29), .ZN(new_n363));
  NAND2_X1  g162(.A1(G228gat), .A2(G233gat), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT79), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n344), .B(new_n365), .C1(KEYINPUT3), .C2(new_n354), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n356), .A2(new_n363), .A3(new_n364), .A4(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n364), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n358), .A2(new_n359), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n330), .A2(new_n335), .B1(new_n341), .B2(new_n342), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n361), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n369), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n358), .A2(new_n372), .A3(new_n359), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n370), .B1(new_n374), .B2(new_n361), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n368), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT31), .B(G50gat), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n367), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n378), .B1(new_n367), .B2(new_n376), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n317), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n367), .A2(new_n376), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n377), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n376), .A3(new_n378), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(new_n316), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n312), .A2(new_n314), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT78), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT6), .ZN(new_n390));
  XNOR2_X1  g189(.A(G1gat), .B(G29gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n391), .B(KEYINPUT0), .ZN(new_n392));
  XNOR2_X1  g191(.A(G57gat), .B(G85gat), .ZN(new_n393));
  XOR2_X1   g192(.A(new_n392), .B(new_n393), .Z(new_n394));
  NAND2_X1  g193(.A1(G225gat), .A2(G233gat), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n215), .A2(new_n228), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n336), .A2(new_n343), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n370), .A2(new_n397), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n396), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT4), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n370), .A2(KEYINPUT4), .A3(new_n397), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n229), .B1(new_n370), .B2(new_n361), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n403), .B(new_n404), .C1(new_n405), .C2(new_n362), .ZN(new_n406));
  OAI211_X1 g205(.A(KEYINPUT5), .B(new_n401), .C1(new_n406), .C2(new_n396), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n403), .A2(new_n404), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT5), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n344), .A2(KEYINPUT3), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n410), .A2(new_n371), .A3(new_n229), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n408), .A2(new_n409), .A3(new_n395), .A4(new_n411), .ZN(new_n412));
  AOI211_X1 g211(.A(new_n390), .B(new_n394), .C1(new_n407), .C2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n407), .A2(new_n412), .ZN(new_n414));
  INV_X1    g213(.A(new_n394), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT6), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n407), .A2(new_n394), .A3(new_n412), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n413), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n260), .B1(new_n275), .B2(new_n279), .ZN(new_n419));
  NAND2_X1  g218(.A1(G226gat), .A2(G233gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n372), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n260), .B(new_n420), .C1(new_n275), .C2(new_n279), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n422), .A2(new_n369), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n369), .B1(new_n422), .B2(new_n423), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT74), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G8gat), .B(G36gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(G64gat), .B(G92gat), .ZN(new_n428));
  XOR2_X1   g227(.A(new_n427), .B(new_n428), .Z(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n423), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n286), .A2(new_n260), .B1(new_n372), .B2(new_n420), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n360), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT74), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n422), .A2(new_n369), .A3(new_n423), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n426), .A2(new_n430), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n433), .A2(new_n435), .A3(new_n429), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT30), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n433), .A2(KEYINPUT30), .A3(new_n435), .A4(new_n429), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n437), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n389), .B1(new_n418), .B2(new_n442), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n426), .A2(new_n430), .A3(new_n436), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n440), .A2(new_n441), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n417), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n394), .B1(new_n407), .B2(new_n412), .ZN(new_n448));
  NOR3_X1   g247(.A1(new_n447), .A2(new_n448), .A3(KEYINPUT6), .ZN(new_n449));
  OAI211_X1 g248(.A(KEYINPUT78), .B(new_n446), .C1(new_n449), .C2(new_n413), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n443), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT35), .B1(new_n388), .B2(new_n451), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n442), .A2(KEYINPUT35), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n301), .A2(new_n313), .A3(new_n303), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n313), .B1(new_n301), .B2(new_n303), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n387), .B(new_n453), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n414), .A2(KEYINPUT6), .A3(new_n415), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT83), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT83), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n448), .A2(new_n460), .A3(KEYINPUT6), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n416), .A2(new_n417), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT81), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT81), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n416), .A2(new_n465), .A3(new_n417), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n462), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  OR2_X1    g266(.A1(new_n457), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT80), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n386), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n381), .A2(new_n385), .A3(KEYINPUT80), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n448), .A2(new_n460), .A3(KEYINPUT6), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n460), .B1(new_n448), .B2(KEYINPUT6), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT38), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n426), .A2(KEYINPUT37), .A3(new_n436), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT37), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n433), .A2(new_n479), .A3(new_n435), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n480), .A2(new_n430), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n477), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT37), .B1(new_n435), .B2(KEYINPUT82), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n424), .A2(new_n425), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n483), .B1(new_n484), .B2(KEYINPUT82), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n480), .A2(new_n477), .A3(new_n430), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n438), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n482), .A2(new_n487), .ZN(new_n488));
  NOR4_X1   g287(.A1(new_n447), .A2(new_n448), .A3(KEYINPUT81), .A4(KEYINPUT6), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n465), .B1(new_n416), .B2(new_n417), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n476), .B(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n448), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n442), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT39), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n399), .A2(new_n400), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n495), .B1(new_n496), .B2(new_n395), .ZN(new_n497));
  INV_X1    g296(.A(new_n406), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n497), .B1(new_n498), .B2(new_n395), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n406), .A2(new_n495), .A3(new_n396), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(new_n394), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT40), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n499), .A2(KEYINPUT40), .A3(new_n394), .A4(new_n500), .ZN(new_n504));
  AND2_X1   g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n386), .B1(new_n494), .B2(new_n505), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n451), .A2(new_n473), .B1(new_n491), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n304), .A2(new_n311), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT36), .B1(new_n508), .B2(new_n454), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n312), .A2(new_n314), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n509), .B1(new_n510), .B2(KEYINPUT36), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n452), .A2(new_n468), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(G232gat), .A2(G233gat), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n513), .B(KEYINPUT93), .Z(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n515), .A2(KEYINPUT41), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(KEYINPUT94), .ZN(new_n517));
  XOR2_X1   g316(.A(G134gat), .B(G162gat), .Z(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT100), .ZN(new_n520));
  XOR2_X1   g319(.A(KEYINPUT86), .B(G29gat), .Z(new_n521));
  INV_X1    g320(.A(KEYINPUT87), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(new_n522), .A3(G36gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT86), .B(G29gat), .ZN(new_n524));
  INV_X1    g323(.A(G36gat), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT87), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT14), .ZN(new_n527));
  NOR2_X1   g326(.A1(G29gat), .A2(G36gat), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n527), .B1(new_n528), .B2(KEYINPUT85), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n529), .B1(KEYINPUT85), .B2(new_n528), .ZN(new_n530));
  OR3_X1    g329(.A1(new_n528), .A2(KEYINPUT85), .A3(KEYINPUT14), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n523), .A2(new_n526), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT15), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n528), .A2(KEYINPUT85), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n529), .B(new_n535), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n536), .A2(KEYINPUT15), .A3(new_n523), .A4(new_n526), .ZN(new_n537));
  XNOR2_X1  g336(.A(G43gat), .B(G50gat), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n534), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  OR3_X1    g338(.A1(new_n532), .A2(new_n533), .A3(new_n538), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT17), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT17), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n539), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(G85gat), .ZN(new_n546));
  INV_X1    g345(.A(G92gat), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT95), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT7), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n548), .B(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT8), .ZN(new_n552));
  NAND2_X1  g351(.A1(G99gat), .A2(G106gat), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n552), .B1(new_n553), .B2(KEYINPUT96), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n554), .B1(KEYINPUT96), .B2(new_n553), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT97), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n546), .A2(new_n547), .ZN(new_n557));
  AND3_X1   g356(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n556), .B1(new_n555), .B2(new_n557), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n551), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(G99gat), .B(G106gat), .Z(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n561), .B(new_n551), .C1(new_n558), .C2(new_n559), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT98), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n563), .A2(KEYINPUT98), .A3(new_n564), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n545), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n567), .A2(new_n568), .A3(new_n541), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n515), .A2(KEYINPUT41), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT99), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT99), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n570), .A2(new_n575), .A3(new_n571), .A4(new_n572), .ZN(new_n576));
  XNOR2_X1  g375(.A(G190gat), .B(G218gat), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  AND3_X1   g377(.A1(new_n574), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n578), .B1(new_n574), .B2(new_n576), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n520), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n574), .A2(new_n576), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(new_n577), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n574), .A2(new_n576), .A3(new_n578), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n519), .B(KEYINPUT100), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(G57gat), .B(G64gat), .Z(new_n588));
  XNOR2_X1  g387(.A(G71gat), .B(G78gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(G71gat), .A2(G78gat), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT9), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AND3_X1   g391(.A1(new_n588), .A2(new_n589), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n589), .B1(new_n588), .B2(new_n592), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT90), .ZN(new_n596));
  XOR2_X1   g395(.A(KEYINPUT91), .B(KEYINPUT21), .Z(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G127gat), .B(G155gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(G8gat), .ZN(new_n601));
  INV_X1    g400(.A(G1gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT16), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT88), .ZN(new_n604));
  XNOR2_X1  g403(.A(G15gat), .B(G22gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT89), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n601), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n606), .B1(G1gat), .B2(new_n605), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT21), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n611), .B1(new_n612), .B2(new_n596), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n600), .B(new_n613), .Z(new_n614));
  NAND2_X1  g413(.A1(G231gat), .A2(G233gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT92), .ZN(new_n616));
  XOR2_X1   g415(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G183gat), .B(G211gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n614), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n587), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n512), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G113gat), .B(G141gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(G169gat), .B(G197gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n610), .A2(new_n541), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n632), .B1(new_n545), .B2(new_n611), .ZN(new_n633));
  NAND2_X1  g432(.A1(G229gat), .A2(G233gat), .ZN(new_n634));
  AOI21_X1  g433(.A(KEYINPUT18), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n544), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n543), .B1(new_n539), .B2(new_n540), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n611), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n638), .A2(KEYINPUT18), .A3(new_n634), .A4(new_n631), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n634), .B(KEYINPUT13), .Z(new_n640));
  NOR2_X1   g439(.A1(new_n610), .A2(new_n541), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n640), .B1(new_n632), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n630), .B1(new_n635), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n638), .A2(new_n634), .A3(new_n631), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT18), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n647), .A2(new_n642), .A3(new_n639), .A4(new_n629), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(G120gat), .B(G148gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(G176gat), .B(G204gat), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n650), .B(new_n651), .Z(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(G230gat), .A2(G233gat), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT101), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n560), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(new_n562), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n560), .A2(new_n656), .A3(new_n561), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n658), .A2(new_n595), .A3(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT10), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n596), .A2(new_n563), .A3(new_n564), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n596), .A2(new_n661), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n567), .A2(new_n664), .A3(new_n568), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n655), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n654), .B1(new_n660), .B2(new_n662), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n653), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n663), .A2(new_n665), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n654), .ZN(new_n670));
  INV_X1    g469(.A(new_n667), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n670), .A2(new_n671), .A3(new_n652), .ZN(new_n672));
  AND3_X1   g471(.A1(new_n649), .A2(new_n668), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n623), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n418), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(new_n602), .ZN(G1324gat));
  INV_X1    g476(.A(new_n674), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT16), .B(G8gat), .Z(new_n679));
  NAND3_X1  g478(.A1(new_n678), .A2(new_n442), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT42), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n680), .A2(KEYINPUT102), .A3(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT102), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n601), .B1(new_n678), .B2(new_n442), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n680), .B1(new_n686), .B2(new_n681), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n682), .B1(new_n685), .B2(new_n687), .ZN(G1325gat));
  INV_X1    g487(.A(G15gat), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n674), .A2(new_n689), .A3(new_n511), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n508), .A2(new_n454), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n689), .B1(new_n674), .B2(new_n692), .ZN(new_n693));
  OR2_X1    g492(.A1(new_n693), .A2(KEYINPUT103), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(KEYINPUT103), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n690), .B1(new_n694), .B2(new_n695), .ZN(G1326gat));
  OR3_X1    g495(.A1(new_n674), .A2(KEYINPUT104), .A3(new_n472), .ZN(new_n697));
  OAI21_X1  g496(.A(KEYINPUT104), .B1(new_n674), .B2(new_n472), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT43), .B(G22gat), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1327gat));
  NAND2_X1  g500(.A1(new_n452), .A2(new_n468), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n507), .A2(new_n511), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n587), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n621), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n705), .A2(new_n673), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n708), .A2(new_n418), .A3(new_n524), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT45), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n711), .B1(new_n512), .B2(new_n587), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n581), .A2(new_n586), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT36), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n691), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n313), .B1(new_n304), .B2(KEYINPUT72), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT72), .ZN(new_n717));
  AOI211_X1 g516(.A(new_n717), .B(new_n311), .C1(new_n301), .C2(new_n303), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n715), .B1(new_n719), .B2(new_n714), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n503), .A2(new_n504), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n387), .B1(new_n493), .B2(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n722), .B1(new_n467), .B2(new_n488), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n472), .B1(new_n443), .B2(new_n450), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n720), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n457), .A2(new_n467), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n719), .A2(new_n387), .A3(new_n443), .A4(new_n450), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n726), .B1(new_n727), .B2(KEYINPUT35), .ZN(new_n728));
  OAI211_X1 g527(.A(KEYINPUT44), .B(new_n713), .C1(new_n725), .C2(new_n728), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n712), .A2(new_n729), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n730), .A2(new_n706), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n731), .A2(new_n418), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n710), .B1(new_n732), .B2(new_n524), .ZN(G1328gat));
  NOR3_X1   g532(.A1(new_n707), .A2(G36gat), .A3(new_n446), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT46), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n731), .A2(new_n442), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n735), .B1(new_n736), .B2(new_n525), .ZN(G1329gat));
  INV_X1    g536(.A(KEYINPUT105), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n692), .A2(G43gat), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n704), .A2(new_n706), .A3(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT106), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n712), .A2(new_n720), .A3(new_n706), .A4(new_n729), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(G43gat), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n738), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT47), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1330gat));
  INV_X1    g546(.A(G50gat), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n748), .B1(new_n731), .B2(new_n386), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n473), .A2(new_n748), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT107), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n750), .B1(new_n708), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n707), .A2(KEYINPUT107), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(KEYINPUT48), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n730), .A2(new_n473), .A3(new_n706), .ZN(new_n756));
  AOI22_X1  g555(.A1(new_n756), .A2(G50gat), .B1(new_n752), .B2(new_n753), .ZN(new_n757));
  OAI22_X1  g556(.A1(new_n749), .A2(new_n755), .B1(new_n757), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g557(.A1(new_n672), .A2(new_n668), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n649), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n623), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n418), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(G57gat), .ZN(G1332gat));
  INV_X1    g564(.A(KEYINPUT49), .ZN(new_n766));
  INV_X1    g565(.A(G64gat), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n442), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT108), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n763), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT109), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT109), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n763), .A2(new_n772), .A3(new_n769), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n766), .A2(new_n767), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n774), .B(new_n775), .ZN(G1333gat));
  OAI21_X1  g575(.A(G71gat), .B1(new_n762), .B2(new_n511), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n692), .A2(G71gat), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n762), .B2(new_n778), .ZN(new_n779));
  XOR2_X1   g578(.A(new_n779), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g579(.A1(new_n763), .A2(new_n473), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g581(.A1(new_n675), .A2(new_n760), .A3(G85gat), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n621), .A2(new_n649), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n713), .B(new_n784), .C1(new_n725), .C2(new_n728), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n704), .A2(KEYINPUT51), .A3(new_n784), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n787), .A2(KEYINPUT111), .A3(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT111), .B1(new_n787), .B2(new_n788), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n783), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n621), .A2(new_n649), .A3(new_n760), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(KEYINPUT110), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n730), .A2(new_n418), .A3(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n791), .B1(new_n546), .B2(new_n794), .ZN(G1336gat));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n446), .A2(G92gat), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n785), .A2(new_n786), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT51), .B1(new_n704), .B2(new_n784), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n759), .B(new_n797), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n712), .A2(new_n442), .A3(new_n729), .A4(new_n793), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(G92gat), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n796), .B1(new_n803), .B2(KEYINPUT52), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n805));
  AOI211_X1 g604(.A(KEYINPUT112), .B(new_n805), .C1(new_n800), .C2(new_n802), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n760), .B1(new_n787), .B2(new_n788), .ZN(new_n807));
  AOI22_X1  g606(.A1(new_n807), .A2(new_n797), .B1(G92gat), .B2(new_n801), .ZN(new_n808));
  XNOR2_X1  g607(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT114), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AND4_X1   g609(.A1(KEYINPUT114), .A2(new_n800), .A3(new_n802), .A4(new_n809), .ZN(new_n811));
  OAI22_X1  g610(.A1(new_n804), .A2(new_n806), .B1(new_n810), .B2(new_n811), .ZN(G1337gat));
  INV_X1    g611(.A(G99gat), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n730), .A2(new_n720), .A3(new_n793), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n813), .B1(new_n814), .B2(KEYINPUT115), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n815), .B1(KEYINPUT115), .B2(new_n814), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n691), .A2(new_n813), .A3(new_n759), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(KEYINPUT116), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n818), .B1(new_n789), .B2(new_n790), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n816), .A2(new_n819), .ZN(G1338gat));
  NAND3_X1  g619(.A1(new_n730), .A2(new_n386), .A3(new_n793), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(G106gat), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n387), .A2(G106gat), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT53), .B1(new_n807), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n730), .A2(new_n473), .A3(new_n793), .ZN(new_n826));
  AOI22_X1  g625(.A1(new_n826), .A2(G106gat), .B1(new_n807), .B2(new_n823), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n825), .B1(new_n827), .B2(new_n828), .ZN(G1339gat));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n663), .A2(new_n665), .A3(new_n655), .ZN(new_n831));
  AND3_X1   g630(.A1(new_n670), .A2(KEYINPUT54), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n653), .B1(new_n670), .B2(KEYINPUT54), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n830), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n670), .A2(KEYINPUT54), .A3(new_n831), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n652), .B1(new_n666), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n835), .A2(KEYINPUT55), .A3(new_n837), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n649), .A2(new_n834), .A3(new_n672), .A4(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n633), .A2(new_n634), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n632), .A2(new_n641), .A3(new_n640), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n628), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n759), .A2(new_n648), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n587), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n842), .A2(new_n648), .A3(new_n672), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n835), .A2(KEYINPUT55), .A3(new_n837), .ZN(new_n847));
  AOI21_X1  g646(.A(KEYINPUT55), .B1(new_n835), .B2(new_n837), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n713), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n845), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n705), .ZN(new_n852));
  INV_X1    g651(.A(new_n649), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n587), .A2(new_n621), .A3(new_n853), .A4(new_n760), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n388), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n675), .A2(new_n442), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n204), .A3(new_n649), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n473), .A2(new_n692), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n855), .A2(new_n860), .A3(new_n857), .ZN(new_n861));
  OAI21_X1  g660(.A(G113gat), .B1(new_n861), .B2(new_n853), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  XOR2_X1   g662(.A(new_n863), .B(KEYINPUT117), .Z(G1340gat));
  AOI21_X1  g663(.A(G120gat), .B1(new_n858), .B2(new_n759), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n861), .A2(new_n206), .A3(new_n760), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(G1341gat));
  NAND4_X1  g666(.A1(new_n858), .A2(new_n209), .A3(new_n210), .A4(new_n621), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n209), .A2(new_n210), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n869), .B1(new_n861), .B2(new_n705), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(G1342gat));
  NAND4_X1  g670(.A1(new_n858), .A2(new_n212), .A3(new_n213), .A4(new_n713), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n872), .A2(KEYINPUT56), .ZN(new_n873));
  OAI21_X1  g672(.A(G134gat), .B1(new_n861), .B2(new_n587), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(KEYINPUT56), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(G1343gat));
  XNOR2_X1  g675(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n877), .B1(new_n832), .B2(new_n833), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n649), .A2(new_n878), .A3(new_n672), .A4(new_n838), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT118), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n843), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n759), .A2(new_n842), .A3(KEYINPUT118), .A4(new_n648), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n879), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n587), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n621), .B1(new_n884), .B2(new_n850), .ZN(new_n885));
  INV_X1    g684(.A(new_n854), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n473), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT57), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n621), .B1(new_n845), .B2(new_n850), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n889), .B(new_n386), .C1(new_n890), .C2(new_n886), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n720), .A2(new_n675), .A3(new_n442), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n888), .A2(new_n649), .A3(new_n891), .A4(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(G141gat), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n855), .A2(new_n857), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n720), .A2(new_n387), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n649), .A2(new_n326), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(KEYINPUT58), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT58), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n894), .B(new_n901), .C1(new_n897), .C2(new_n898), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(new_n902), .ZN(G1344gat));
  NAND4_X1  g702(.A1(new_n895), .A2(new_n320), .A3(new_n759), .A4(new_n896), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n892), .A2(new_n759), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n887), .A2(new_n889), .ZN(new_n907));
  OAI211_X1 g706(.A(KEYINPUT57), .B(new_n386), .C1(new_n890), .C2(new_n886), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT120), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n320), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n906), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n713), .A2(new_n849), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n913), .B1(new_n587), .B2(new_n883), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n854), .B1(new_n914), .B2(new_n621), .ZN(new_n915));
  AOI21_X1  g714(.A(KEYINPUT57), .B1(new_n915), .B2(new_n473), .ZN(new_n916));
  INV_X1    g715(.A(new_n908), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n912), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(KEYINPUT120), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n905), .B1(new_n911), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n888), .A2(new_n891), .A3(new_n892), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n921), .A2(new_n760), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n922), .A2(KEYINPUT59), .A3(new_n320), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n904), .B1(new_n920), .B2(new_n923), .ZN(G1345gat));
  NAND4_X1  g723(.A1(new_n888), .A2(new_n621), .A3(new_n891), .A4(new_n892), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(G155gat), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n705), .A2(G155gat), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n926), .B1(new_n897), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(KEYINPUT121), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT121), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n926), .B(new_n930), .C1(new_n897), .C2(new_n927), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(G1346gat));
  INV_X1    g731(.A(G162gat), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n921), .A2(new_n933), .A3(new_n587), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n895), .A2(new_n713), .A3(new_n896), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n934), .B1(new_n933), .B2(new_n935), .ZN(G1347gat));
  NOR2_X1   g735(.A1(new_n418), .A2(new_n446), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n855), .A2(new_n860), .A3(new_n937), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n938), .A2(new_n245), .A3(new_n853), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n855), .A2(new_n937), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(new_n856), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(new_n649), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n939), .B1(new_n943), .B2(new_n245), .ZN(G1348gat));
  OAI21_X1  g743(.A(G176gat), .B1(new_n938), .B2(new_n760), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n759), .A2(new_n246), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n945), .B1(new_n941), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT122), .ZN(G1349gat));
  OAI21_X1  g747(.A(G183gat), .B1(new_n938), .B2(new_n705), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n621), .A2(new_n231), .A3(new_n233), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n949), .B1(new_n941), .B2(new_n950), .ZN(new_n951));
  XNOR2_X1  g750(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n952));
  XOR2_X1   g751(.A(new_n951), .B(new_n952), .Z(G1350gat));
  NAND3_X1  g752(.A1(new_n942), .A2(new_n234), .A3(new_n713), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n940), .A2(new_n713), .A3(new_n860), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n955), .A2(new_n956), .A3(G190gat), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n956), .B1(new_n955), .B2(G190gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n954), .B1(new_n958), .B2(new_n959), .ZN(G1351gat));
  AOI21_X1  g759(.A(new_n387), .B1(new_n852), .B2(new_n854), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n511), .A2(new_n937), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  XNOR2_X1  g764(.A(KEYINPUT124), .B(G197gat), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n965), .A2(new_n649), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n962), .B1(new_n907), .B2(new_n908), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n969), .A2(new_n853), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n967), .B1(new_n970), .B2(new_n966), .ZN(G1352gat));
  OAI21_X1  g770(.A(G204gat), .B1(new_n969), .B2(new_n760), .ZN(new_n972));
  OR2_X1    g771(.A1(new_n760), .A2(G204gat), .ZN(new_n973));
  OAI21_X1  g772(.A(KEYINPUT62), .B1(new_n964), .B2(new_n973), .ZN(new_n974));
  OR3_X1    g773(.A1(new_n964), .A2(KEYINPUT62), .A3(new_n973), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n972), .A2(new_n974), .A3(new_n975), .ZN(G1353gat));
  AND4_X1   g775(.A1(new_n346), .A2(new_n961), .A3(new_n621), .A4(new_n963), .ZN(new_n977));
  XOR2_X1   g776(.A(new_n977), .B(KEYINPUT125), .Z(new_n978));
  NAND2_X1  g777(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n346), .B1(new_n968), .B2(new_n621), .ZN(new_n980));
  NOR2_X1   g779(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n981));
  INV_X1    g780(.A(new_n981), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n979), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  AOI211_X1 g782(.A(new_n346), .B(new_n981), .C1(new_n968), .C2(new_n621), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n978), .B1(new_n983), .B2(new_n984), .ZN(G1354gat));
  OAI21_X1  g784(.A(G218gat), .B1(new_n969), .B2(new_n587), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n965), .A2(new_n347), .A3(new_n713), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n986), .A2(new_n987), .ZN(G1355gat));
endmodule


