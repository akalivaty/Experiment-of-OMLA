

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753;

  AND2_X1 U365 ( .A1(n598), .A2(KEYINPUT44), .ZN(n389) );
  XNOR2_X1 U366 ( .A(KEYINPUT32), .B(n593), .ZN(n751) );
  NOR2_X1 U367 ( .A1(n662), .A2(n646), .ZN(n607) );
  XNOR2_X1 U368 ( .A(n602), .B(n601), .ZN(n662) );
  NAND2_X1 U369 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U370 ( .A1(n386), .A2(n385), .ZN(n384) );
  NOR2_X1 U371 ( .A1(n692), .A2(n691), .ZN(n553) );
  NAND2_X1 U372 ( .A1(n688), .A2(n689), .ZN(n692) );
  NAND2_X1 U373 ( .A1(n396), .A2(n689), .ZN(n546) );
  INV_X1 U374 ( .A(n536), .ZN(n678) );
  XNOR2_X1 U375 ( .A(n471), .B(n470), .ZN(n513) );
  XOR2_X1 U376 ( .A(G116), .B(G107), .Z(n489) );
  INV_X1 U377 ( .A(n473), .ZN(n508) );
  XNOR2_X2 U378 ( .A(n394), .B(n441), .ZN(n688) );
  XNOR2_X2 U379 ( .A(n520), .B(n419), .ZN(n562) );
  NOR2_X1 U380 ( .A1(n364), .A2(n749), .ZN(n613) );
  XNOR2_X1 U381 ( .A(n469), .B(n468), .ZN(n471) );
  XOR2_X1 U382 ( .A(G140), .B(G107), .Z(n525) );
  XNOR2_X1 U383 ( .A(n516), .B(n439), .ZN(n736) );
  NAND2_X1 U384 ( .A1(n426), .A2(n424), .ZN(n666) );
  AND2_X4 U385 ( .A1(n444), .A2(n619), .ZN(n719) );
  AND2_X2 U386 ( .A1(n672), .A2(n616), .ZN(n444) );
  XNOR2_X2 U387 ( .A(G119), .B(G113), .ZN(n469) );
  NOR2_X1 U388 ( .A1(G953), .A2(G237), .ZN(n494) );
  NOR2_X1 U389 ( .A1(n621), .A2(G902), .ZN(n481) );
  XNOR2_X1 U390 ( .A(n472), .B(KEYINPUT69), .ZN(n495) );
  XOR2_X1 U391 ( .A(G146), .B(G125), .Z(n516) );
  INV_X1 U392 ( .A(G137), .ZN(n362) );
  OR2_X1 U393 ( .A1(n443), .A2(n655), .ZN(n344) );
  XNOR2_X1 U394 ( .A(n589), .B(n588), .ZN(n594) );
  XNOR2_X1 U395 ( .A(n681), .B(n408), .ZN(n608) );
  XNOR2_X1 U396 ( .A(n629), .B(n628), .ZN(n631) );
  XNOR2_X1 U397 ( .A(n636), .B(n635), .ZN(n638) );
  XNOR2_X1 U398 ( .A(n485), .B(n495), .ZN(n363) );
  NAND2_X1 U399 ( .A1(n379), .A2(n378), .ZN(n485) );
  XNOR2_X1 U400 ( .A(n517), .B(n362), .ZN(n361) );
  INV_X2 U401 ( .A(G953), .ZN(n740) );
  XNOR2_X1 U402 ( .A(G131), .B(KEYINPUT70), .ZN(n472) );
  XOR2_X1 U403 ( .A(KEYINPUT4), .B(KEYINPUT64), .Z(n517) );
  NOR2_X1 U404 ( .A1(n594), .A2(n590), .ZN(n592) );
  AND2_X1 U405 ( .A1(n613), .A2(n597), .ZN(n388) );
  BUF_X2 U406 ( .A(n562), .Z(n394) );
  OR2_X2 U407 ( .A1(n673), .A2(n554), .ZN(n349) );
  NAND2_X1 U408 ( .A1(n710), .A2(n359), .ZN(n358) );
  XNOR2_X1 U409 ( .A(n410), .B(G101), .ZN(n504) );
  INV_X1 U410 ( .A(KEYINPUT68), .ZN(n410) );
  OR2_X1 U411 ( .A1(G237), .A2(G902), .ZN(n521) );
  NAND2_X1 U412 ( .A1(n356), .A2(n353), .ZN(n360) );
  AND2_X1 U413 ( .A1(n358), .A2(n357), .ZN(n356) );
  NAND2_X1 U414 ( .A1(n529), .A2(n355), .ZN(n354) );
  XOR2_X1 U415 ( .A(G140), .B(KEYINPUT10), .Z(n439) );
  INV_X1 U416 ( .A(KEYINPUT102), .ZN(n368) );
  NAND2_X1 U417 ( .A1(n435), .A2(n433), .ZN(n432) );
  NAND2_X1 U418 ( .A1(KEYINPUT89), .A2(KEYINPUT48), .ZN(n435) );
  NAND2_X1 U419 ( .A1(n434), .A2(n436), .ZN(n433) );
  AND2_X1 U420 ( .A1(n565), .A2(n429), .ZN(n425) );
  NAND2_X1 U421 ( .A1(n431), .A2(n430), .ZN(n429) );
  NAND2_X1 U422 ( .A1(KEYINPUT89), .A2(n434), .ZN(n431) );
  NAND2_X1 U423 ( .A1(n436), .A2(KEYINPUT48), .ZN(n430) );
  XOR2_X1 U424 ( .A(KEYINPUT98), .B(KEYINPUT100), .Z(n477) );
  XNOR2_X1 U425 ( .A(n411), .B(n504), .ZN(n409) );
  XNOR2_X1 U426 ( .A(n475), .B(KEYINPUT99), .ZN(n411) );
  XNOR2_X1 U427 ( .A(KEYINPUT85), .B(KEYINPUT8), .ZN(n454) );
  INV_X1 U428 ( .A(G146), .ZN(n422) );
  XNOR2_X1 U429 ( .A(n504), .B(n725), .ZN(n523) );
  XNOR2_X1 U430 ( .A(n402), .B(n401), .ZN(n691) );
  INV_X1 U431 ( .A(KEYINPUT109), .ZN(n401) );
  NAND2_X1 U432 ( .A1(n390), .A2(n547), .ZN(n402) );
  INV_X1 U433 ( .A(KEYINPUT22), .ZN(n586) );
  XNOR2_X1 U434 ( .A(n519), .B(KEYINPUT82), .ZN(n419) );
  BUF_X1 U435 ( .A(n666), .Z(n738) );
  NAND2_X1 U436 ( .A1(n413), .A2(n388), .ZN(n412) );
  XNOR2_X1 U437 ( .A(G119), .B(G128), .ZN(n450) );
  XNOR2_X1 U438 ( .A(KEYINPUT84), .B(KEYINPUT23), .ZN(n452) );
  XOR2_X1 U439 ( .A(KEYINPUT7), .B(KEYINPUT105), .Z(n483) );
  XNOR2_X1 U440 ( .A(KEYINPUT106), .B(KEYINPUT9), .ZN(n482) );
  XNOR2_X1 U441 ( .A(n404), .B(n403), .ZN(n497) );
  XNOR2_X1 U442 ( .A(KEYINPUT15), .B(G902), .ZN(n615) );
  XNOR2_X1 U443 ( .A(n407), .B(n578), .ZN(n702) );
  NOR2_X1 U444 ( .A1(n577), .A2(n600), .ZN(n407) );
  INV_X1 U445 ( .A(n608), .ZN(n577) );
  NOR2_X1 U446 ( .A1(n373), .A2(n657), .ZN(n372) );
  NAND2_X1 U447 ( .A1(n371), .A2(n370), .ZN(n369) );
  INV_X1 U448 ( .A(n603), .ZN(n370) );
  INV_X1 U449 ( .A(n600), .ZN(n371) );
  XNOR2_X1 U450 ( .A(n544), .B(KEYINPUT116), .ZN(n554) );
  AND2_X1 U451 ( .A1(n681), .A2(n541), .ZN(n542) );
  XNOR2_X1 U452 ( .A(n420), .B(KEYINPUT47), .ZN(n443) );
  NAND2_X1 U453 ( .A1(n393), .A2(n392), .ZN(n420) );
  INV_X1 U454 ( .A(KEYINPUT48), .ZN(n434) );
  INV_X1 U455 ( .A(G902), .ZN(n355) );
  NAND2_X1 U456 ( .A1(n359), .A2(G902), .ZN(n357) );
  NOR2_X1 U457 ( .A1(n598), .A2(n397), .ZN(n599) );
  NAND2_X1 U458 ( .A1(n406), .A2(n398), .ZN(n397) );
  INV_X1 U459 ( .A(KEYINPUT44), .ZN(n398) );
  XNOR2_X1 U460 ( .A(n366), .B(n365), .ZN(n364) );
  INV_X1 U461 ( .A(KEYINPUT108), .ZN(n365) );
  XNOR2_X1 U462 ( .A(n492), .B(KEYINPUT12), .ZN(n403) );
  XNOR2_X1 U463 ( .A(G113), .B(G122), .ZN(n492) );
  XNOR2_X1 U464 ( .A(n493), .B(n405), .ZN(n404) );
  XNOR2_X1 U465 ( .A(G143), .B(G104), .ZN(n493) );
  XNOR2_X1 U466 ( .A(KEYINPUT103), .B(KEYINPUT11), .ZN(n405) );
  XNOR2_X1 U467 ( .A(n507), .B(KEYINPUT80), .ZN(n399) );
  INV_X1 U468 ( .A(KEYINPUT18), .ZN(n505) );
  NAND2_X1 U469 ( .A1(G234), .A2(G237), .ZN(n445) );
  AND2_X1 U470 ( .A1(n565), .A2(n432), .ZN(n428) );
  XNOR2_X1 U471 ( .A(n360), .B(n530), .ZN(n675) );
  XNOR2_X1 U472 ( .A(n380), .B(n423), .ZN(n621) );
  XNOR2_X1 U473 ( .A(n479), .B(n513), .ZN(n423) );
  XNOR2_X1 U474 ( .A(n478), .B(n409), .ZN(n479) );
  XNOR2_X1 U475 ( .A(n515), .B(n514), .ZN(n724) );
  XNOR2_X1 U476 ( .A(n513), .B(KEYINPUT76), .ZN(n514) );
  XOR2_X1 U477 ( .A(n512), .B(KEYINPUT16), .Z(n515) );
  XNOR2_X1 U478 ( .A(n380), .B(n528), .ZN(n710) );
  XNOR2_X1 U479 ( .A(n724), .B(n416), .ZN(n627) );
  XNOR2_X1 U480 ( .A(n510), .B(n417), .ZN(n416) );
  XNOR2_X1 U481 ( .A(n518), .B(n509), .ZN(n417) );
  XNOR2_X1 U482 ( .A(n399), .B(n523), .ZN(n510) );
  NAND2_X1 U483 ( .A1(n685), .A2(n369), .ZN(n686) );
  NOR2_X1 U484 ( .A1(n548), .A2(KEYINPUT39), .ZN(n382) );
  BUF_X1 U485 ( .A(n675), .Z(n400) );
  XNOR2_X1 U486 ( .A(n352), .B(n580), .ZN(n351) );
  OR2_X1 U487 ( .A1(n702), .A2(n606), .ZN(n352) );
  INV_X1 U488 ( .A(KEYINPUT34), .ZN(n579) );
  INV_X1 U489 ( .A(n581), .ZN(n414) );
  XNOR2_X1 U490 ( .A(n587), .B(n586), .ZN(n588) );
  NOR2_X1 U491 ( .A1(n535), .A2(n534), .ZN(n538) );
  XNOR2_X1 U492 ( .A(n546), .B(n545), .ZN(n567) );
  XNOR2_X1 U493 ( .A(n500), .B(n499), .ZN(n501) );
  INV_X1 U494 ( .A(KEYINPUT6), .ZN(n408) );
  XNOR2_X1 U495 ( .A(G110), .B(G104), .ZN(n725) );
  XNOR2_X1 U496 ( .A(n736), .B(n437), .ZN(n459) );
  XNOR2_X1 U497 ( .A(n488), .B(n391), .ZN(n717) );
  NOR2_X1 U498 ( .A1(G952), .A2(n740), .ZN(n723) );
  NAND2_X1 U499 ( .A1(n374), .A2(n394), .ZN(n665) );
  XNOR2_X1 U500 ( .A(n375), .B(KEYINPUT43), .ZN(n374) );
  NAND2_X1 U501 ( .A1(n377), .A2(n376), .ZN(n375) );
  NOR2_X1 U502 ( .A1(n400), .A2(n418), .ZN(n376) );
  INV_X1 U503 ( .A(KEYINPUT42), .ZN(n348) );
  NOR2_X1 U504 ( .A1(n606), .A2(n369), .ZN(n602) );
  NOR2_X1 U505 ( .A1(n708), .A2(G953), .ZN(n709) );
  XNOR2_X1 U506 ( .A(n490), .B(n491), .ZN(n552) );
  INV_X1 U507 ( .A(n552), .ZN(n390) );
  INV_X1 U508 ( .A(n689), .ZN(n418) );
  XOR2_X1 U509 ( .A(n582), .B(KEYINPUT88), .Z(n345) );
  NOR2_X2 U510 ( .A1(n346), .A2(n344), .ZN(n560) );
  NAND2_X1 U511 ( .A1(n395), .A2(n347), .ZN(n346) );
  INV_X1 U512 ( .A(n747), .ZN(n347) );
  XNOR2_X2 U513 ( .A(n349), .B(n348), .ZN(n752) );
  XNOR2_X2 U514 ( .A(n350), .B(n345), .ZN(n750) );
  NAND2_X1 U515 ( .A1(n351), .A2(n414), .ZN(n350) );
  OR2_X1 U516 ( .A1(n710), .A2(n354), .ZN(n353) );
  INV_X1 U517 ( .A(n529), .ZN(n359) );
  NAND2_X1 U518 ( .A1(n674), .A2(n360), .ZN(n537) );
  NAND2_X1 U519 ( .A1(n543), .A2(n360), .ZN(n544) );
  XNOR2_X2 U520 ( .A(n363), .B(n361), .ZN(n737) );
  NAND2_X1 U521 ( .A1(n367), .A2(n392), .ZN(n366) );
  XNOR2_X1 U522 ( .A(n607), .B(n368), .ZN(n367) );
  NAND2_X1 U523 ( .A1(n608), .A2(n372), .ZN(n503) );
  INV_X1 U524 ( .A(n541), .ZN(n373) );
  INV_X1 U525 ( .A(n561), .ZN(n377) );
  NAND2_X1 U526 ( .A1(n473), .A2(G134), .ZN(n378) );
  NAND2_X1 U527 ( .A1(n508), .A2(n474), .ZN(n379) );
  XNOR2_X2 U528 ( .A(n737), .B(n422), .ZN(n380) );
  NAND2_X1 U529 ( .A1(n384), .A2(n381), .ZN(n563) );
  NAND2_X1 U530 ( .A1(n383), .A2(n382), .ZN(n381) );
  INV_X1 U531 ( .A(n549), .ZN(n383) );
  NAND2_X1 U532 ( .A1(n548), .A2(KEYINPUT39), .ZN(n385) );
  NAND2_X1 U533 ( .A1(n549), .A2(KEYINPUT39), .ZN(n386) );
  XNOR2_X2 U534 ( .A(n387), .B(n550), .ZN(n753) );
  NAND2_X1 U535 ( .A1(n563), .A2(n659), .ZN(n387) );
  INV_X1 U536 ( .A(G134), .ZN(n474) );
  NAND2_X1 U537 ( .A1(n427), .A2(n428), .ZN(n426) );
  NOR2_X2 U538 ( .A1(n599), .A2(n389), .ZN(n413) );
  XNOR2_X1 U539 ( .A(n511), .B(n487), .ZN(n391) );
  INV_X1 U540 ( .A(n693), .ZN(n392) );
  INV_X1 U541 ( .A(n656), .ZN(n393) );
  NAND2_X1 U542 ( .A1(n559), .A2(n558), .ZN(n395) );
  NOR2_X2 U543 ( .A1(n753), .A2(n752), .ZN(n557) );
  NOR2_X2 U544 ( .A1(n594), .A2(n400), .ZN(n611) );
  INV_X1 U545 ( .A(n562), .ZN(n396) );
  INV_X1 U546 ( .A(n547), .ZN(n551) );
  NOR2_X1 U547 ( .A1(n691), .A2(n584), .ZN(n585) );
  INV_X1 U548 ( .A(n750), .ZN(n406) );
  XNOR2_X2 U549 ( .A(n412), .B(KEYINPUT45), .ZN(n415) );
  NAND2_X1 U550 ( .A1(n415), .A2(n614), .ZN(n672) );
  NOR2_X1 U551 ( .A1(n415), .A2(KEYINPUT2), .ZN(n668) );
  NAND2_X1 U552 ( .A1(n415), .A2(n738), .ZN(n618) );
  NAND2_X1 U553 ( .A1(n415), .A2(n740), .ZN(n732) );
  NAND2_X1 U554 ( .A1(n649), .A2(n751), .ZN(n598) );
  XNOR2_X2 U555 ( .A(G122), .B(n489), .ZN(n511) );
  XNOR2_X2 U556 ( .A(G128), .B(G143), .ZN(n473) );
  XNOR2_X1 U557 ( .A(n421), .B(KEYINPUT81), .ZN(n656) );
  NOR2_X1 U558 ( .A1(n554), .A2(n567), .ZN(n421) );
  NAND2_X1 U559 ( .A1(n560), .A2(n425), .ZN(n424) );
  INV_X1 U560 ( .A(n560), .ZN(n427) );
  INV_X1 U561 ( .A(KEYINPUT89), .ZN(n436) );
  XNOR2_X2 U562 ( .A(n576), .B(KEYINPUT0), .ZN(n606) );
  XOR2_X1 U563 ( .A(n451), .B(n450), .Z(n437) );
  XOR2_X1 U564 ( .A(KEYINPUT79), .B(n461), .Z(n438) );
  AND2_X1 U565 ( .A1(G214), .A2(n494), .ZN(n440) );
  XOR2_X1 U566 ( .A(KEYINPUT38), .B(KEYINPUT77), .Z(n441) );
  XOR2_X1 U567 ( .A(KEYINPUT110), .B(n585), .Z(n442) );
  XNOR2_X1 U568 ( .A(n506), .B(n505), .ZN(n507) );
  INV_X1 U569 ( .A(KEYINPUT72), .ZN(n468) );
  INV_X1 U570 ( .A(n664), .ZN(n564) );
  XNOR2_X1 U571 ( .A(n497), .B(n496), .ZN(n498) );
  NOR2_X1 U572 ( .A1(n584), .A2(n609), .ZN(n674) );
  AND2_X1 U573 ( .A1(n665), .A2(n564), .ZN(n565) );
  XNOR2_X1 U574 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U575 ( .A(n464), .B(n463), .ZN(n536) );
  XNOR2_X1 U576 ( .A(n579), .B(KEYINPUT74), .ZN(n580) );
  XNOR2_X1 U577 ( .A(n502), .B(n501), .ZN(n547) );
  XNOR2_X1 U578 ( .A(n621), .B(n620), .ZN(n622) );
  XNOR2_X1 U579 ( .A(n445), .B(KEYINPUT14), .ZN(n446) );
  NAND2_X1 U580 ( .A1(G952), .A2(n446), .ZN(n701) );
  NOR2_X1 U581 ( .A1(G953), .A2(n701), .ZN(n572) );
  NAND2_X1 U582 ( .A1(G902), .A2(n446), .ZN(n568) );
  NOR2_X1 U583 ( .A1(G900), .A2(n568), .ZN(n447) );
  NAND2_X1 U584 ( .A1(G953), .A2(n447), .ZN(n448) );
  XNOR2_X1 U585 ( .A(KEYINPUT113), .B(n448), .ZN(n449) );
  NOR2_X1 U586 ( .A1(n572), .A2(n449), .ZN(n534) );
  XOR2_X1 U587 ( .A(G110), .B(G137), .Z(n451) );
  XNOR2_X1 U588 ( .A(n452), .B(KEYINPUT24), .ZN(n453) );
  XOR2_X1 U589 ( .A(KEYINPUT73), .B(n453), .Z(n457) );
  NAND2_X1 U590 ( .A1(n740), .A2(G234), .ZN(n455) );
  XNOR2_X1 U591 ( .A(n455), .B(n454), .ZN(n486) );
  NAND2_X1 U592 ( .A1(G221), .A2(n486), .ZN(n456) );
  XNOR2_X1 U593 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U594 ( .A(n459), .B(n458), .ZN(n721) );
  NOR2_X1 U595 ( .A1(G902), .A2(n721), .ZN(n464) );
  NAND2_X1 U596 ( .A1(G234), .A2(n615), .ZN(n460) );
  XNOR2_X1 U597 ( .A(KEYINPUT20), .B(n460), .ZN(n465) );
  NAND2_X1 U598 ( .A1(G217), .A2(n465), .ZN(n462) );
  XOR2_X1 U599 ( .A(KEYINPUT25), .B(KEYINPUT96), .Z(n461) );
  XNOR2_X1 U600 ( .A(n462), .B(n438), .ZN(n463) );
  NAND2_X1 U601 ( .A1(n465), .A2(G221), .ZN(n466) );
  XNOR2_X1 U602 ( .A(n466), .B(KEYINPUT21), .ZN(n584) );
  INV_X1 U603 ( .A(n584), .ZN(n677) );
  NAND2_X1 U604 ( .A1(n536), .A2(n677), .ZN(n467) );
  NOR2_X1 U605 ( .A1(n534), .A2(n467), .ZN(n541) );
  XOR2_X1 U606 ( .A(KEYINPUT93), .B(KEYINPUT3), .Z(n470) );
  NAND2_X1 U607 ( .A1(n494), .A2(G210), .ZN(n475) );
  XNOR2_X1 U608 ( .A(G116), .B(KEYINPUT5), .ZN(n476) );
  XNOR2_X1 U609 ( .A(n477), .B(n476), .ZN(n478) );
  INV_X1 U610 ( .A(G472), .ZN(n480) );
  XNOR2_X2 U611 ( .A(n481), .B(n480), .ZN(n681) );
  XNOR2_X1 U612 ( .A(KEYINPUT107), .B(G478), .ZN(n491) );
  XNOR2_X1 U613 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U614 ( .A(n485), .B(n484), .Z(n488) );
  NAND2_X1 U615 ( .A1(G217), .A2(n486), .ZN(n487) );
  NOR2_X1 U616 ( .A1(G902), .A2(n717), .ZN(n490) );
  XNOR2_X1 U617 ( .A(n495), .B(n440), .ZN(n496) );
  XNOR2_X1 U618 ( .A(n498), .B(n736), .ZN(n634) );
  NOR2_X1 U619 ( .A1(G902), .A2(n634), .ZN(n502) );
  XNOR2_X1 U620 ( .A(KEYINPUT104), .B(KEYINPUT13), .ZN(n500) );
  INV_X1 U621 ( .A(G475), .ZN(n499) );
  NAND2_X1 U622 ( .A1(n390), .A2(n551), .ZN(n657) );
  XNOR2_X1 U623 ( .A(KEYINPUT114), .B(n503), .ZN(n561) );
  NAND2_X1 U624 ( .A1(G224), .A2(n740), .ZN(n506) );
  XOR2_X1 U625 ( .A(n508), .B(KEYINPUT17), .Z(n509) );
  INV_X1 U626 ( .A(n511), .ZN(n512) );
  XOR2_X1 U627 ( .A(n517), .B(n516), .Z(n518) );
  NAND2_X1 U628 ( .A1(n615), .A2(n627), .ZN(n520) );
  NAND2_X1 U629 ( .A1(n521), .A2(G210), .ZN(n519) );
  NAND2_X1 U630 ( .A1(G214), .A2(n521), .ZN(n689) );
  NOR2_X1 U631 ( .A1(n561), .A2(n546), .ZN(n522) );
  XNOR2_X1 U632 ( .A(KEYINPUT36), .B(n522), .ZN(n531) );
  INV_X1 U633 ( .A(n523), .ZN(n527) );
  NAND2_X1 U634 ( .A1(G227), .A2(n740), .ZN(n524) );
  XNOR2_X1 U635 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U636 ( .A(KEYINPUT71), .B(G469), .ZN(n529) );
  XNOR2_X1 U637 ( .A(KEYINPUT1), .B(KEYINPUT66), .ZN(n530) );
  NAND2_X1 U638 ( .A1(n531), .A2(n400), .ZN(n532) );
  XNOR2_X1 U639 ( .A(n532), .B(KEYINPUT117), .ZN(n747) );
  NAND2_X1 U640 ( .A1(n552), .A2(n551), .ZN(n581) );
  NAND2_X1 U641 ( .A1(n681), .A2(n689), .ZN(n533) );
  XNOR2_X1 U642 ( .A(KEYINPUT30), .B(n533), .ZN(n535) );
  INV_X1 U643 ( .A(n678), .ZN(n609) );
  XNOR2_X1 U644 ( .A(n537), .B(KEYINPUT97), .ZN(n604) );
  NAND2_X1 U645 ( .A1(n538), .A2(n604), .ZN(n549) );
  NOR2_X1 U646 ( .A1(n394), .A2(n549), .ZN(n539) );
  XNOR2_X1 U647 ( .A(n539), .B(KEYINPUT115), .ZN(n540) );
  NOR2_X1 U648 ( .A1(n581), .A2(n540), .ZN(n655) );
  XNOR2_X1 U649 ( .A(n542), .B(KEYINPUT28), .ZN(n543) );
  XOR2_X1 U650 ( .A(KEYINPUT78), .B(KEYINPUT19), .Z(n545) );
  INV_X1 U651 ( .A(n657), .ZN(n659) );
  NAND2_X1 U652 ( .A1(n552), .A2(n547), .ZN(n651) );
  INV_X1 U653 ( .A(n651), .ZN(n661) );
  NOR2_X1 U654 ( .A1(n659), .A2(n661), .ZN(n693) );
  INV_X1 U655 ( .A(n688), .ZN(n548) );
  INV_X1 U656 ( .A(KEYINPUT40), .ZN(n550) );
  XNOR2_X1 U657 ( .A(n553), .B(KEYINPUT41), .ZN(n673) );
  INV_X1 U658 ( .A(n557), .ZN(n556) );
  INV_X1 U659 ( .A(KEYINPUT46), .ZN(n555) );
  NAND2_X1 U660 ( .A1(n556), .A2(n555), .ZN(n559) );
  NAND2_X1 U661 ( .A1(n557), .A2(KEYINPUT46), .ZN(n558) );
  AND2_X1 U662 ( .A1(n661), .A2(n563), .ZN(n664) );
  NAND2_X1 U663 ( .A1(n666), .A2(KEYINPUT2), .ZN(n566) );
  XNOR2_X1 U664 ( .A(n566), .B(KEYINPUT87), .ZN(n614) );
  INV_X1 U665 ( .A(n567), .ZN(n575) );
  NOR2_X1 U666 ( .A1(G898), .A2(n740), .ZN(n727) );
  INV_X1 U667 ( .A(n568), .ZN(n569) );
  NAND2_X1 U668 ( .A1(n727), .A2(n569), .ZN(n570) );
  XOR2_X1 U669 ( .A(KEYINPUT94), .B(n570), .Z(n571) );
  NOR2_X1 U670 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U671 ( .A(KEYINPUT95), .B(n573), .ZN(n574) );
  NAND2_X1 U672 ( .A1(n675), .A2(n674), .ZN(n600) );
  XNOR2_X1 U673 ( .A(KEYINPUT112), .B(KEYINPUT33), .ZN(n578) );
  INV_X1 U674 ( .A(KEYINPUT35), .ZN(n582) );
  NAND2_X1 U675 ( .A1(n750), .A2(KEYINPUT44), .ZN(n583) );
  XNOR2_X1 U676 ( .A(n583), .B(KEYINPUT90), .ZN(n597) );
  NOR2_X1 U677 ( .A1(n606), .A2(n442), .ZN(n589) );
  INV_X1 U678 ( .A(KEYINPUT75), .ZN(n587) );
  INV_X1 U679 ( .A(n400), .ZN(n590) );
  NOR2_X1 U680 ( .A1(n608), .A2(n678), .ZN(n591) );
  NAND2_X1 U681 ( .A1(n592), .A2(n591), .ZN(n593) );
  INV_X1 U682 ( .A(n681), .ZN(n603) );
  NAND2_X1 U683 ( .A1(n611), .A2(n603), .ZN(n595) );
  XNOR2_X1 U684 ( .A(n595), .B(KEYINPUT65), .ZN(n596) );
  NAND2_X1 U685 ( .A1(n596), .A2(n609), .ZN(n649) );
  XNOR2_X1 U686 ( .A(KEYINPUT31), .B(KEYINPUT101), .ZN(n601) );
  NAND2_X1 U687 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U688 ( .A1(n606), .A2(n605), .ZN(n646) );
  NOR2_X1 U689 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X1 U690 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U691 ( .A(KEYINPUT111), .B(n612), .ZN(n749) );
  INV_X1 U692 ( .A(n615), .ZN(n616) );
  INV_X1 U693 ( .A(KEYINPUT2), .ZN(n617) );
  NAND2_X1 U694 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U695 ( .A1(n719), .A2(G472), .ZN(n623) );
  XOR2_X1 U696 ( .A(KEYINPUT62), .B(KEYINPUT92), .Z(n620) );
  XNOR2_X1 U697 ( .A(n623), .B(n622), .ZN(n625) );
  INV_X1 U698 ( .A(n723), .ZN(n624) );
  NAND2_X1 U699 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U700 ( .A(n626), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U701 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n629) );
  XNOR2_X1 U702 ( .A(n627), .B(KEYINPUT91), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n719), .A2(G210), .ZN(n630) );
  XNOR2_X1 U704 ( .A(n631), .B(n630), .ZN(n632) );
  NOR2_X2 U705 ( .A1(n632), .A2(n723), .ZN(n633) );
  XNOR2_X1 U706 ( .A(n633), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U707 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n636) );
  XNOR2_X1 U708 ( .A(n634), .B(KEYINPUT67), .ZN(n635) );
  NAND2_X1 U709 ( .A1(n719), .A2(G475), .ZN(n637) );
  XNOR2_X1 U710 ( .A(n638), .B(n637), .ZN(n639) );
  NOR2_X2 U711 ( .A1(n639), .A2(n723), .ZN(n640) );
  XNOR2_X1 U712 ( .A(n640), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U713 ( .A1(n646), .A2(n659), .ZN(n641) );
  XNOR2_X1 U714 ( .A(n641), .B(KEYINPUT118), .ZN(n642) );
  XNOR2_X1 U715 ( .A(G104), .B(n642), .ZN(G6) );
  XOR2_X1 U716 ( .A(KEYINPUT120), .B(KEYINPUT27), .Z(n644) );
  XNOR2_X1 U717 ( .A(G107), .B(KEYINPUT26), .ZN(n643) );
  XNOR2_X1 U718 ( .A(n644), .B(n643), .ZN(n645) );
  XOR2_X1 U719 ( .A(KEYINPUT119), .B(n645), .Z(n648) );
  NAND2_X1 U720 ( .A1(n646), .A2(n661), .ZN(n647) );
  XNOR2_X1 U721 ( .A(n648), .B(n647), .ZN(G9) );
  BUF_X1 U722 ( .A(n649), .Z(n650) );
  XNOR2_X1 U723 ( .A(G110), .B(n650), .ZN(G12) );
  NOR2_X1 U724 ( .A1(n651), .A2(n656), .ZN(n653) );
  XNOR2_X1 U725 ( .A(KEYINPUT121), .B(KEYINPUT29), .ZN(n652) );
  XNOR2_X1 U726 ( .A(n653), .B(n652), .ZN(n654) );
  XOR2_X1 U727 ( .A(G128), .B(n654), .Z(G30) );
  XOR2_X1 U728 ( .A(G143), .B(n655), .Z(G45) );
  NOR2_X1 U729 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U730 ( .A(G146), .B(n658), .Z(G48) );
  NAND2_X1 U731 ( .A1(n662), .A2(n659), .ZN(n660) );
  XNOR2_X1 U732 ( .A(n660), .B(G113), .ZN(G15) );
  NAND2_X1 U733 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U734 ( .A(n663), .B(G116), .ZN(G18) );
  XOR2_X1 U735 ( .A(G134), .B(n664), .Z(G36) );
  XNOR2_X1 U736 ( .A(G140), .B(n665), .ZN(G42) );
  NOR2_X1 U737 ( .A1(n666), .A2(KEYINPUT2), .ZN(n667) );
  XNOR2_X1 U738 ( .A(n667), .B(KEYINPUT86), .ZN(n669) );
  NOR2_X1 U739 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U740 ( .A(KEYINPUT83), .B(n670), .Z(n671) );
  NAND2_X1 U741 ( .A1(n672), .A2(n671), .ZN(n707) );
  NOR2_X1 U742 ( .A1(n400), .A2(n674), .ZN(n676) );
  XOR2_X1 U743 ( .A(KEYINPUT50), .B(n676), .Z(n684) );
  NOR2_X1 U744 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U745 ( .A(KEYINPUT49), .B(n679), .Z(n680) );
  NOR2_X1 U746 ( .A1(n370), .A2(n680), .ZN(n682) );
  XNOR2_X1 U747 ( .A(KEYINPUT122), .B(n682), .ZN(n683) );
  NAND2_X1 U748 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U749 ( .A(KEYINPUT51), .B(n686), .ZN(n687) );
  NOR2_X1 U750 ( .A1(n673), .A2(n687), .ZN(n698) );
  NOR2_X1 U751 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U752 ( .A1(n691), .A2(n690), .ZN(n695) );
  NOR2_X1 U753 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U754 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U755 ( .A1(n702), .A2(n696), .ZN(n697) );
  NOR2_X1 U756 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U757 ( .A(n699), .B(KEYINPUT52), .ZN(n700) );
  NOR2_X1 U758 ( .A1(n701), .A2(n700), .ZN(n705) );
  NOR2_X1 U759 ( .A1(n673), .A2(n702), .ZN(n703) );
  XOR2_X1 U760 ( .A(KEYINPUT123), .B(n703), .Z(n704) );
  NOR2_X1 U761 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U762 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U763 ( .A(n709), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U764 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n712) );
  XNOR2_X1 U765 ( .A(n710), .B(KEYINPUT57), .ZN(n711) );
  XNOR2_X1 U766 ( .A(n712), .B(n711), .ZN(n714) );
  NAND2_X1 U767 ( .A1(n719), .A2(G469), .ZN(n713) );
  XOR2_X1 U768 ( .A(n714), .B(n713), .Z(n715) );
  NOR2_X1 U769 ( .A1(n723), .A2(n715), .ZN(G54) );
  NAND2_X1 U770 ( .A1(G478), .A2(n719), .ZN(n716) );
  XNOR2_X1 U771 ( .A(n717), .B(n716), .ZN(n718) );
  NOR2_X1 U772 ( .A1(n723), .A2(n718), .ZN(G63) );
  NAND2_X1 U773 ( .A1(G217), .A2(n719), .ZN(n720) );
  XNOR2_X1 U774 ( .A(n721), .B(n720), .ZN(n722) );
  NOR2_X1 U775 ( .A1(n723), .A2(n722), .ZN(G66) );
  XNOR2_X1 U776 ( .A(G101), .B(n724), .ZN(n726) );
  XNOR2_X1 U777 ( .A(n726), .B(n725), .ZN(n728) );
  NOR2_X1 U778 ( .A1(n728), .A2(n727), .ZN(n735) );
  NAND2_X1 U779 ( .A1(G953), .A2(G224), .ZN(n729) );
  XNOR2_X1 U780 ( .A(KEYINPUT61), .B(n729), .ZN(n730) );
  NAND2_X1 U781 ( .A1(n730), .A2(G898), .ZN(n731) );
  XNOR2_X1 U782 ( .A(n731), .B(KEYINPUT126), .ZN(n733) );
  NAND2_X1 U783 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U784 ( .A(n735), .B(n734), .ZN(G69) );
  XNOR2_X1 U785 ( .A(n737), .B(n736), .ZN(n742) );
  INV_X1 U786 ( .A(n742), .ZN(n739) );
  XNOR2_X1 U787 ( .A(n739), .B(n738), .ZN(n741) );
  NAND2_X1 U788 ( .A1(n741), .A2(n740), .ZN(n746) );
  XNOR2_X1 U789 ( .A(G227), .B(n742), .ZN(n743) );
  NAND2_X1 U790 ( .A1(n743), .A2(G900), .ZN(n744) );
  NAND2_X1 U791 ( .A1(n744), .A2(G953), .ZN(n745) );
  NAND2_X1 U792 ( .A1(n746), .A2(n745), .ZN(G72) );
  XNOR2_X1 U793 ( .A(G125), .B(n747), .ZN(n748) );
  XNOR2_X1 U794 ( .A(n748), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U795 ( .A(G101), .B(n749), .Z(G3) );
  XOR2_X1 U796 ( .A(n750), .B(G122), .Z(G24) );
  XNOR2_X1 U797 ( .A(n751), .B(G119), .ZN(G21) );
  XOR2_X1 U798 ( .A(n752), .B(G137), .Z(G39) );
  XOR2_X1 U799 ( .A(n753), .B(G131), .Z(G33) );
endmodule

