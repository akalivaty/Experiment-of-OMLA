//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 1 0 0 1 0 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994;
  NAND2_X1  g000(.A1(KEYINPUT0), .A2(G128), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(G143), .B(G146), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n190), .B1(KEYINPUT0), .B2(G128), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n188), .B1(new_n189), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT0), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  AOI21_X1  g013(.A(KEYINPUT64), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n197), .A2(new_n187), .A3(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n192), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT69), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n192), .A2(new_n201), .A3(KEYINPUT69), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G131), .ZN(new_n207));
  INV_X1    g021(.A(G134), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT65), .B1(new_n208), .B2(G137), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT11), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT11), .ZN(new_n211));
  OAI211_X1 g025(.A(KEYINPUT65), .B(new_n211), .C1(new_n208), .C2(G137), .ZN(new_n212));
  INV_X1    g026(.A(G137), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(G134), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  AND4_X1   g029(.A1(new_n207), .A2(new_n210), .A3(new_n212), .A4(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n214), .B1(new_n209), .B2(KEYINPUT11), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n207), .B1(new_n217), .B2(new_n212), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT70), .ZN(new_n219));
  NOR3_X1   g033(.A1(new_n216), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n210), .A2(new_n212), .A3(new_n215), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G131), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n217), .A2(new_n207), .A3(new_n212), .ZN(new_n223));
  AOI21_X1  g037(.A(KEYINPUT70), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n206), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n194), .A2(KEYINPUT1), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n197), .A2(new_n226), .A3(G128), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n194), .B(new_n196), .C1(KEYINPUT1), .C2(new_n199), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n213), .A2(KEYINPUT66), .A3(G134), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n231), .B1(new_n208), .B2(G137), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n215), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G131), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n229), .A2(new_n223), .A3(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n225), .A2(KEYINPUT30), .A3(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(KEYINPUT2), .A2(G113), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT68), .B(G116), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G119), .ZN(new_n241));
  NAND2_X1  g055(.A1(KEYINPUT2), .A2(G113), .ZN(new_n242));
  INV_X1    g056(.A(G119), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G116), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n239), .A2(new_n241), .A3(new_n242), .A4(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  AOI22_X1  g060(.A1(new_n239), .A2(new_n242), .B1(new_n241), .B2(new_n244), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n216), .A2(new_n218), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n235), .B1(new_n250), .B2(new_n202), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT30), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n236), .A2(new_n249), .A3(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n225), .A2(new_n248), .A3(new_n235), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g072(.A1(G237), .A2(G953), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G210), .ZN(new_n260));
  INV_X1    g074(.A(G101), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n260), .B(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n263));
  XOR2_X1   g077(.A(new_n262), .B(new_n263), .Z(new_n264));
  NAND4_X1  g078(.A1(new_n236), .A2(new_n253), .A3(new_n256), .A4(new_n249), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n258), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT31), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n219), .B1(new_n216), .B2(new_n218), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n222), .A2(KEYINPUT70), .A3(new_n223), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n268), .A2(new_n269), .B1(new_n205), .B2(new_n204), .ZN(new_n270));
  INV_X1    g084(.A(new_n235), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n272), .A2(KEYINPUT28), .A3(new_n248), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT28), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n255), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n251), .A2(new_n249), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n273), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n264), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT31), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n258), .A2(new_n280), .A3(new_n264), .A4(new_n265), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n267), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(G472), .A2(G902), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n283), .B(KEYINPUT72), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT32), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n282), .A2(KEYINPUT32), .A3(new_n284), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n249), .B1(new_n270), .B2(new_n271), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT73), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n289), .A2(new_n255), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n272), .A2(KEYINPUT73), .A3(new_n248), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n293), .A2(new_n274), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n275), .B(KEYINPUT74), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n264), .A2(KEYINPUT29), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G902), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT29), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n299), .B1(new_n277), .B2(new_n278), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n264), .B1(new_n258), .B2(new_n265), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n298), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(G472), .B1(new_n297), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n287), .A2(new_n288), .A3(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT22), .B(G137), .ZN(new_n305));
  INV_X1    g119(.A(G953), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n306), .A2(G221), .A3(G234), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n305), .B(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G140), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G125), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n311), .A2(KEYINPUT16), .ZN(new_n312));
  INV_X1    g126(.A(G125), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G140), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n311), .A2(new_n314), .A3(KEYINPUT16), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n312), .B1(new_n315), .B2(KEYINPUT78), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT78), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n311), .A2(new_n317), .A3(KEYINPUT16), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n193), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n318), .ZN(new_n320));
  XNOR2_X1  g134(.A(G125), .B(G140), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n317), .B1(new_n321), .B2(KEYINPUT16), .ZN(new_n322));
  OAI211_X1 g136(.A(G146), .B(new_n320), .C1(new_n322), .C2(new_n312), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G110), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT76), .ZN(new_n326));
  OAI211_X1 g140(.A(G119), .B(new_n199), .C1(new_n326), .C2(KEYINPUT23), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT23), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n328), .B1(new_n243), .B2(G128), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT76), .B1(new_n243), .B2(G128), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n327), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT77), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n325), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI211_X1 g147(.A(KEYINPUT77), .B(new_n327), .C1(new_n329), .C2(new_n330), .ZN(new_n334));
  OR2_X1    g148(.A1(KEYINPUT24), .A2(G110), .ZN(new_n335));
  NAND2_X1  g149(.A1(KEYINPUT24), .A2(G110), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n199), .A2(G119), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n243), .A2(G128), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(KEYINPUT75), .B1(new_n337), .B2(new_n340), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n338), .A2(new_n339), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT75), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n342), .A2(new_n343), .A3(new_n335), .A4(new_n336), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n333), .A2(new_n334), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n324), .A2(new_n345), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n325), .B(new_n327), .C1(new_n329), .C2(new_n330), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n337), .A2(new_n340), .ZN(new_n348));
  AOI22_X1  g162(.A1(new_n347), .A2(new_n348), .B1(new_n193), .B2(new_n321), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n323), .A2(new_n349), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n346), .A2(KEYINPUT79), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT79), .B1(new_n346), .B2(new_n350), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n309), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT80), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI211_X1 g169(.A(KEYINPUT80), .B(new_n309), .C1(new_n351), .C2(new_n352), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n324), .A2(new_n345), .B1(new_n323), .B2(new_n349), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT81), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n358), .A2(new_n359), .A3(new_n308), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n359), .B1(new_n358), .B2(new_n308), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n357), .A2(new_n298), .A3(new_n363), .A4(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G217), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n369), .B1(G234), .B2(new_n298), .ZN(new_n370));
  AOI211_X1 g184(.A(G902), .B(new_n362), .C1(new_n355), .C2(new_n356), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n368), .B(new_n370), .C1(new_n371), .C2(new_n364), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n370), .A2(G902), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n357), .A2(new_n363), .A3(new_n373), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(G214), .B1(G237), .B2(G902), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(G110), .B(G122), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G104), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G107), .ZN(new_n381));
  INV_X1    g195(.A(G107), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n382), .A2(KEYINPUT3), .A3(G104), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT3), .B1(new_n382), .B2(G104), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n261), .B(new_n381), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n382), .A2(G104), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT3), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n387), .B1(new_n380), .B2(G107), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n382), .A2(KEYINPUT3), .A3(G104), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n386), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT87), .ZN(new_n391));
  OAI21_X1  g205(.A(G101), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AOI211_X1 g206(.A(KEYINPUT87), .B(new_n386), .C1(new_n388), .C2(new_n389), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n385), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT4), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n381), .B1(new_n383), .B2(new_n384), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT87), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n390), .A2(new_n391), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(G101), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT4), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n248), .B1(new_n395), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n241), .A2(KEYINPUT5), .A3(new_n244), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n244), .A2(KEYINPUT5), .ZN(new_n404));
  INV_X1    g218(.A(G113), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n382), .A2(G104), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n261), .B1(new_n381), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n409), .B1(new_n390), .B2(new_n261), .ZN(new_n410));
  AND3_X1   g224(.A1(new_n407), .A2(new_n245), .A3(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n379), .B1(new_n402), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n411), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n261), .B1(new_n396), .B2(KEYINPUT87), .ZN(new_n414));
  AOI21_X1  g228(.A(KEYINPUT4), .B1(new_n414), .B2(new_n398), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n415), .B1(KEYINPUT4), .B2(new_n394), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n378), .B(new_n413), .C1(new_n416), .C2(new_n248), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n412), .A2(new_n417), .A3(KEYINPUT6), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n192), .A2(new_n201), .A3(G125), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n227), .A2(new_n313), .A3(new_n228), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n306), .A2(G224), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n421), .B(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT6), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n424), .B(new_n379), .C1(new_n402), .C2(new_n411), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n418), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n378), .B(KEYINPUT8), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n410), .B1(new_n407), .B2(new_n245), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n427), .B1(new_n411), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n422), .A2(KEYINPUT7), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n419), .A2(new_n420), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n430), .B1(new_n419), .B2(new_n420), .ZN(new_n433));
  XOR2_X1   g247(.A(new_n433), .B(KEYINPUT91), .Z(new_n434));
  NOR2_X1   g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(G902), .B1(new_n435), .B2(new_n417), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n426), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(G210), .B1(G237), .B2(G902), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n426), .A2(new_n436), .A3(new_n438), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n377), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(KEYINPUT9), .B(G234), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n443), .B(KEYINPUT83), .ZN(new_n444));
  OAI21_X1  g258(.A(G221), .B1(new_n444), .B2(G902), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n445), .B(KEYINPUT84), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n400), .B1(new_n399), .B2(new_n385), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n206), .B1(new_n447), .B2(new_n415), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n268), .A2(new_n269), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n229), .A2(KEYINPUT10), .A3(new_n410), .ZN(new_n451));
  INV_X1    g265(.A(new_n409), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n385), .A2(new_n227), .A3(new_n452), .A4(new_n228), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT10), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n448), .A2(new_n450), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n385), .A2(new_n452), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n227), .A2(new_n228), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n453), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT89), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n462), .A2(new_n463), .B1(new_n268), .B2(new_n269), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n459), .A2(new_n460), .ZN(new_n465));
  AOI22_X1  g279(.A1(new_n385), .A2(new_n452), .B1(new_n227), .B2(new_n228), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(KEYINPUT89), .ZN(new_n468));
  AOI21_X1  g282(.A(KEYINPUT12), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n222), .A2(new_n223), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(KEYINPUT12), .ZN(new_n471));
  OAI21_X1  g285(.A(KEYINPUT88), .B1(new_n467), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT88), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n462), .A2(new_n470), .A3(new_n473), .A4(KEYINPUT12), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n458), .B1(new_n469), .B2(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(G110), .B(G140), .ZN(new_n477));
  INV_X1    g291(.A(G227), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n478), .A2(G953), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n477), .B(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(KEYINPUT85), .B(KEYINPUT86), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n480), .B(new_n481), .ZN(new_n482));
  AOI22_X1  g296(.A1(new_n414), .A2(new_n398), .B1(new_n261), .B2(new_n390), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n401), .B1(new_n483), .B2(new_n400), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n456), .B1(new_n484), .B2(new_n206), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n482), .B1(new_n485), .B2(new_n450), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n448), .A2(new_n457), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n449), .ZN(new_n488));
  AOI22_X1  g302(.A1(new_n476), .A2(new_n482), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(G469), .B1(new_n489), .B2(G902), .ZN(new_n490));
  AOI211_X1 g304(.A(new_n449), .B(new_n456), .C1(new_n484), .C2(new_n206), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n450), .B1(new_n448), .B2(new_n457), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n482), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n482), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n458), .B(new_n494), .C1(new_n469), .C2(new_n475), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  XOR2_X1   g310(.A(KEYINPUT90), .B(G469), .Z(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n298), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n446), .B1(new_n490), .B2(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(G113), .B(G122), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n500), .B(new_n380), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n321), .B(new_n193), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n195), .A2(KEYINPUT92), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT92), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G143), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n259), .A2(G214), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT18), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n503), .A2(G214), .A3(new_n259), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n508), .A2(new_n207), .A3(new_n510), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n502), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n510), .ZN(new_n514));
  AOI22_X1  g328(.A1(new_n503), .A2(new_n505), .B1(new_n259), .B2(G214), .ZN(new_n515));
  OAI21_X1  g329(.A(G131), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT93), .ZN(new_n517));
  NOR3_X1   g331(.A1(new_n516), .A2(new_n517), .A3(new_n509), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n207), .B1(new_n508), .B2(new_n510), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT93), .B1(new_n519), .B2(KEYINPUT18), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n513), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT17), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n516), .A2(new_n512), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT95), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT95), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n516), .A2(new_n512), .A3(new_n525), .A4(new_n522), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n519), .A2(KEYINPUT17), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(new_n319), .A3(new_n323), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n501), .B(new_n521), .C1(new_n527), .C2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n324), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n532), .A2(new_n524), .A3(new_n528), .A4(new_n526), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n501), .B1(new_n533), .B2(new_n521), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n298), .B1(new_n531), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(G475), .ZN(new_n536));
  INV_X1    g350(.A(new_n501), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n516), .A2(new_n512), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n311), .A2(new_n314), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT19), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT19), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n321), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n540), .A2(new_n542), .A3(new_n193), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT94), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT94), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n540), .A2(new_n542), .A3(new_n545), .A4(new_n193), .ZN(new_n546));
  AND4_X1   g360(.A1(new_n323), .A2(new_n538), .A3(new_n544), .A4(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n502), .A2(new_n511), .A3(new_n512), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n517), .B1(new_n516), .B2(new_n509), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n519), .A2(KEYINPUT93), .A3(KEYINPUT18), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n537), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n530), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT96), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT20), .ZN(new_n556));
  NOR2_X1   g370(.A1(G475), .A2(G902), .ZN(new_n557));
  AOI22_X1  g371(.A1(new_n555), .A2(new_n556), .B1(new_n553), .B2(new_n557), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n553), .A2(KEYINPUT96), .A3(new_n556), .A4(new_n557), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n536), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n240), .A2(G122), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(G116), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(G122), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT97), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(new_n195), .B2(G128), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n199), .A2(KEYINPUT97), .A3(G143), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n195), .A2(G128), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G134), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n570), .A2(new_n208), .A3(new_n571), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n566), .A2(new_n382), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n562), .A2(KEYINPUT100), .A3(KEYINPUT14), .ZN(new_n576));
  INV_X1    g390(.A(new_n565), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(new_n562), .B2(KEYINPUT14), .ZN(new_n578));
  AOI21_X1  g392(.A(KEYINPUT100), .B1(new_n562), .B2(KEYINPUT14), .ZN(new_n579));
  NOR3_X1   g393(.A1(new_n576), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n575), .B1(new_n580), .B2(new_n382), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n444), .A2(new_n369), .A3(G953), .ZN(new_n582));
  INV_X1    g396(.A(new_n574), .ZN(new_n583));
  OAI21_X1  g397(.A(G107), .B1(new_n563), .B2(new_n565), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n562), .A2(new_n382), .A3(new_n577), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT13), .ZN(new_n587));
  AOI22_X1  g401(.A1(new_n568), .A2(new_n569), .B1(new_n571), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT98), .ZN(new_n589));
  OR2_X1    g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n571), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n588), .A2(new_n589), .B1(KEYINPUT13), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n208), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT99), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n586), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n588), .A2(new_n589), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n591), .A2(KEYINPUT13), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n588), .A2(new_n589), .ZN(new_n599));
  OAI21_X1  g413(.A(G134), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n600), .A2(KEYINPUT99), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n581), .B(new_n582), .C1(new_n595), .C2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n600), .A2(KEYINPUT99), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n593), .A2(new_n594), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(new_n605), .A3(new_n586), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n582), .B1(new_n606), .B2(new_n581), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n298), .B1(new_n603), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(G478), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(KEYINPUT15), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(G234), .A2(G237), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(G952), .A3(new_n306), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT21), .B(G898), .Z(new_n614));
  NAND3_X1  g428(.A1(new_n612), .A2(G902), .A3(G953), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n581), .B1(new_n595), .B2(new_n601), .ZN(new_n617));
  INV_X1    g431(.A(new_n582), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n602), .ZN(new_n620));
  INV_X1    g434(.A(new_n610), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n620), .A2(new_n298), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n611), .A2(new_n616), .A3(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n561), .A2(new_n623), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n442), .A2(new_n499), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n304), .A2(new_n375), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G101), .ZN(G3));
  AND3_X1   g441(.A1(new_n372), .A2(new_n499), .A3(new_n374), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n282), .A2(new_n298), .ZN(new_n629));
  AOI22_X1  g443(.A1(new_n629), .A2(G472), .B1(new_n282), .B2(new_n284), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n426), .A2(new_n436), .A3(new_n438), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n438), .B1(new_n426), .B2(new_n436), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n376), .B(new_n616), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT33), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n634), .B1(new_n603), .B2(new_n607), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n619), .A2(KEYINPUT33), .A3(new_n602), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n609), .A2(G902), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n608), .A2(new_n609), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n561), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n633), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n628), .A2(new_n630), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT34), .B(G104), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G6));
  NAND2_X1  g459(.A1(new_n611), .A2(new_n622), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n553), .A2(KEYINPUT20), .A3(new_n557), .ZN(new_n647));
  AOI21_X1  g461(.A(KEYINPUT20), .B1(new_n553), .B2(new_n557), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n648), .B1(G475), .B2(new_n535), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n646), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n633), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n628), .A2(new_n630), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT35), .B(G107), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  NOR2_X1   g468(.A1(new_n351), .A2(new_n352), .ZN(new_n655));
  OR2_X1    g469(.A1(new_n309), .A2(KEYINPUT36), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n373), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n372), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n625), .A2(new_n630), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT37), .B(G110), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT101), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n660), .B(new_n662), .ZN(G12));
  INV_X1    g477(.A(new_n658), .ZN(new_n664));
  INV_X1    g478(.A(new_n370), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n346), .A2(new_n350), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT79), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n358), .A2(KEYINPUT79), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(KEYINPUT80), .B1(new_n670), .B2(new_n309), .ZN(new_n671));
  INV_X1    g485(.A(new_n356), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n298), .B(new_n363), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n665), .B1(new_n673), .B2(new_n365), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n664), .B1(new_n674), .B2(new_n368), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n490), .A2(new_n498), .ZN(new_n676));
  INV_X1    g490(.A(new_n446), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n376), .B1(new_n631), .B2(new_n632), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n675), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n680), .A2(new_n304), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n613), .B1(new_n615), .B2(G900), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n650), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G128), .ZN(G30));
  NAND2_X1  g500(.A1(new_n440), .A2(new_n441), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT38), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT40), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT102), .B(KEYINPUT39), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n682), .B(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n499), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n689), .B1(new_n690), .B2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n266), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n293), .A2(new_n264), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n298), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(G472), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n287), .A2(new_n288), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n693), .A2(KEYINPUT40), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n561), .A2(new_n646), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n659), .A2(new_n377), .A3(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n695), .A2(new_n700), .A3(new_n701), .A4(new_n703), .ZN(new_n704));
  XOR2_X1   g518(.A(KEYINPUT103), .B(G143), .Z(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G45));
  NAND3_X1  g520(.A1(new_n561), .A2(new_n640), .A3(new_n682), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n681), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G146), .ZN(G48));
  INV_X1    g524(.A(G469), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n711), .B1(new_n496), .B2(new_n298), .ZN(new_n712));
  INV_X1    g526(.A(new_n497), .ZN(new_n713));
  AOI211_X1 g527(.A(G902), .B(new_n713), .C1(new_n493), .C2(new_n495), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n715), .A2(KEYINPUT104), .A3(new_n677), .ZN(new_n716));
  AOI21_X1  g530(.A(G902), .B1(new_n493), .B2(new_n495), .ZN(new_n717));
  OAI211_X1 g531(.A(new_n498), .B(new_n677), .C1(new_n711), .C2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT104), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n304), .A2(new_n375), .A3(new_n642), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT41), .B(G113), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G15));
  NAND4_X1  g538(.A1(new_n304), .A2(new_n375), .A3(new_n651), .A4(new_n721), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G116), .ZN(G18));
  NAND4_X1  g540(.A1(new_n715), .A2(new_n687), .A3(new_n376), .A4(new_n677), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n727), .A2(new_n675), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n304), .A3(new_n624), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  OAI21_X1  g544(.A(new_n278), .B1(new_n294), .B2(new_n295), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(new_n267), .A3(new_n281), .ZN(new_n732));
  AOI22_X1  g546(.A1(new_n629), .A2(G472), .B1(new_n732), .B2(new_n284), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n633), .A2(new_n702), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n733), .A2(new_n721), .A3(new_n375), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G122), .ZN(G24));
  NOR3_X1   g550(.A1(new_n727), .A2(new_n675), .A3(new_n707), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n737), .A2(KEYINPUT105), .A3(new_n733), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT105), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n679), .A2(new_n718), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n659), .A3(new_n708), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n629), .A2(G472), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n732), .A2(new_n284), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n739), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n738), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G125), .ZN(G27));
  NAND2_X1  g561(.A1(new_n287), .A2(KEYINPUT107), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(new_n288), .A3(new_n303), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n287), .A2(KEYINPUT107), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n375), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n440), .A2(new_n376), .A3(new_n441), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n678), .A2(new_n707), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT42), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n304), .A2(new_n753), .A3(new_n375), .ZN(new_n756));
  AOI21_X1  g570(.A(KEYINPUT42), .B1(new_n756), .B2(KEYINPUT106), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n757), .B1(KEYINPUT106), .B2(new_n756), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G131), .ZN(G33));
  AND2_X1   g574(.A1(new_n304), .A2(new_n375), .ZN(new_n761));
  INV_X1    g575(.A(new_n752), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n684), .A2(new_n762), .A3(new_n499), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G134), .ZN(G36));
  NAND2_X1  g579(.A1(new_n489), .A2(KEYINPUT45), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT108), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT108), .B1(new_n489), .B2(KEYINPUT45), .ZN(new_n769));
  OAI21_X1  g583(.A(G469), .B1(new_n489), .B2(KEYINPUT45), .ZN(new_n770));
  OR3_X1    g584(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(G469), .A2(G902), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT46), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n771), .A2(KEYINPUT46), .A3(new_n772), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n498), .A3(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n677), .A3(new_n692), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT109), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n630), .A2(new_n675), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n780), .B(new_n781), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n638), .A2(new_n639), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n561), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n784), .B1(new_n785), .B2(KEYINPUT43), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(KEYINPUT43), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n784), .A2(new_n785), .A3(KEYINPUT43), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n782), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT44), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n752), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n792), .A2(new_n793), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(KEYINPUT112), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT112), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n792), .A2(new_n797), .A3(new_n793), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n779), .B(new_n794), .C1(new_n796), .C2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G137), .ZN(G39));
  NAND2_X1  g614(.A1(new_n777), .A2(new_n677), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT47), .ZN(new_n802));
  INV_X1    g616(.A(new_n375), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n803), .A2(new_n708), .A3(new_n762), .ZN(new_n804));
  OR3_X1    g618(.A1(new_n802), .A2(new_n304), .A3(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G140), .ZN(G42));
  OR2_X1    g620(.A1(new_n558), .A2(new_n560), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n807), .A2(new_n808), .A3(new_n536), .A4(new_n646), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n621), .B1(new_n620), .B2(new_n298), .ZN(new_n810));
  AOI211_X1 g624(.A(G902), .B(new_n610), .C1(new_n619), .C2(new_n602), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(KEYINPUT114), .B1(new_n561), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n633), .B1(new_n809), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(new_n628), .A3(new_n630), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT115), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n815), .A2(new_n660), .A3(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n817), .A2(new_n626), .A3(new_n643), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n722), .A2(new_n725), .A3(new_n729), .A4(new_n735), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n816), .B1(new_n815), .B2(new_n660), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n304), .A2(new_n812), .A3(new_n647), .A4(new_n649), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n822), .B1(new_n641), .B2(new_n744), .ZN(new_n823));
  NOR4_X1   g637(.A1(new_n675), .A2(new_n678), .A3(new_n683), .A4(new_n752), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT52), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n680), .B(new_n304), .C1(new_n684), .C2(new_n708), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n659), .A2(new_n678), .A3(new_n683), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n679), .A2(new_n702), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(new_n700), .A3(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n746), .A2(new_n826), .A3(new_n827), .A4(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(KEYINPUT105), .B1(new_n737), .B2(new_n733), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n741), .A2(new_n744), .A3(new_n739), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n827), .B(new_n830), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT52), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n821), .A2(new_n825), .A3(new_n831), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n759), .A2(new_n764), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n838));
  OR3_X1    g652(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n838), .B1(new_n836), .B2(new_n837), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(KEYINPUT54), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n843));
  OR2_X1    g657(.A1(new_n819), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n819), .A2(new_n843), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n844), .A2(new_n835), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n818), .A2(new_n820), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n838), .B1(new_n823), .B2(new_n824), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n847), .A2(new_n831), .A3(new_n848), .ZN(new_n849));
  AOI22_X1  g663(.A1(new_n755), .A2(new_n758), .B1(new_n761), .B2(new_n763), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n846), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n840), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n842), .B1(KEYINPUT54), .B2(new_n852), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n752), .A2(new_n718), .A3(new_n613), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n855), .A2(new_n700), .A3(new_n803), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n856), .A2(KEYINPUT119), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(KEYINPUT119), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n857), .A2(new_n561), .A3(new_n640), .A4(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n790), .A2(new_n613), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n803), .A2(new_n744), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n862), .A2(new_n727), .ZN(new_n863));
  INV_X1    g677(.A(G952), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n863), .A2(new_n864), .A3(G953), .ZN(new_n865));
  AND2_X1   g679(.A1(KEYINPUT120), .A2(KEYINPUT48), .ZN(new_n866));
  NOR4_X1   g680(.A1(new_n751), .A2(new_n790), .A3(new_n855), .A4(new_n866), .ZN(new_n867));
  OR3_X1    g681(.A1(new_n867), .A2(KEYINPUT120), .A3(KEYINPUT48), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n867), .B1(KEYINPUT120), .B2(KEYINPUT48), .ZN(new_n869));
  AND4_X1   g683(.A1(new_n859), .A2(new_n865), .A3(new_n868), .A4(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT51), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n791), .A2(new_n659), .A3(new_n733), .A4(new_n854), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(KEYINPUT118), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n561), .A2(new_n640), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n857), .A2(new_n858), .A3(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n689), .A2(new_n377), .A3(new_n677), .A4(new_n715), .ZN(new_n876));
  OAI21_X1  g690(.A(KEYINPUT50), .B1(new_n862), .B2(new_n876), .ZN(new_n877));
  OR3_X1    g691(.A1(new_n862), .A2(KEYINPUT50), .A3(new_n876), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n873), .A2(new_n875), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n677), .B1(new_n715), .B2(KEYINPUT117), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n881), .B1(KEYINPUT117), .B2(new_n715), .ZN(new_n882));
  AOI211_X1 g696(.A(new_n752), .B(new_n862), .C1(new_n802), .C2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n871), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n879), .A2(new_n883), .A3(KEYINPUT51), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n870), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n853), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(G952), .A2(G953), .ZN(new_n889));
  NOR4_X1   g703(.A1(new_n783), .A2(new_n561), .A3(new_n377), .A4(new_n446), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT49), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n375), .B(new_n890), .C1(new_n891), .C2(new_n715), .ZN(new_n892));
  OR2_X1    g706(.A1(new_n892), .A2(KEYINPUT113), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(KEYINPUT113), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n715), .A2(new_n891), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n893), .A2(new_n689), .A3(new_n894), .A4(new_n895), .ZN(new_n896));
  OAI22_X1  g710(.A1(new_n888), .A2(new_n889), .B1(new_n700), .B2(new_n896), .ZN(G75));
  AOI21_X1  g711(.A(new_n298), .B1(new_n840), .B2(new_n851), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT56), .B1(new_n898), .B2(G210), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n418), .A2(new_n425), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(new_n423), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT55), .Z(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(KEYINPUT121), .B1(new_n899), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n905));
  INV_X1    g719(.A(G210), .ZN(new_n906));
  AOI211_X1 g720(.A(new_n906), .B(new_n298), .C1(new_n840), .C2(new_n851), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n905), .B(new_n902), .C1(new_n907), .C2(KEYINPUT56), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n864), .A2(G953), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT123), .Z(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  OR2_X1    g726(.A1(new_n902), .A2(KEYINPUT56), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n852), .A2(G210), .A3(G902), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT122), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n907), .A2(KEYINPUT122), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n912), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n909), .A2(new_n918), .ZN(G51));
  INV_X1    g733(.A(KEYINPUT54), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n852), .B(new_n920), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n772), .B(KEYINPUT57), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n496), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n771), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n898), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n912), .B1(new_n923), .B2(new_n925), .ZN(G54));
  INV_X1    g740(.A(new_n553), .ZN(new_n927));
  AND2_X1   g741(.A1(KEYINPUT58), .A2(G475), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n898), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n927), .B1(new_n898), .B2(new_n928), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n911), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT124), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI211_X1 g747(.A(KEYINPUT124), .B(new_n911), .C1(new_n929), .C2(new_n930), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(G60));
  AND2_X1   g749(.A1(new_n635), .A2(new_n636), .ZN(new_n936));
  NAND2_X1  g750(.A1(G478), .A2(G902), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT59), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n936), .B1(new_n853), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n936), .A2(new_n938), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n911), .B1(new_n921), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n939), .A2(new_n941), .ZN(G63));
  XNOR2_X1  g756(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n369), .A2(new_n298), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n852), .A2(new_n657), .A3(new_n945), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n852), .A2(new_n945), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n362), .B1(new_n355), .B2(new_n356), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n911), .B(new_n946), .C1(new_n947), .C2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n949), .B(new_n950), .ZN(G66));
  NAND2_X1  g765(.A1(new_n614), .A2(G224), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(G953), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(new_n821), .B2(G953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n900), .B1(G898), .B2(new_n306), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n954), .B(new_n955), .ZN(G69));
  INV_X1    g770(.A(G900), .ZN(new_n957));
  OAI21_X1  g771(.A(G953), .B1(new_n478), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n236), .A2(new_n253), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n540), .A2(new_n542), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n959), .B(new_n960), .Z(new_n961));
  AOI21_X1  g775(.A(new_n961), .B1(G900), .B2(G953), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n746), .A2(new_n827), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n375), .B(new_n829), .C1(new_n749), .C2(new_n750), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n964), .B1(new_n779), .B2(new_n966), .ZN(new_n967));
  AND4_X1   g781(.A1(new_n799), .A2(new_n967), .A3(new_n805), .A4(new_n850), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n963), .B1(new_n968), .B2(new_n306), .ZN(new_n969));
  INV_X1    g783(.A(new_n961), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n809), .A2(new_n641), .A3(new_n813), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n761), .A2(new_n694), .A3(new_n762), .A4(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n704), .A2(new_n746), .A3(new_n827), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT62), .Z(new_n974));
  NAND4_X1  g788(.A1(new_n799), .A2(new_n805), .A3(new_n972), .A4(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n970), .B1(new_n975), .B2(new_n306), .ZN(new_n976));
  OAI211_X1 g790(.A(KEYINPUT126), .B(new_n958), .C1(new_n969), .C2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n976), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n958), .A2(KEYINPUT126), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n799), .A2(new_n805), .A3(new_n850), .A4(new_n967), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n962), .B1(new_n980), .B2(G953), .ZN(new_n981));
  OR2_X1    g795(.A1(new_n958), .A2(KEYINPUT126), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n978), .A2(new_n979), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n977), .A2(new_n983), .ZN(G72));
  XNOR2_X1  g798(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n985));
  NAND2_X1  g799(.A1(G472), .A2(G902), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n985), .B(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(new_n821), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n987), .B1(new_n980), .B2(new_n988), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n989), .A2(new_n278), .A3(new_n258), .A4(new_n265), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n841), .B(new_n987), .C1(new_n696), .C2(new_n301), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n987), .B1(new_n975), .B2(new_n988), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n278), .B1(new_n258), .B2(new_n265), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AND4_X1   g808(.A1(new_n911), .A2(new_n990), .A3(new_n991), .A4(new_n994), .ZN(G57));
endmodule


