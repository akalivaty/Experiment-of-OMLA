//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 1 1 0 0 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1255, new_n1256, new_n1257, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n208), .B1(new_n211), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT1), .ZN(new_n216));
  OR3_X1    g0016(.A1(new_n208), .A2(KEYINPUT64), .A3(G13), .ZN(new_n217));
  OAI21_X1  g0017(.A(KEYINPUT64), .B1(new_n208), .B2(G13), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n219), .B(G250), .C1(G257), .C2(G264), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT0), .Z(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(G58), .A2(G68), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G50), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  AOI211_X1 g0028(.A(new_n216), .B(new_n221), .C1(new_n224), .C2(new_n228), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G226), .B(G232), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT66), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n234), .B(new_n238), .Z(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT67), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  XNOR2_X1  g0047(.A(KEYINPUT71), .B(G200), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT3), .B(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G1698), .ZN(new_n250));
  INV_X1    g0050(.A(G223), .ZN(new_n251));
  OAI22_X1  g0051(.A1(new_n250), .A2(new_n251), .B1(new_n202), .B2(new_n249), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n249), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G222), .ZN(new_n255));
  OR3_X1    g0055(.A1(new_n254), .A2(KEYINPUT68), .A3(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(KEYINPUT68), .B1(new_n254), .B2(new_n255), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n252), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G1), .A3(G13), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  INV_X1    g0062(.A(G45), .ZN(new_n263));
  AOI21_X1  g0063(.A(G1), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(new_n260), .A3(G274), .ZN(new_n265));
  INV_X1    g0065(.A(G226), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n260), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n265), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n248), .B1(new_n261), .B2(new_n270), .ZN(new_n271));
  OAI221_X1 g0071(.A(new_n265), .B1(new_n266), .B2(new_n269), .C1(new_n258), .C2(new_n260), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n271), .B1(G190), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT74), .ZN(new_n274));
  AOI21_X1  g0074(.A(KEYINPUT10), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n223), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G150), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT8), .B(G58), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n223), .A2(G33), .ZN(new_n281));
  OAI221_X1 g0081(.A(new_n279), .B1(new_n201), .B2(new_n223), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT69), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n283), .B1(new_n208), .B2(new_n276), .ZN(new_n284));
  NAND4_X1  g0084(.A1(KEYINPUT69), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(new_n222), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G50), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n267), .A2(G13), .A3(G20), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n282), .A2(new_n286), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n286), .A2(new_n289), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n267), .A2(G20), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n291), .A2(G50), .A3(new_n292), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT9), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n294), .B(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n273), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n275), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n296), .B(new_n273), .C1(new_n274), .C2(KEYINPUT10), .ZN(new_n299));
  INV_X1    g0099(.A(G169), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n294), .B1(new_n272), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n301), .B1(G179), .B2(new_n272), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n298), .A2(new_n299), .A3(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n291), .A2(G77), .A3(new_n292), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n289), .A2(new_n202), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G20), .A2(G77), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(new_n280), .B2(new_n277), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n276), .A2(G20), .ZN(new_n308));
  XNOR2_X1  g0108(.A(KEYINPUT15), .B(G87), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n307), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n286), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n304), .B(new_n305), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G244), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n265), .B1(new_n314), .B2(new_n269), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n249), .A2(G232), .A3(new_n253), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n249), .A2(G238), .A3(G1698), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n316), .B(new_n317), .C1(new_n205), .C2(new_n249), .ZN(new_n318));
  INV_X1    g0118(.A(new_n260), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n315), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G190), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n313), .B1(new_n323), .B2(KEYINPUT70), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT70), .B1(new_n320), .B2(new_n248), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(new_n322), .B2(new_n321), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n313), .B1(G169), .B2(new_n320), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT72), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT72), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n313), .B(new_n330), .C1(G169), .C2(new_n320), .ZN(new_n331));
  INV_X1    g0131(.A(G179), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n320), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n329), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n327), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g0135(.A(new_n335), .B(KEYINPUT73), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n276), .A2(KEYINPUT3), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT3), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(G33), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT7), .B1(new_n340), .B2(new_n223), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT7), .ZN(new_n342));
  AOI211_X1 g0142(.A(new_n342), .B(G20), .C1(new_n337), .C2(new_n339), .ZN(new_n343));
  OAI21_X1  g0143(.A(G68), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G58), .ZN(new_n345));
  INV_X1    g0145(.A(G68), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(G20), .B1(new_n347), .B2(new_n225), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n278), .A2(G159), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n344), .A2(KEYINPUT16), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT16), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n342), .B1(new_n249), .B2(G20), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n338), .A2(G33), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n276), .A2(KEYINPUT3), .ZN(new_n356));
  OAI211_X1 g0156(.A(KEYINPUT7), .B(new_n223), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n346), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n353), .B1(new_n358), .B2(new_n350), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n352), .A2(new_n359), .A3(new_n286), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n280), .B1(new_n267), .B2(G20), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n291), .A2(new_n361), .B1(new_n289), .B2(new_n280), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n337), .A2(new_n339), .A3(G226), .A4(G1698), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n337), .A2(new_n339), .A3(G223), .A4(new_n253), .ZN(new_n364));
  NAND2_X1  g0164(.A1(G33), .A2(G87), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n319), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n260), .A2(G232), .A3(new_n268), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n265), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n367), .A2(new_n322), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n369), .B1(new_n319), .B2(new_n366), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n371), .B1(G200), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n360), .A2(new_n362), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT77), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n360), .A2(new_n373), .A3(KEYINPUT77), .A4(new_n362), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT17), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT17), .ZN(new_n380));
  AND2_X1   g0180(.A1(new_n374), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n367), .A2(new_n332), .A3(new_n370), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(G169), .B2(new_n372), .ZN(new_n384));
  AOI211_X1 g0184(.A(KEYINPUT18), .B(new_n384), .C1(new_n360), .C2(new_n362), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT18), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n360), .A2(new_n362), .ZN(new_n387));
  INV_X1    g0187(.A(new_n384), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n379), .A2(new_n382), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n346), .A2(G20), .ZN(new_n392));
  OAI221_X1 g0192(.A(new_n392), .B1(new_n281), .B2(new_n202), .C1(new_n287), .C2(new_n277), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n286), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n394), .A2(KEYINPUT75), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(KEYINPUT75), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT11), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT11), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n395), .A2(new_n399), .A3(new_n396), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT76), .B1(new_n288), .B2(G68), .ZN(new_n401));
  XNOR2_X1  g0201(.A(new_n401), .B(KEYINPUT12), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n346), .B1(new_n267), .B2(G20), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n402), .B1(new_n291), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n398), .A2(new_n400), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT14), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n249), .A2(G232), .A3(G1698), .ZN(new_n407));
  NAND2_X1  g0207(.A1(G33), .A2(G97), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n337), .A2(new_n339), .A3(G226), .A4(new_n253), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n319), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT13), .ZN(new_n412));
  INV_X1    g0212(.A(new_n269), .ZN(new_n413));
  INV_X1    g0213(.A(G274), .ZN(new_n414));
  INV_X1    g0214(.A(new_n222), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n414), .B1(new_n415), .B2(new_n259), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n413), .A2(G238), .B1(new_n264), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n411), .A2(new_n412), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n412), .B1(new_n411), .B2(new_n417), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n406), .B(G169), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n411), .A2(new_n417), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT13), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n423), .A2(G179), .A3(new_n418), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n418), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n406), .B1(new_n426), .B2(G169), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n405), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n398), .A2(new_n400), .A3(new_n404), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n423), .A2(G190), .A3(new_n418), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n426), .A2(G200), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  NOR4_X1   g0233(.A1(new_n303), .A2(new_n336), .A3(new_n391), .A4(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n337), .A2(new_n339), .A3(G238), .A4(new_n253), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT80), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT80), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n249), .A2(new_n437), .A3(G238), .A4(new_n253), .ZN(new_n438));
  NAND2_X1  g0238(.A1(G33), .A2(G116), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n249), .A2(G244), .A3(G1698), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n436), .A2(new_n438), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n319), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n263), .A2(G1), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n416), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n267), .A2(G45), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n260), .A2(G250), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n248), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AND2_X1   g0251(.A1(KEYINPUT78), .A2(G97), .ZN(new_n452));
  NOR2_X1   g0252(.A1(KEYINPUT78), .A2(G97), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n308), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT19), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OR2_X1    g0256(.A1(KEYINPUT78), .A2(G97), .ZN(new_n457));
  NAND2_X1  g0257(.A1(KEYINPUT78), .A2(G97), .ZN(new_n458));
  NOR2_X1   g0258(.A1(G87), .A2(G107), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n223), .B1(new_n408), .B2(new_n455), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n249), .A2(new_n223), .A3(G68), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n456), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n286), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n267), .A2(G33), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n291), .A2(G87), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n309), .A2(new_n289), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n451), .A2(new_n470), .A3(KEYINPUT81), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT81), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n248), .B1(new_n442), .B2(new_n448), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n472), .B1(new_n473), .B2(new_n469), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n447), .B1(new_n441), .B2(new_n319), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G190), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n471), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n464), .A2(new_n286), .B1(new_n289), .B2(new_n309), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n291), .A2(new_n310), .A3(new_n466), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n332), .A2(new_n475), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n449), .A2(new_n300), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n337), .A2(new_n339), .A3(new_n223), .A4(G87), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT22), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT22), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n249), .A2(new_n486), .A3(new_n223), .A4(G87), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT24), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n439), .A2(G20), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT23), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(new_n223), .B2(G107), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n205), .A2(KEYINPUT23), .A3(G20), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n490), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n488), .A2(new_n489), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n489), .B1(new_n488), .B2(new_n494), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n286), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n289), .A2(new_n205), .ZN(new_n498));
  XNOR2_X1  g0298(.A(new_n498), .B(KEYINPUT25), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n285), .A2(new_n222), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n500), .A2(new_n284), .A3(new_n288), .A4(new_n466), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(new_n205), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n497), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n337), .A2(new_n339), .A3(G257), .A4(G1698), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n337), .A2(new_n339), .A3(G250), .A4(new_n253), .ZN(new_n506));
  NAND2_X1  g0306(.A1(G33), .A2(G294), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  XNOR2_X1  g0308(.A(KEYINPUT5), .B(G41), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n509), .A2(new_n443), .B1(new_n415), .B2(new_n259), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n508), .A2(new_n319), .B1(new_n510), .B2(G264), .ZN(new_n511));
  OR2_X1    g0311(.A1(KEYINPUT5), .A2(G41), .ZN(new_n512));
  NAND2_X1  g0312(.A1(KEYINPUT5), .A2(G41), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n445), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n416), .ZN(new_n515));
  AOI21_X1  g0315(.A(G169), .B1(new_n511), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n511), .A2(new_n515), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n516), .B1(new_n518), .B2(new_n332), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n504), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n278), .A2(G77), .ZN(new_n521));
  NAND2_X1  g0321(.A1(G97), .A2(G107), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT6), .B1(new_n206), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n457), .A2(new_n458), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT6), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n525), .A2(G107), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n523), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n521), .B1(new_n527), .B2(new_n223), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n205), .B1(new_n354), .B2(new_n357), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n286), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n291), .A2(G97), .A3(new_n466), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n289), .A2(new_n204), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n513), .ZN(new_n534));
  NOR2_X1   g0334(.A1(KEYINPUT5), .A2(G41), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n443), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n536), .A2(G257), .A3(new_n260), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n515), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n337), .A2(new_n339), .A3(G244), .A4(new_n253), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT4), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n249), .A2(KEYINPUT4), .A3(G244), .A4(new_n253), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G283), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n337), .A2(new_n339), .A3(G250), .A4(G1698), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n541), .A2(new_n542), .A3(new_n543), .A4(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n538), .B1(new_n545), .B2(new_n319), .ZN(new_n546));
  OR2_X1    g0346(.A1(new_n546), .A2(G169), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT79), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n537), .A2(new_n515), .A3(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n548), .B1(new_n537), .B2(new_n515), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n543), .B(new_n544), .C1(new_n539), .C2(new_n540), .ZN(new_n553));
  AND2_X1   g0353(.A1(new_n539), .A2(new_n540), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n319), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n552), .A2(new_n332), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n533), .A2(new_n547), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n538), .A2(KEYINPUT79), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n555), .A2(new_n558), .A3(new_n549), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(G200), .ZN(new_n560));
  OAI21_X1  g0360(.A(G107), .B1(new_n341), .B2(new_n343), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n524), .A2(new_n526), .ZN(new_n562));
  INV_X1    g0362(.A(new_n522), .ZN(new_n563));
  NOR2_X1   g0363(.A1(G97), .A2(G107), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n525), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G20), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n561), .A2(new_n567), .A3(new_n521), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n568), .A2(new_n286), .B1(new_n204), .B2(new_n289), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n546), .A2(G190), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n560), .A2(new_n569), .A3(new_n531), .A4(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n517), .A2(G190), .ZN(new_n572));
  AOI21_X1  g0372(.A(G200), .B1(new_n511), .B2(new_n515), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n497), .B(new_n503), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n520), .A2(new_n557), .A3(new_n571), .A4(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n288), .A2(G116), .ZN(new_n576));
  INV_X1    g0376(.A(G116), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(G20), .ZN(new_n578));
  AOI21_X1  g0378(.A(G33), .B1(new_n457), .B2(new_n458), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n543), .A2(new_n223), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n286), .B(new_n578), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  XOR2_X1   g0381(.A(KEYINPUT83), .B(KEYINPUT20), .Z(new_n582));
  AOI21_X1  g0382(.A(new_n576), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n291), .A2(KEYINPUT82), .A3(G116), .A4(new_n466), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT82), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n501), .B2(new_n577), .ZN(new_n586));
  OR2_X1    g0386(.A1(new_n579), .A2(new_n580), .ZN(new_n587));
  NOR2_X1   g0387(.A1(KEYINPUT83), .A2(KEYINPUT20), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n587), .A2(new_n286), .A3(new_n578), .A4(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n583), .A2(new_n584), .A3(new_n586), .A4(new_n589), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n510), .A2(G270), .B1(new_n416), .B2(new_n514), .ZN(new_n591));
  OAI21_X1  g0391(.A(G303), .B1(new_n355), .B2(new_n356), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n337), .A2(new_n339), .A3(G264), .A4(G1698), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n337), .A2(new_n339), .A3(G257), .A4(new_n253), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n319), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n300), .B1(new_n591), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n590), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT84), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n599), .A2(KEYINPUT21), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n583), .A2(new_n586), .A3(new_n589), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n591), .A2(new_n596), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(G200), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n591), .A2(new_n596), .A3(G190), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n602), .A2(new_n584), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n591), .A2(new_n596), .A3(G179), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n590), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n600), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n590), .A2(new_n597), .A3(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n601), .A2(new_n606), .A3(new_n609), .A4(new_n611), .ZN(new_n612));
  NOR3_X1   g0412(.A1(new_n483), .A2(new_n575), .A3(new_n612), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n434), .A2(new_n613), .ZN(G372));
  NAND2_X1  g0414(.A1(new_n469), .A2(KEYINPUT85), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT85), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n478), .A2(new_n616), .A3(new_n467), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  AOI211_X1 g0418(.A(new_n322), .B(new_n447), .C1(new_n441), .C2(new_n319), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n473), .A2(new_n619), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n618), .A2(new_n620), .B1(new_n481), .B2(new_n480), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n621), .A2(new_n574), .A3(new_n557), .A4(new_n571), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT86), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n611), .A2(new_n609), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n610), .B1(new_n590), .B2(new_n597), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n601), .A2(KEYINPUT86), .A3(new_n609), .A4(new_n611), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n622), .B1(new_n628), .B2(new_n520), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT26), .ZN(new_n630));
  AND4_X1   g0430(.A1(new_n616), .A2(new_n465), .A3(new_n468), .A4(new_n467), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n616), .B1(new_n478), .B2(new_n467), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n476), .B1(new_n248), .B2(new_n475), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n482), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n630), .B1(new_n635), .B2(new_n557), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n533), .A2(new_n547), .A3(new_n556), .ZN(new_n637));
  XOR2_X1   g0437(.A(KEYINPUT87), .B(KEYINPUT26), .Z(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n477), .A2(new_n637), .A3(new_n482), .A4(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n482), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n434), .B1(new_n629), .B2(new_n642), .ZN(new_n643));
  XOR2_X1   g0443(.A(new_n643), .B(KEYINPUT88), .Z(new_n644));
  INV_X1    g0444(.A(new_n432), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n428), .B1(new_n645), .B2(new_n334), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n381), .B1(new_n378), .B2(KEYINPUT17), .ZN(new_n647));
  AOI211_X1 g0447(.A(new_n389), .B(new_n385), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n298), .A2(new_n299), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n302), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n644), .A2(new_n650), .ZN(G369));
  INV_X1    g0451(.A(G330), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n612), .A2(KEYINPUT89), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n612), .A2(KEYINPUT89), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n267), .A2(new_n223), .A3(G13), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(G213), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(G343), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n590), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n655), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT90), .ZN(new_n664));
  INV_X1    g0464(.A(new_n662), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n628), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n663), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n665), .B1(new_n653), .B2(new_n654), .ZN(new_n668));
  INV_X1    g0468(.A(new_n666), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT90), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n652), .B1(new_n667), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n504), .A2(new_n661), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n574), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n673), .A2(new_n520), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n520), .A2(new_n661), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n661), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n624), .B2(new_n625), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n673), .A2(new_n520), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n675), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n677), .A2(new_n682), .ZN(G399));
  INV_X1    g0483(.A(new_n219), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(G41), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n460), .A2(G116), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n685), .A2(new_n267), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n688), .B1(new_n228), .B2(new_n685), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT28), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT93), .ZN(new_n691));
  INV_X1    g0491(.A(new_n629), .ZN(new_n692));
  INV_X1    g0492(.A(new_n482), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n693), .B1(new_n636), .B2(new_n640), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n661), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n691), .B1(new_n695), .B2(KEYINPUT29), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n678), .B1(new_n642), .B2(new_n629), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT29), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(KEYINPUT93), .A3(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n557), .A2(new_n571), .A3(new_n574), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(new_n635), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n520), .A2(new_n601), .A3(new_n609), .A4(new_n611), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n693), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n477), .A2(new_n637), .A3(new_n482), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n638), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n621), .A2(new_n637), .A3(KEYINPUT26), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n708), .A2(KEYINPUT29), .A3(new_n678), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(KEYINPUT94), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n661), .B1(new_n703), .B2(new_n707), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT94), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(new_n712), .A3(KEYINPUT29), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n696), .A2(new_n699), .B1(new_n710), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n538), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n555), .A2(new_n511), .A3(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT91), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n607), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n591), .A2(new_n596), .A3(KEYINPUT91), .A4(G179), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n716), .A2(new_n718), .A3(new_n475), .A4(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT30), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n517), .A2(new_n332), .A3(new_n603), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n475), .B1(new_n552), .B2(new_n555), .ZN(new_n723));
  AOI22_X1  g0523(.A1(new_n720), .A2(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT92), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(new_n720), .B2(new_n721), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n718), .A2(new_n719), .ZN(new_n727));
  AND3_X1   g0527(.A1(new_n546), .A2(new_n475), .A3(new_n511), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n727), .A2(KEYINPUT92), .A3(KEYINPUT30), .A4(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n724), .A2(new_n726), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(new_n661), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT31), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n575), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n477), .A2(new_n482), .ZN(new_n735));
  INV_X1    g0535(.A(new_n612), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n734), .A2(new_n735), .A3(new_n736), .A4(new_n678), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n730), .A2(KEYINPUT31), .A3(new_n661), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n733), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G330), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n714), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n690), .B1(new_n743), .B2(new_n267), .ZN(new_n744));
  XOR2_X1   g0544(.A(new_n744), .B(KEYINPUT95), .Z(G364));
  INV_X1    g0545(.A(new_n670), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n668), .A2(new_n669), .A3(KEYINPUT90), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G13), .A2(G33), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  AND2_X1   g0552(.A1(new_n223), .A2(G13), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n267), .B1(new_n753), .B2(G45), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n685), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n223), .A2(G179), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n450), .A2(new_n322), .A3(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT98), .ZN(new_n759));
  OR2_X1    g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G283), .ZN(new_n764));
  NOR4_X1   g0564(.A1(new_n223), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n249), .B1(new_n765), .B2(G329), .ZN(new_n766));
  INV_X1    g0566(.A(G294), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n322), .A2(G179), .A3(G200), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n223), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n766), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(G20), .A2(G179), .ZN(new_n771));
  XOR2_X1   g0571(.A(new_n771), .B(KEYINPUT96), .Z(new_n772));
  NOR2_X1   g0572(.A1(G190), .A2(G200), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n770), .B1(new_n775), .B2(G311), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n322), .A2(G200), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n772), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n450), .A2(G190), .A3(new_n757), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n779), .A2(G322), .B1(new_n781), .B2(G303), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n772), .A2(G200), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n322), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(G190), .ZN(new_n785));
  XNOR2_X1  g0585(.A(KEYINPUT33), .B(G317), .ZN(new_n786));
  AOI22_X1  g0586(.A1(G326), .A2(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n764), .A2(new_n776), .A3(new_n782), .A4(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n785), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n789), .A2(new_n346), .B1(new_n204), .B2(new_n769), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n790), .A2(KEYINPUT99), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(KEYINPUT99), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n762), .A2(new_n205), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n765), .A2(G159), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT32), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n340), .B(new_n796), .C1(G87), .C2(new_n781), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n791), .A2(new_n792), .A3(new_n794), .A4(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(G58), .A2(new_n779), .B1(new_n775), .B2(G77), .ZN(new_n799));
  INV_X1    g0599(.A(new_n784), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n799), .B1(new_n287), .B2(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT97), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n788), .B1(new_n798), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n222), .B1(G20), .B2(new_n300), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n751), .A2(new_n804), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n684), .A2(new_n249), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(G45), .B2(new_n227), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(G45), .B2(new_n242), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n219), .A2(new_n249), .ZN(new_n810));
  INV_X1    g0610(.A(G355), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n810), .A2(new_n811), .B1(G116), .B2(new_n219), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n806), .B1(new_n809), .B2(new_n812), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n752), .A2(new_n756), .A3(new_n805), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n748), .A2(new_n652), .ZN(new_n815));
  OAI21_X1  g0615(.A(G330), .B1(new_n746), .B2(new_n747), .ZN(new_n816));
  INV_X1    g0616(.A(new_n756), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(G396));
  NAND2_X1  g0620(.A1(new_n313), .A2(new_n661), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AND4_X1   g0622(.A1(new_n331), .A2(new_n329), .A3(new_n333), .A4(new_n822), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n328), .A2(KEYINPUT72), .B1(new_n332), .B2(new_n320), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n824), .A2(new_n331), .B1(new_n324), .B2(new_n326), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n823), .B1(new_n825), .B2(new_n821), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n697), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n823), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n335), .B2(new_n822), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n678), .B(new_n829), .C1(new_n642), .C2(new_n629), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n756), .B1(new_n831), .B2(new_n740), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n740), .B2(new_n831), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n804), .A2(new_n749), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT100), .Z(new_n835));
  OAI21_X1  g0635(.A(new_n756), .B1(new_n835), .B2(G77), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n763), .A2(G87), .ZN(new_n837));
  INV_X1    g0637(.A(G311), .ZN(new_n838));
  INV_X1    g0638(.A(new_n765), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n340), .B1(new_n769), .B2(new_n204), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(new_n779), .B2(G294), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n775), .A2(G116), .B1(new_n781), .B2(G107), .ZN(new_n842));
  AOI22_X1  g0642(.A1(G283), .A2(new_n785), .B1(new_n784), .B2(G303), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n837), .A2(new_n841), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n763), .A2(G68), .ZN(new_n845));
  INV_X1    g0645(.A(G132), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n249), .B1(new_n769), .B2(new_n345), .C1(new_n846), .C2(new_n839), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(G50), .B2(new_n781), .ZN(new_n848));
  AOI22_X1  g0648(.A1(G143), .A2(new_n779), .B1(new_n775), .B2(G159), .ZN(new_n849));
  INV_X1    g0649(.A(G150), .ZN(new_n850));
  INV_X1    g0650(.A(G137), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n849), .B1(new_n789), .B2(new_n850), .C1(new_n851), .C2(new_n800), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT34), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n845), .B(new_n848), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n852), .A2(new_n853), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n844), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n836), .B1(new_n856), .B2(new_n804), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(new_n750), .B2(new_n829), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n833), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(G384));
  OR2_X1    g0660(.A1(new_n566), .A2(KEYINPUT35), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n566), .A2(KEYINPUT35), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n861), .A2(G116), .A3(new_n862), .A4(new_n224), .ZN(new_n863));
  XOR2_X1   g0663(.A(new_n863), .B(KEYINPUT36), .Z(new_n864));
  NOR3_X1   g0664(.A1(new_n227), .A2(new_n202), .A3(new_n347), .ZN(new_n865));
  OR2_X1    g0665(.A1(new_n865), .A2(KEYINPUT101), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n865), .A2(KEYINPUT101), .B1(new_n287), .B2(G68), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n267), .B(G13), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n864), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n405), .A2(new_n661), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n428), .A2(new_n432), .A3(new_n870), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n405), .B(new_n661), .C1(new_n425), .C2(new_n427), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n826), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n659), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT37), .B1(new_n387), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n387), .A2(new_n388), .ZN(new_n876));
  AND4_X1   g0676(.A1(new_n376), .A2(new_n875), .A3(new_n377), .A4(new_n876), .ZN(new_n877));
  AND3_X1   g0677(.A1(new_n376), .A2(new_n377), .A3(new_n876), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT102), .ZN(new_n879));
  INV_X1    g0679(.A(new_n362), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n344), .A2(new_n351), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n312), .B1(new_n881), .B2(new_n353), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n880), .B1(new_n882), .B2(new_n352), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n879), .B1(new_n883), .B2(new_n659), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n387), .A2(KEYINPUT102), .A3(new_n874), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n878), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n877), .B1(new_n887), .B2(KEYINPUT37), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n886), .B1(new_n647), .B2(new_n390), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT38), .ZN(new_n890));
  NOR3_X1   g0690(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT102), .B1(new_n387), .B2(new_n874), .ZN(new_n892));
  AOI211_X1 g0692(.A(new_n879), .B(new_n659), .C1(new_n360), .C2(new_n362), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n391), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n376), .A2(new_n377), .A3(new_n876), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT37), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n878), .A2(new_n875), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT38), .B1(new_n895), .B2(new_n899), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n739), .B(new_n873), .C1(new_n891), .C2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT40), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n871), .A2(new_n872), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n829), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n613), .A2(new_n678), .B1(new_n731), .B2(new_n732), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n904), .B1(new_n905), .B2(new_n738), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n387), .A2(new_n874), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n647), .B2(new_n390), .ZN(new_n908));
  AND3_X1   g0708(.A1(new_n360), .A2(new_n362), .A3(new_n373), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n384), .B1(new_n360), .B2(new_n362), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT103), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT103), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n912), .B(new_n374), .C1(new_n883), .C2(new_n384), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n911), .A2(new_n913), .A3(new_n907), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n914), .A2(KEYINPUT37), .B1(new_n878), .B2(new_n875), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n890), .B1(new_n908), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n895), .A2(KEYINPUT38), .A3(new_n899), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n902), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n901), .A2(new_n902), .B1(new_n906), .B2(new_n918), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n919), .A2(new_n434), .A3(new_n739), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n919), .B1(new_n434), .B2(new_n739), .ZN(new_n921));
  OR3_X1    g0721(.A1(new_n920), .A2(new_n921), .A3(new_n652), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT39), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n914), .A2(KEYINPUT37), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n898), .ZN(new_n925));
  INV_X1    g0725(.A(new_n907), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n391), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT38), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n923), .B1(new_n891), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n428), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n678), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n890), .B1(new_n888), .B2(new_n889), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n933), .A2(KEYINPUT39), .A3(new_n917), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n929), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n903), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n334), .A2(new_n661), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n936), .B1(new_n830), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n891), .B2(new_n900), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n390), .A2(new_n874), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  AND3_X1   g0742(.A1(new_n935), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n650), .B1(new_n714), .B2(new_n434), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n943), .B(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n922), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n267), .B2(new_n753), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n922), .A2(new_n945), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n869), .B1(new_n947), .B2(new_n948), .ZN(G367));
  INV_X1    g0749(.A(new_n807), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n238), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n806), .B1(new_n219), .B2(new_n309), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n756), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n249), .B1(new_n765), .B2(G317), .ZN(new_n954));
  INV_X1    g0754(.A(G283), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n954), .B1(new_n205), .B2(new_n769), .C1(new_n774), .C2(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(G303), .B2(new_n779), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n763), .A2(new_n524), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n780), .A2(new_n577), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n959), .A2(KEYINPUT46), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(G311), .B2(new_n784), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n785), .A2(G294), .B1(new_n959), .B2(KEYINPUT46), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n957), .A2(new_n958), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n763), .A2(G77), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n249), .B1(new_n769), .B2(new_n346), .C1(new_n851), .C2(new_n839), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n965), .B1(G58), .B2(new_n781), .ZN(new_n966));
  AOI22_X1  g0766(.A1(G50), .A2(new_n775), .B1(new_n779), .B2(G150), .ZN(new_n967));
  AOI22_X1  g0767(.A1(G143), .A2(new_n784), .B1(new_n785), .B2(G159), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n964), .A2(new_n966), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n963), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT47), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n953), .B1(new_n971), .B2(new_n804), .ZN(new_n972));
  INV_X1    g0772(.A(new_n751), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n621), .B1(new_n618), .B2(new_n678), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n693), .A2(new_n633), .A3(new_n661), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n972), .B1(new_n973), .B2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT45), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n674), .A2(new_n679), .B1(new_n520), .B2(new_n661), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n637), .A2(new_n661), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n533), .A2(new_n661), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n557), .A2(new_n571), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n978), .B1(new_n979), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n682), .A2(KEYINPUT45), .A3(new_n983), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n979), .A2(KEYINPUT44), .A3(new_n984), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT44), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n682), .B2(new_n983), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n987), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT107), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n993), .B1(new_n677), .B2(new_n994), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n671), .A2(new_n992), .A3(KEYINPUT107), .A4(new_n676), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n676), .B(new_n680), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n816), .B(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n742), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n685), .B(KEYINPUT41), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n755), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n677), .A2(new_n984), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(KEYINPUT106), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n976), .ZN(new_n1005));
  XOR2_X1   g0805(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n676), .A2(new_n680), .A3(new_n983), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT42), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n557), .B1(new_n982), .B2(new_n520), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT105), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1013), .A2(new_n678), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1007), .B1(new_n1010), .B2(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n1010), .A2(new_n1015), .B1(KEYINPUT43), .B2(new_n976), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1016), .B1(new_n1018), .B2(new_n1007), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1003), .A2(KEYINPUT106), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1004), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1007), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1017), .A2(new_n1022), .ZN(new_n1023));
  OAI211_X1 g0823(.A(KEYINPUT106), .B(new_n1003), .C1(new_n1023), .C2(new_n1016), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n977), .B1(new_n1002), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT108), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n1028), .A2(new_n1029), .ZN(G387));
  NAND2_X1  g0830(.A1(new_n743), .A2(new_n999), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n671), .B(new_n998), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n742), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1031), .A2(new_n1033), .A3(new_n685), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n804), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n249), .B1(new_n765), .B2(G326), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n762), .B2(new_n577), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT112), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G303), .A2(new_n775), .B1(new_n779), .B2(G317), .ZN(new_n1039));
  INV_X1    g0839(.A(G322), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1039), .B1(new_n789), .B2(new_n838), .C1(new_n1040), .C2(new_n800), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT48), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n769), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n781), .A2(G294), .B1(G283), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1043), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT49), .Z(new_n1048));
  AOI21_X1  g0848(.A(new_n1038), .B1(new_n1048), .B2(KEYINPUT111), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(KEYINPUT111), .B2(new_n1048), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n762), .A2(new_n204), .ZN(new_n1051));
  INV_X1    g0851(.A(G159), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n1052), .A2(new_n800), .B1(new_n789), .B2(new_n280), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1045), .A2(new_n310), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(KEYINPUT110), .B(G150), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n340), .B1(new_n765), .B2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1054), .B(new_n1056), .C1(new_n778), .C2(new_n287), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n774), .A2(new_n346), .B1(new_n780), .B2(new_n202), .ZN(new_n1058));
  OR4_X1    g0858(.A1(new_n1051), .A2(new_n1053), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1035), .B1(new_n1050), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n806), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n810), .A2(new_n686), .B1(G107), .B2(new_n219), .ZN(new_n1062));
  AOI211_X1 g0862(.A(G45), .B(new_n687), .C1(G68), .C2(G77), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n280), .A2(G50), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT50), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n950), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1066), .A2(KEYINPUT109), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1066), .A2(KEYINPUT109), .B1(G45), .B2(new_n234), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1062), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n756), .B1(new_n1061), .B2(new_n1069), .C1(new_n676), .C2(new_n973), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1034), .B1(new_n754), .B2(new_n999), .C1(new_n1060), .C2(new_n1070), .ZN(G393));
  NAND2_X1  g0871(.A1(new_n677), .A2(new_n993), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n671), .A2(new_n992), .A3(new_n676), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1072), .A2(new_n755), .A3(new_n1073), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n800), .A2(new_n850), .B1(new_n778), .B2(new_n1052), .ZN(new_n1075));
  XOR2_X1   g0875(.A(new_n1075), .B(KEYINPUT51), .Z(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(G77), .B2(new_n1045), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n340), .B1(new_n765), .B2(G143), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n837), .B(new_n1078), .C1(new_n346), .C2(new_n780), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n1079), .A2(KEYINPUT114), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n280), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n785), .A2(G50), .B1(new_n775), .B2(new_n1081), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT115), .Z(new_n1083));
  NAND2_X1  g0883(.A1(new_n1079), .A2(KEYINPUT114), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1077), .A2(new_n1080), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n784), .A2(G317), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n838), .B2(new_n778), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT116), .Z(new_n1088));
  NOR2_X1   g0888(.A1(new_n1088), .A2(KEYINPUT52), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(KEYINPUT52), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n775), .A2(G294), .B1(G116), .B2(new_n1045), .ZN(new_n1091));
  INV_X1    g0891(.A(G303), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1091), .B1(new_n1092), .B2(new_n789), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n1093), .B(KEYINPUT117), .Z(new_n1094));
  OAI21_X1  g0894(.A(new_n340), .B1(new_n839), .B2(new_n1040), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1095), .B(new_n793), .C1(G283), .C2(new_n781), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1090), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1085), .B1(new_n1089), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n804), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n983), .A2(new_n973), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT113), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n807), .A2(new_n246), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1061), .B1(new_n684), .B2(new_n524), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n817), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1099), .A2(new_n1101), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1074), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1033), .A2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n742), .A2(new_n1032), .A3(new_n995), .A4(new_n996), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1108), .A2(new_n685), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT118), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1108), .A2(new_n1109), .A3(KEYINPUT118), .A4(new_n685), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1106), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(G390));
  INV_X1    g0915(.A(new_n685), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n739), .A2(G330), .A3(new_n829), .A4(new_n903), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n830), .A2(new_n938), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n903), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n1120), .A2(new_n931), .B1(new_n929), .B2(new_n934), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n916), .A2(new_n917), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n937), .B1(new_n711), .B2(new_n829), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n931), .B(new_n1122), .C1(new_n1123), .C2(new_n936), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1118), .B1(new_n1121), .B2(new_n1125), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n933), .A2(KEYINPUT39), .A3(new_n917), .ZN(new_n1127));
  AOI21_X1  g0927(.A(KEYINPUT39), .B1(new_n916), .B2(new_n917), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n1127), .A2(new_n1128), .B1(new_n939), .B2(new_n932), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1129), .A2(new_n1117), .A3(new_n1124), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1126), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n936), .B1(new_n740), .B2(new_n826), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n1117), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n1119), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1132), .A2(new_n1117), .A3(new_n1123), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n434), .A2(new_n741), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1136), .A2(new_n944), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1116), .B1(new_n1131), .B2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n1131), .B2(new_n1138), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n756), .B1(new_n835), .B2(new_n1081), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1142), .A2(new_n750), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n340), .B1(new_n769), .B2(new_n202), .C1(new_n767), .C2(new_n839), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(G87), .B2(new_n781), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(G116), .A2(new_n779), .B1(new_n775), .B2(new_n524), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(G107), .A2(new_n785), .B1(new_n784), .B2(G283), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n845), .A2(new_n1145), .A3(new_n1146), .A4(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT54), .B(G143), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n785), .A2(G137), .B1(new_n775), .B2(new_n1150), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1151), .B(KEYINPUT119), .Z(new_n1152));
  NAND2_X1  g0952(.A1(new_n763), .A2(G50), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n781), .A2(new_n1055), .ZN(new_n1154));
  OR2_X1    g0954(.A1(new_n1154), .A2(KEYINPUT53), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n340), .B1(new_n765), .B2(G125), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n1052), .B2(new_n769), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n779), .B2(G132), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(KEYINPUT53), .A2(new_n1154), .B1(new_n784), .B2(G128), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1153), .A2(new_n1155), .A3(new_n1158), .A4(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1148), .B1(new_n1152), .B2(new_n1160), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n1141), .B(new_n1143), .C1(new_n804), .C2(new_n1161), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n1129), .A2(new_n1117), .A3(new_n1124), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1117), .B1(new_n1129), .B2(new_n1124), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1162), .B1(new_n1165), .B2(new_n755), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1140), .A2(new_n1166), .ZN(G378));
  NAND3_X1  g0967(.A1(new_n935), .A2(new_n940), .A3(new_n942), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1122), .A2(new_n906), .A3(KEYINPUT40), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n739), .A2(new_n873), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(new_n917), .B2(new_n933), .ZN(new_n1171));
  OAI211_X1 g0971(.A(G330), .B(new_n1169), .C1(new_n1171), .C2(KEYINPUT40), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n294), .A2(new_n659), .ZN(new_n1173));
  OR2_X1    g0973(.A1(new_n303), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n303), .A2(new_n1173), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1174), .A2(new_n1175), .A3(new_n1177), .ZN(new_n1180));
  AND2_X1   g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1172), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n919), .B2(G330), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1168), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1172), .A2(new_n1181), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n901), .A2(new_n902), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1183), .A2(new_n1187), .A3(G330), .A4(new_n1169), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1186), .A2(new_n943), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1185), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1181), .A2(new_n749), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n756), .B1(new_n835), .B2(G50), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n249), .A2(G41), .ZN(new_n1193));
  AOI211_X1 g0993(.A(G50), .B(new_n1193), .C1(new_n276), .C2(new_n262), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n763), .A2(G58), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1193), .B1(new_n769), .B2(new_n346), .C1(new_n955), .C2(new_n839), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(G77), .B2(new_n781), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(G107), .A2(new_n779), .B1(new_n775), .B2(new_n310), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(G97), .A2(new_n785), .B1(new_n784), .B2(G116), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1195), .A2(new_n1197), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT58), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1194), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(G125), .A2(new_n784), .B1(new_n785), .B2(G132), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n781), .A2(new_n1150), .B1(G150), .B2(new_n1045), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(G128), .A2(new_n779), .B1(new_n775), .B2(G137), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1207));
  AOI211_X1 g1007(.A(G33), .B(G41), .C1(new_n765), .C2(G124), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1207), .B(new_n1208), .C1(new_n1052), .C2(new_n762), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1202), .B1(new_n1201), .B2(new_n1200), .C1(new_n1209), .C2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1192), .B1(new_n1211), .B2(new_n804), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1190), .A2(new_n755), .B1(new_n1191), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT57), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n1186), .A2(new_n943), .A3(new_n1188), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n941), .B1(new_n1142), .B2(new_n932), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n1186), .A2(new_n1188), .B1(new_n1216), .B2(new_n940), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n944), .A2(new_n1137), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n1165), .B2(new_n1136), .ZN(new_n1220));
  OAI211_X1 g1020(.A(KEYINPUT121), .B(new_n1214), .C1(new_n1218), .C2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(KEYINPUT57), .B1(new_n1215), .B2(new_n1217), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT120), .ZN(new_n1223));
  NOR3_X1   g1023(.A1(new_n1222), .A2(new_n1220), .A3(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1214), .B1(new_n1185), .B2(new_n1189), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n944), .A2(new_n1137), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1136), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1226), .B1(new_n1131), .B2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(KEYINPUT120), .B1(new_n1225), .B2(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1221), .B1(new_n1224), .B2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(KEYINPUT57), .B1(new_n1228), .B2(new_n1190), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n685), .B1(new_n1231), .B2(KEYINPUT121), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1213), .B1(new_n1230), .B2(new_n1232), .ZN(G375));
  NAND2_X1  g1033(.A1(new_n1219), .A2(new_n1227), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1234), .A2(new_n1001), .A3(new_n1138), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1235), .B(KEYINPUT122), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1195), .A2(new_n249), .ZN(new_n1237));
  XOR2_X1   g1037(.A(new_n1237), .B(KEYINPUT124), .Z(new_n1238));
  AOI22_X1  g1038(.A1(new_n1045), .A2(G50), .B1(G128), .B2(new_n765), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n850), .B2(new_n774), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n778), .A2(new_n851), .B1(new_n780), .B2(new_n1052), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n846), .A2(new_n800), .B1(new_n789), .B2(new_n1149), .ZN(new_n1242));
  NOR4_X1   g1042(.A1(new_n1238), .A2(new_n1240), .A3(new_n1241), .A4(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n964), .A2(new_n340), .ZN(new_n1244));
  XOR2_X1   g1044(.A(new_n1244), .B(KEYINPUT123), .Z(new_n1245));
  OAI221_X1 g1045(.A(new_n1054), .B1(new_n1092), .B2(new_n839), .C1(new_n774), .C2(new_n205), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n778), .A2(new_n955), .B1(new_n780), .B2(new_n204), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n577), .A2(new_n789), .B1(new_n800), .B2(new_n767), .ZN(new_n1248));
  NOR4_X1   g1048(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n804), .B1(new_n1243), .B2(new_n1249), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1250), .B(new_n756), .C1(G68), .C2(new_n835), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n749), .B2(new_n936), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n1136), .B2(new_n755), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1236), .A2(new_n1253), .ZN(G381));
  NOR3_X1   g1054(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1255));
  INV_X1    g1055(.A(G378), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1255), .A2(new_n1114), .A3(new_n1256), .ZN(new_n1257));
  OR4_X1    g1057(.A1(G387), .A2(G375), .A3(new_n1257), .A4(G381), .ZN(G407));
  INV_X1    g1058(.A(new_n1213), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1223), .B1(new_n1222), .B2(new_n1220), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1225), .A2(KEYINPUT120), .A3(new_n1228), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n1260), .A2(new_n1261), .B1(new_n1231), .B2(KEYINPUT121), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1214), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT121), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1116), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1259), .B1(new_n1262), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(G213), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1267), .A2(G343), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1266), .A2(new_n1256), .A3(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(G407), .A2(G213), .A3(new_n1269), .ZN(G409));
  XNOR2_X1  g1070(.A(G393), .B(new_n819), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT125), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1106), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1272), .A2(new_n1026), .A3(new_n1273), .A4(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1275), .B1(new_n1026), .B2(new_n1114), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1273), .B1(new_n1114), .B2(new_n1026), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1271), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1028), .A2(new_n1029), .A3(new_n1114), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(G393), .B(G396), .ZN(new_n1280));
  OR2_X1    g1080(.A1(new_n1114), .A2(new_n1026), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1279), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1278), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  OAI211_X1 g1084(.A(G378), .B(new_n1213), .C1(new_n1230), .C2(new_n1232), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1228), .A2(new_n1190), .A3(new_n1001), .ZN(new_n1286));
  AOI21_X1  g1086(.A(G378), .B1(new_n1286), .B2(new_n1213), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1285), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1268), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT60), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1234), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n685), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1291), .B1(new_n1234), .B2(new_n1138), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1253), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n859), .ZN(new_n1296));
  OAI211_X1 g1096(.A(G384), .B(new_n1253), .C1(new_n1293), .C2(new_n1294), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1289), .A2(new_n1290), .A3(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(KEYINPUT62), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1268), .B1(new_n1285), .B2(new_n1288), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT62), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1302), .A2(new_n1303), .A3(new_n1299), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1301), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1268), .A2(G2897), .ZN(new_n1306));
  AND3_X1   g1106(.A1(new_n1296), .A2(new_n1297), .A3(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1306), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1287), .B1(new_n1266), .B2(G378), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1309), .B1(new_n1310), .B2(new_n1268), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT61), .ZN(new_n1312));
  AOI21_X1  g1112(.A(KEYINPUT126), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1284), .B1(new_n1305), .B2(new_n1313), .ZN(new_n1314));
  AND4_X1   g1114(.A1(KEYINPUT63), .A2(new_n1289), .A3(new_n1290), .A4(new_n1299), .ZN(new_n1315));
  AOI21_X1  g1115(.A(KEYINPUT63), .B1(new_n1302), .B2(new_n1299), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1283), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT126), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1278), .A2(new_n1318), .A3(new_n1282), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1309), .ZN(new_n1320));
  OAI211_X1 g1120(.A(new_n1319), .B(new_n1312), .C1(new_n1320), .C2(new_n1302), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1317), .A2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1314), .A2(new_n1323), .ZN(G405));
  NAND2_X1  g1124(.A1(G375), .A2(new_n1256), .ZN(new_n1325));
  AND3_X1   g1125(.A1(new_n1325), .A2(new_n1285), .A3(new_n1298), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1298), .B1(new_n1325), .B2(new_n1285), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT127), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1328), .A2(new_n1329), .A3(new_n1283), .ZN(new_n1330));
  XNOR2_X1  g1130(.A(new_n1283), .B(new_n1329), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1330), .B1(new_n1328), .B2(new_n1331), .ZN(G402));
endmodule


