//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1246, new_n1247, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  INV_X1    g0009(.A(G77), .ZN(new_n210));
  INV_X1    g0010(.A(G244), .ZN(new_n211));
  INV_X1    g0011(.A(G97), .ZN(new_n212));
  INV_X1    g0012(.A(G257), .ZN(new_n213));
  OAI22_X1  g0013(.A1(new_n210), .A2(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT64), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n214), .B(new_n216), .C1(G50), .C2(G226), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G116), .A2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n217), .B(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n206), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(new_n201), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n209), .B(new_n226), .C1(new_n229), .C2(new_n232), .ZN(G361));
  XOR2_X1   g0033(.A(KEYINPUT65), .B(KEYINPUT66), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  INV_X1    g0039(.A(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(KEYINPUT2), .B(G226), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n238), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  NAND2_X1  g0051(.A1(new_n228), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G116), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n228), .A2(G107), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n255), .B(KEYINPUT23), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT22), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT3), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  AOI21_X1  g0061(.A(G20), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n257), .B1(new_n262), .B2(G87), .ZN(new_n263));
  AND2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n228), .B(G87), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(KEYINPUT22), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n254), .B(new_n256), .C1(new_n263), .C2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT24), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n266), .B(KEYINPUT22), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n271), .A2(KEYINPUT24), .A3(new_n254), .A4(new_n256), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n227), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n270), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G1), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(G13), .A3(G20), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT67), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT67), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n279), .A2(new_n276), .A3(G13), .A4(G20), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n274), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n276), .A2(G33), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n281), .A2(G107), .A3(new_n282), .A4(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G107), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n278), .A2(new_n285), .A3(new_n280), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT25), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT25), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n278), .A2(new_n288), .A3(new_n285), .A4(new_n280), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n284), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(KEYINPUT84), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT84), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n284), .A2(new_n287), .A3(new_n292), .A4(new_n289), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n275), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n213), .A2(G1698), .ZN(new_n296));
  OAI221_X1 g0096(.A(new_n296), .B1(G250), .B2(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n297));
  NAND2_X1  g0097(.A1(G33), .A2(G294), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n300));
  INV_X1    g0100(.A(G45), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n301), .A2(G1), .ZN(new_n302));
  XNOR2_X1  g0102(.A(KEYINPUT5), .B(G41), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n300), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n299), .A2(new_n300), .B1(new_n304), .B2(G264), .ZN(new_n305));
  INV_X1    g0105(.A(G41), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT5), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT5), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G41), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n302), .A2(new_n307), .A3(new_n309), .A4(G274), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT79), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT79), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n303), .A2(new_n312), .A3(G274), .A4(new_n302), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n305), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G169), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n305), .A2(G179), .A3(new_n314), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n295), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n315), .A2(G200), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n305), .A2(G190), .A3(new_n314), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n275), .A2(new_n294), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT75), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n260), .A2(new_n261), .B1(new_n240), .B2(G1698), .ZN(new_n326));
  INV_X1    g0126(.A(G226), .ZN(new_n327));
  INV_X1    g0127(.A(G1698), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n326), .A2(new_n329), .B1(G33), .B2(G97), .ZN(new_n330));
  NAND2_X1  g0130(.A1(G33), .A2(G41), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(G1), .A3(G13), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n325), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  OAI221_X1 g0133(.A(new_n329), .B1(G232), .B2(new_n328), .C1(new_n264), .C2(new_n265), .ZN(new_n334));
  NAND2_X1  g0134(.A1(G33), .A2(G97), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(KEYINPUT75), .A3(new_n300), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n276), .B1(G41), .B2(G45), .ZN(new_n338));
  INV_X1    g0138(.A(G274), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n332), .A2(new_n338), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n340), .B1(new_n341), .B2(G238), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n333), .A2(new_n337), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(KEYINPUT13), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT13), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n333), .A2(new_n337), .A3(new_n345), .A4(new_n342), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT76), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT14), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n347), .A2(G179), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n348), .A2(new_n349), .ZN(new_n351));
  INV_X1    g0151(.A(G169), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n351), .B1(new_n347), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n344), .A2(new_n346), .ZN(new_n354));
  INV_X1    g0154(.A(new_n351), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(G169), .A3(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n350), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n278), .A2(new_n280), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n222), .ZN(new_n359));
  XNOR2_X1  g0159(.A(new_n359), .B(KEYINPUT12), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n274), .B1(new_n278), .B2(new_n280), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n276), .A2(G20), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(G68), .ZN(new_n364));
  NOR2_X1   g0164(.A1(G20), .A2(G33), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n366), .A2(new_n202), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n252), .A2(new_n210), .B1(new_n228), .B2(G68), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n274), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  XNOR2_X1  g0169(.A(new_n369), .B(KEYINPUT11), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n360), .A2(new_n364), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n357), .A2(new_n371), .ZN(new_n372));
  XNOR2_X1  g0172(.A(KEYINPUT3), .B(G33), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n373), .A2(G232), .A3(new_n328), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(G238), .A3(G1698), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n374), .B(new_n375), .C1(new_n285), .C2(new_n373), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n340), .B1(new_n376), .B2(new_n300), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n341), .A2(G244), .ZN(new_n378));
  AND2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G179), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n377), .A2(new_n378), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n352), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT70), .ZN(new_n384));
  XOR2_X1   g0184(.A(KEYINPUT8), .B(G58), .Z(new_n385));
  AOI22_X1  g0185(.A1(new_n385), .A2(new_n365), .B1(G20), .B2(G77), .ZN(new_n386));
  NOR2_X1   g0186(.A1(KEYINPUT15), .A2(G87), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(KEYINPUT15), .A2(G87), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(KEYINPUT69), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT69), .ZN(new_n391));
  INV_X1    g0191(.A(new_n389), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n391), .B1(new_n392), .B2(new_n387), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n386), .B1(new_n252), .B2(new_n394), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n274), .A2(new_n395), .B1(new_n363), .B2(G77), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n358), .A2(new_n210), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n384), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n395), .A2(new_n274), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n363), .A2(G77), .ZN(new_n400));
  AND4_X1   g0200(.A1(new_n384), .A2(new_n399), .A3(new_n397), .A4(new_n400), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n381), .B(new_n383), .C1(new_n398), .C2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n372), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(G222), .A2(G1698), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n328), .A2(G223), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n373), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n406), .B(new_n300), .C1(G77), .C2(new_n373), .ZN(new_n407));
  INV_X1    g0207(.A(new_n340), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n341), .A2(G226), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(G190), .ZN(new_n411));
  OR2_X1    g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g0212(.A(KEYINPUT72), .B(G200), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n203), .A2(G20), .ZN(new_n416));
  INV_X1    g0216(.A(G150), .ZN(new_n417));
  XNOR2_X1  g0217(.A(KEYINPUT8), .B(G58), .ZN(new_n418));
  OAI221_X1 g0218(.A(new_n416), .B1(new_n417), .B2(new_n366), .C1(new_n252), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n274), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n358), .A2(new_n202), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT68), .ZN(new_n422));
  INV_X1    g0222(.A(new_n362), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n422), .B1(new_n423), .B2(new_n202), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n362), .A2(KEYINPUT68), .A3(G50), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n361), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n420), .A2(KEYINPUT9), .A3(new_n421), .A4(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n420), .A2(new_n421), .A3(new_n426), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT9), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT73), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n428), .A2(KEYINPUT73), .A3(new_n429), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n415), .A2(new_n427), .A3(new_n432), .A4(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n412), .A2(KEYINPUT74), .A3(new_n414), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT10), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g0237(.A(new_n434), .B(new_n437), .ZN(new_n438));
  OR2_X1    g0238(.A1(new_n410), .A2(G179), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n410), .A2(new_n352), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n439), .A2(new_n428), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT17), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n264), .A2(new_n265), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT7), .B1(new_n444), .B2(new_n228), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n260), .A2(KEYINPUT7), .A3(new_n228), .A4(new_n261), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(G68), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(G58), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(new_n222), .ZN(new_n450));
  OAI21_X1  g0250(.A(G20), .B1(new_n450), .B2(new_n201), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n365), .A2(G159), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n448), .A2(KEYINPUT16), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT77), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT16), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n260), .A2(new_n228), .A3(new_n261), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT7), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n222), .B1(new_n460), .B2(new_n446), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n457), .B1(new_n461), .B2(new_n453), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT77), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n448), .A2(new_n463), .A3(KEYINPUT16), .A4(new_n454), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n456), .A2(new_n274), .A3(new_n462), .A4(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n281), .A2(new_n385), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n466), .B1(new_n363), .B2(new_n385), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  AND3_X1   g0268(.A1(new_n332), .A2(G232), .A3(new_n338), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  OR2_X1    g0270(.A1(G223), .A2(G1698), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n327), .A2(G1698), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n471), .B(new_n472), .C1(new_n264), .C2(new_n265), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G87), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n408), .B(new_n470), .C1(new_n475), .C2(new_n332), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(G190), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT78), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n332), .B1(new_n473), .B2(new_n474), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(new_n340), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n478), .B1(new_n480), .B2(new_n470), .ZN(new_n481));
  NOR4_X1   g0281(.A1(new_n479), .A2(KEYINPUT78), .A3(new_n469), .A4(new_n340), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G200), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n477), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n443), .B1(new_n468), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n476), .A2(KEYINPUT78), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n480), .A2(new_n478), .A3(new_n470), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n487), .A2(new_n484), .A3(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n489), .B1(G190), .B2(new_n476), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n490), .A2(KEYINPUT17), .A3(new_n465), .A4(new_n467), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n476), .A2(G179), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n493), .B1(new_n483), .B2(new_n352), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT18), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n468), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n495), .B1(new_n468), .B2(new_n494), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT71), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(new_n398), .B2(new_n401), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n399), .A2(new_n400), .A3(new_n397), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT70), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n396), .A2(new_n384), .A3(new_n397), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT71), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n382), .A2(new_n413), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n379), .A2(G190), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n347), .A2(G190), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n371), .B1(new_n354), .B2(G200), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n492), .A2(new_n498), .A3(new_n508), .A4(new_n511), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n403), .A2(new_n442), .A3(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n413), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n223), .A2(new_n328), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n211), .A2(G1698), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n515), .B(new_n516), .C1(new_n264), .C2(new_n265), .ZN(new_n517));
  INV_X1    g0317(.A(G116), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n259), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n220), .B1(new_n302), .B2(KEYINPUT80), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT80), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n301), .B2(G1), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n332), .A2(new_n524), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n521), .A2(new_n300), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n302), .A2(G274), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n514), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n332), .B1(new_n517), .B2(new_n520), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n276), .A2(KEYINPUT80), .A3(G45), .ZN(new_n530));
  AND4_X1   g0330(.A1(G250), .A2(new_n332), .A3(new_n524), .A4(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n527), .ZN(new_n532));
  NOR4_X1   g0332(.A1(new_n529), .A2(new_n531), .A3(new_n411), .A4(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT19), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n228), .B1(new_n335), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(G97), .A2(G107), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n219), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n228), .B(G68), .C1(new_n264), .C2(new_n265), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n535), .B1(new_n252), .B2(new_n212), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n274), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n358), .A2(new_n394), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n281), .A2(G87), .A3(new_n282), .A4(new_n283), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT81), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT81), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n361), .A2(new_n548), .A3(G87), .A4(new_n283), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n545), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n542), .A2(new_n274), .B1(new_n358), .B2(new_n394), .ZN(new_n551));
  INV_X1    g0351(.A(new_n394), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n552), .A2(new_n361), .A3(new_n283), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n522), .A2(new_n332), .A3(new_n524), .ZN(new_n554));
  NOR2_X1   g0354(.A1(G238), .A2(G1698), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n555), .B1(new_n211), .B2(G1698), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n519), .B1(new_n556), .B2(new_n373), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n554), .B(new_n527), .C1(new_n557), .C2(new_n332), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n551), .A2(new_n553), .B1(new_n558), .B2(new_n352), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n526), .A2(new_n380), .A3(new_n527), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n534), .A2(new_n550), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(G244), .B(new_n328), .C1(new_n264), .C2(new_n265), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT4), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n373), .A2(KEYINPUT4), .A3(G244), .A4(new_n328), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n373), .A2(G250), .A3(G1698), .ZN(new_n567));
  NAND2_X1  g0367(.A1(G33), .A2(G283), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n300), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g0370(.A1(G257), .A2(new_n304), .B1(new_n311), .B2(new_n313), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(G200), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n281), .A2(G97), .ZN(new_n574));
  OAI21_X1  g0374(.A(G107), .B1(new_n445), .B2(new_n447), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n366), .A2(new_n210), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT6), .ZN(new_n578));
  AND2_X1   g0378(.A1(G97), .A2(G107), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n578), .B1(new_n579), .B2(new_n537), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n285), .A2(KEYINPUT6), .A3(G97), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n228), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n575), .A2(new_n577), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n574), .B1(new_n584), .B2(new_n274), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n361), .A2(G97), .A3(new_n283), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n570), .A2(G190), .A3(new_n571), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n573), .A2(new_n585), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n574), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n285), .B1(new_n460), .B2(new_n446), .ZN(new_n590));
  NOR3_X1   g0390(.A1(new_n590), .A2(new_n576), .A3(new_n582), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n589), .B(new_n586), .C1(new_n591), .C2(new_n282), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n572), .A2(new_n352), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n570), .A2(new_n380), .A3(new_n571), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n561), .A2(new_n588), .A3(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT21), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n303), .A2(new_n302), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n599), .A2(G270), .A3(new_n332), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n314), .A2(new_n600), .ZN(new_n601));
  OAI211_X1 g0401(.A(G264), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT82), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT82), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n373), .A2(new_n604), .A3(G264), .A4(G1698), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n373), .A2(G257), .A3(new_n328), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n444), .A2(G303), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n603), .A2(new_n605), .A3(new_n606), .A4(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n601), .B1(new_n300), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n273), .A2(new_n227), .B1(G20), .B2(new_n518), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n568), .B(new_n228), .C1(G33), .C2(new_n212), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n610), .A2(KEYINPUT20), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT20), .B1(new_n610), .B2(new_n611), .ZN(new_n613));
  OAI22_X1  g0413(.A1(new_n612), .A2(new_n613), .B1(G116), .B2(new_n281), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n361), .A2(G116), .A3(new_n283), .ZN(new_n615));
  OAI21_X1  g0415(.A(G169), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n598), .B1(new_n609), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n361), .A2(G116), .A3(new_n283), .ZN(new_n618));
  OAI221_X1 g0418(.A(new_n618), .B1(G116), .B2(new_n281), .C1(new_n613), .C2(new_n612), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n608), .A2(new_n300), .ZN(new_n620));
  AOI22_X1  g0420(.A1(G270), .A2(new_n304), .B1(new_n311), .B2(new_n313), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n619), .A2(new_n622), .A3(KEYINPUT21), .A4(G169), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n609), .A2(G179), .A3(new_n619), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n617), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT83), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n614), .A2(new_n615), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n626), .B(new_n627), .C1(new_n609), .C2(new_n484), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n484), .B1(new_n620), .B2(new_n621), .ZN(new_n629));
  OAI21_X1  g0429(.A(KEYINPUT83), .B1(new_n629), .B2(new_n619), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n609), .A2(G190), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n628), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n625), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  AND4_X1   g0434(.A1(new_n324), .A2(new_n513), .A3(new_n597), .A4(new_n634), .ZN(G372));
  NAND3_X1  g0435(.A1(new_n617), .A2(new_n623), .A3(new_n624), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT85), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT86), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n319), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT85), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n617), .A2(new_n623), .A3(new_n624), .A4(new_n640), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n275), .A2(new_n294), .B1(new_n316), .B2(new_n317), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(KEYINPUT86), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n637), .A2(new_n639), .A3(new_n641), .A4(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n561), .A2(new_n322), .A3(new_n588), .A4(new_n595), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n547), .A2(new_n549), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n558), .A2(new_n413), .ZN(new_n649));
  INV_X1    g0449(.A(new_n529), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n650), .A2(G190), .A3(new_n527), .A4(new_n554), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n648), .A2(new_n649), .A3(new_n651), .A4(new_n551), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n551), .A2(new_n553), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n558), .A2(new_n352), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(new_n560), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n595), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n657), .B1(new_n595), .B2(new_n656), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n659), .A2(new_n660), .B1(new_n560), .B2(new_n559), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n647), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n513), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g0463(.A(new_n663), .B(KEYINPUT87), .Z(new_n664));
  INV_X1    g0464(.A(new_n441), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n403), .A2(new_n492), .A3(new_n511), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n498), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n665), .B1(new_n667), .B2(new_n438), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n664), .A2(new_n668), .ZN(G369));
  INV_X1    g0469(.A(G13), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(G20), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  OR3_X1    g0472(.A1(new_n672), .A2(KEYINPUT27), .A3(G1), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT27), .B1(new_n672), .B2(G1), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G213), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G343), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  AOI211_X1 g0478(.A(new_n627), .B(new_n678), .C1(new_n637), .C2(new_n641), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n633), .B1(new_n619), .B2(new_n677), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G330), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n642), .A2(KEYINPUT88), .A3(new_n677), .ZN(new_n684));
  AOI21_X1  g0484(.A(KEYINPUT88), .B1(new_n642), .B2(new_n677), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n678), .B1(new_n275), .B2(new_n294), .ZN(new_n686));
  OAI22_X1  g0486(.A1(new_n684), .A2(new_n685), .B1(new_n323), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n677), .B1(new_n639), .B2(new_n643), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n625), .A2(new_n677), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n689), .B1(new_n687), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n688), .A2(new_n691), .ZN(G399));
  NOR2_X1   g0492(.A1(new_n538), .A2(G116), .ZN(new_n693));
  XOR2_X1   g0493(.A(new_n693), .B(KEYINPUT89), .Z(new_n694));
  INV_X1    g0494(.A(new_n207), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G41), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n694), .A2(G1), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n231), .B2(new_n697), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n699), .B(KEYINPUT28), .Z(new_n700));
  AOI21_X1  g0500(.A(KEYINPUT91), .B1(KEYINPUT92), .B2(KEYINPUT30), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n570), .A2(new_n571), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n299), .A2(new_n300), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n304), .A2(G264), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(KEYINPUT90), .B1(new_n705), .B2(new_n558), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n705), .A2(new_n558), .A3(KEYINPUT90), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n620), .A2(G179), .A3(new_n621), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n701), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n620), .A2(G179), .A3(new_n621), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT90), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n305), .A2(new_n713), .A3(new_n527), .A4(new_n526), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n712), .A2(new_n702), .A3(new_n706), .A4(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(KEYINPUT92), .B1(new_n715), .B2(KEYINPUT91), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT30), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n711), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(G179), .B1(new_n305), .B2(new_n314), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n719), .A2(new_n622), .A3(new_n572), .A4(new_n558), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n677), .B1(new_n718), .B2(new_n721), .ZN(new_n722));
  NOR4_X1   g0522(.A1(new_n633), .A2(new_n323), .A3(new_n596), .A4(new_n677), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT31), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n722), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI211_X1 g0525(.A(KEYINPUT31), .B(new_n677), .C1(new_n718), .C2(new_n721), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(KEYINPUT93), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT91), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n707), .A2(new_n728), .A3(new_n710), .ZN(new_n729));
  AOI21_X1  g0529(.A(KEYINPUT30), .B1(new_n729), .B2(KEYINPUT92), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n720), .B1(new_n730), .B2(new_n711), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT93), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n731), .A2(new_n732), .A3(KEYINPUT31), .A4(new_n677), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n725), .A2(new_n727), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G330), .ZN(new_n735));
  AOI211_X1 g0535(.A(KEYINPUT29), .B(new_n677), .C1(new_n647), .C2(new_n661), .ZN(new_n736));
  AND3_X1   g0536(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n737));
  AOI21_X1  g0537(.A(KEYINPUT26), .B1(new_n737), .B2(new_n561), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n655), .B1(new_n738), .B2(new_n658), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n636), .A2(new_n642), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n645), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n678), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n742), .A2(KEYINPUT29), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n736), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n735), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n700), .B1(new_n745), .B2(new_n276), .ZN(new_n746));
  XOR2_X1   g0546(.A(new_n746), .B(KEYINPUT94), .Z(G364));
  AOI21_X1  g0547(.A(new_n276), .B1(new_n671), .B2(G45), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n696), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n683), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n681), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n751), .B1(G330), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n750), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n227), .B1(G20), .B2(new_n352), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(G20), .A2(G179), .A3(G190), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G322), .ZN(new_n759));
  NAND2_X1  g0559(.A1(G20), .A2(G179), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n760), .A2(G190), .A3(G200), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G311), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G179), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G190), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G20), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G294), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n759), .B1(new_n762), .B2(new_n763), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n413), .A2(G20), .A3(new_n380), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G190), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n411), .ZN(new_n772));
  AOI22_X1  g0572(.A1(G283), .A2(new_n771), .B1(new_n772), .B2(G303), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n764), .A2(G20), .A3(new_n411), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G329), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n773), .A2(new_n444), .A3(new_n776), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n760), .A2(new_n484), .A3(G190), .ZN(new_n778));
  XNOR2_X1  g0578(.A(KEYINPUT33), .B(G317), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n769), .B(new_n777), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G326), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n757), .A2(new_n484), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n780), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n373), .B1(new_n762), .B2(new_n210), .ZN(new_n785));
  INV_X1    g0585(.A(new_n778), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n767), .A2(new_n212), .B1(new_n786), .B2(new_n222), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n785), .B(new_n787), .C1(G50), .C2(new_n782), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n772), .A2(G87), .B1(G58), .B2(new_n758), .ZN(new_n789));
  INV_X1    g0589(.A(new_n771), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n285), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G159), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n774), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g0594(.A(KEYINPUT95), .B(KEYINPUT32), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n788), .A2(new_n789), .A3(new_n792), .A4(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n756), .B1(new_n784), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(G13), .A2(G33), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(G20), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n755), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n232), .A2(new_n301), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n695), .A2(new_n373), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n803), .B(new_n804), .C1(new_n250), .C2(new_n301), .ZN(new_n805));
  INV_X1    g0605(.A(G355), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n373), .A2(new_n207), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n805), .B1(G116), .B2(new_n207), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n754), .B(new_n798), .C1(new_n802), .C2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n801), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n809), .B1(new_n752), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n753), .A2(new_n811), .ZN(G396));
  AOI21_X1  g0612(.A(new_n677), .B1(new_n647), .B2(new_n661), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT98), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n402), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n502), .A2(new_n503), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n816), .A2(KEYINPUT98), .A3(new_n383), .A4(new_n381), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n678), .B1(new_n502), .B2(new_n503), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(KEYINPUT99), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(KEYINPUT99), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n818), .A2(new_n508), .A3(new_n820), .A4(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n813), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n823), .B1(new_n402), .B2(new_n678), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n825), .B1(new_n813), .B2(new_n826), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n735), .B(new_n827), .Z(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n754), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n373), .B1(new_n772), .B2(G107), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT96), .Z(new_n831));
  AOI22_X1  g0631(.A1(new_n771), .A2(G87), .B1(G311), .B2(new_n775), .ZN(new_n832));
  AOI22_X1  g0632(.A1(G283), .A2(new_n778), .B1(new_n758), .B2(G294), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n766), .A2(G97), .B1(G303), .B2(new_n782), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n831), .A2(new_n832), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n762), .A2(new_n518), .ZN(new_n836));
  AOI22_X1  g0636(.A1(G159), .A2(new_n761), .B1(new_n758), .B2(G143), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n782), .A2(G137), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n837), .B(new_n838), .C1(new_n417), .C2(new_n786), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT34), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n766), .A2(G58), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n771), .A2(G68), .B1(G132), .B2(new_n775), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n840), .A2(new_n373), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n772), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n844), .A2(new_n202), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n835), .A2(new_n836), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n754), .B1(new_n846), .B2(new_n755), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n755), .A2(new_n799), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n847), .B1(G77), .B2(new_n849), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n850), .B(KEYINPUT97), .Z(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n800), .B2(new_n826), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n829), .A2(new_n852), .ZN(G384));
  INV_X1    g0653(.A(KEYINPUT40), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n402), .A2(new_n678), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n500), .A2(new_n504), .B1(new_n413), .B2(new_n382), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n821), .B1(new_n856), .B2(new_n507), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n815), .A2(new_n817), .B1(new_n819), .B2(KEYINPUT99), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n855), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n357), .A2(new_n371), .A3(new_n678), .ZN(new_n860));
  INV_X1    g0660(.A(new_n371), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n355), .B1(new_n354), .B2(G169), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n352), .B(new_n351), .C1(new_n344), .C2(new_n346), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n861), .B1(new_n864), .B2(new_n350), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n509), .A2(new_n510), .B1(new_n371), .B2(new_n677), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n860), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n859), .B(new_n867), .C1(new_n726), .C2(new_n725), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT102), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n461), .B2(new_n453), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n448), .A2(KEYINPUT102), .A3(new_n454), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n870), .A2(new_n871), .A3(new_n457), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n872), .A2(new_n274), .A3(new_n456), .A4(new_n464), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n467), .ZN(new_n874));
  INV_X1    g0674(.A(new_n675), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n468), .A2(new_n494), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT18), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n468), .A2(new_n494), .A3(new_n495), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n486), .A2(new_n491), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n877), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n487), .A2(new_n352), .A3(new_n488), .ZN(new_n884));
  INV_X1    g0684(.A(new_n493), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n886), .A2(new_n675), .B1(new_n873), .B2(new_n467), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n468), .A2(new_n485), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT37), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n468), .B1(new_n494), .B2(new_n875), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n490), .A2(new_n465), .A3(new_n467), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n889), .B1(KEYINPUT37), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n883), .A2(new_n893), .A3(KEYINPUT38), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n886), .A2(new_n675), .B1(new_n465), .B2(new_n467), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT37), .B1(new_n895), .B2(KEYINPUT104), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n892), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n890), .A2(new_n891), .A3(KEYINPUT104), .A4(KEYINPUT37), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT105), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n882), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n486), .A2(KEYINPUT105), .A3(new_n491), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n901), .A2(new_n498), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n468), .A2(new_n875), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n899), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n894), .B1(new_n906), .B2(KEYINPUT38), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n854), .B1(new_n868), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT38), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n876), .B1(new_n492), .B2(new_n498), .ZN(new_n910));
  NOR3_X1   g0710(.A1(new_n888), .A2(new_n895), .A3(KEYINPUT37), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT37), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n886), .A2(new_n675), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n874), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n912), .B1(new_n914), .B2(new_n891), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n909), .B1(new_n910), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT103), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n917), .A2(new_n918), .A3(new_n894), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n883), .A2(new_n893), .A3(KEYINPUT103), .A4(KEYINPUT38), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n725), .A2(new_n726), .ZN(new_n922));
  INV_X1    g0722(.A(new_n867), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n922), .A2(new_n854), .A3(new_n826), .A4(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(G330), .B1(new_n908), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n513), .A2(new_n922), .A3(G330), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n894), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n903), .A2(new_n905), .ZN(new_n930));
  INV_X1    g0730(.A(new_n899), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n929), .B1(new_n932), .B2(new_n909), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n922), .A2(new_n826), .A3(new_n923), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT40), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n868), .A2(new_n854), .A3(new_n920), .A4(new_n919), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n937), .A2(new_n513), .A3(new_n922), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n928), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT101), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n818), .A2(new_n677), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n825), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n940), .B1(new_n943), .B2(new_n923), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n941), .B1(new_n813), .B2(new_n824), .ZN(new_n945));
  NOR3_X1   g0745(.A1(new_n945), .A2(KEYINPUT101), .A3(new_n867), .ZN(new_n946));
  NOR3_X1   g0746(.A1(new_n944), .A2(new_n946), .A3(new_n921), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n919), .A2(KEYINPUT39), .A3(new_n920), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT39), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n949), .B(new_n894), .C1(new_n906), .C2(KEYINPUT38), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n860), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n498), .A2(new_n875), .ZN(new_n952));
  NOR3_X1   g0752(.A1(new_n947), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n939), .B(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n513), .B1(new_n736), .B2(new_n743), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n668), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n954), .B(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n276), .B2(new_n671), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n580), .A2(new_n581), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT100), .Z(new_n960));
  AOI21_X1  g0760(.A(new_n518), .B1(new_n960), .B2(KEYINPUT35), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n961), .B(new_n229), .C1(KEYINPUT35), .C2(new_n960), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT36), .ZN(new_n963));
  OAI21_X1  g0763(.A(G77), .B1(new_n449), .B2(new_n222), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n231), .A2(new_n964), .B1(G50), .B2(new_n222), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n965), .A2(G1), .A3(new_n670), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n958), .A2(new_n963), .A3(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT106), .Z(G367));
  AND2_X1   g0768(.A1(new_n687), .A2(new_n690), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n595), .A2(new_n678), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT107), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n592), .A2(new_n677), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n588), .A2(new_n595), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n969), .A2(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n976));
  XNOR2_X1  g0776(.A(new_n975), .B(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n974), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n595), .B1(new_n978), .B2(new_n319), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n678), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n550), .A2(new_n678), .ZN(new_n982));
  MUX2_X1   g0782(.A(new_n656), .B(new_n655), .S(new_n982), .Z(new_n983));
  INV_X1    g0783(.A(KEYINPUT43), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n983), .A2(new_n984), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n981), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n977), .A2(new_n984), .A3(new_n983), .A4(new_n980), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n688), .A2(new_n978), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n989), .B(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n691), .A2(new_n974), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT109), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT44), .ZN(new_n995));
  NOR3_X1   g0795(.A1(new_n691), .A2(new_n974), .A3(KEYINPUT109), .ZN(new_n996));
  OR3_X1    g0796(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n691), .A2(new_n974), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT45), .Z(new_n999));
  OAI21_X1  g0799(.A(new_n995), .B1(new_n994), .B2(new_n996), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n997), .A2(new_n688), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n683), .A2(new_n690), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(new_n687), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n745), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n696), .B(KEYINPUT41), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n748), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n991), .A2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(KEYINPUT112), .B(G137), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n775), .A2(new_n1009), .B1(G143), .B2(new_n782), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n771), .A2(G77), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n373), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT111), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1010), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n1012), .A2(new_n1013), .B1(G150), .B2(new_n758), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G50), .A2(new_n761), .B1(new_n778), .B2(G159), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n766), .A2(G68), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n1014), .B(new_n1018), .C1(G58), .C2(new_n772), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n790), .A2(new_n212), .ZN(new_n1020));
  INV_X1    g0820(.A(G317), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n444), .B1(new_n774), .B2(new_n1021), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n766), .A2(G107), .B1(G283), .B2(new_n761), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n758), .ZN(new_n1024));
  INV_X1    g0824(.A(G303), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1023), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NOR3_X1   g0826(.A1(new_n1020), .A2(new_n1022), .A3(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n763), .B2(new_n783), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G294), .B2(new_n778), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n772), .A2(G116), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT46), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1019), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT47), .Z(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n755), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n983), .A2(new_n801), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n804), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n802), .B1(new_n207), .B2(new_n394), .C1(new_n238), .C2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1034), .A2(new_n750), .A3(new_n1035), .A4(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT113), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1008), .A2(new_n1039), .ZN(G387));
  OR2_X1    g0840(.A1(new_n687), .A2(new_n810), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(G311), .A2(new_n778), .B1(new_n782), .B2(G322), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n1025), .B2(new_n762), .C1(new_n1021), .C2(new_n1024), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT48), .ZN(new_n1044));
  INV_X1    g0844(.A(G283), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1044), .B1(new_n1045), .B2(new_n767), .C1(new_n768), .C2(new_n844), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT49), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n771), .A2(G116), .B1(G326), .B2(new_n775), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1047), .A2(new_n444), .A3(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n844), .A2(new_n210), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n552), .A2(new_n766), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n202), .B2(new_n1024), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1050), .B(new_n1052), .C1(G150), .C2(new_n775), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n786), .A2(new_n418), .B1(new_n783), .B2(new_n793), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1020), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n761), .A2(G68), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1053), .A2(new_n373), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n756), .B1(new_n1049), .B2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n243), .A2(new_n301), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT114), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n418), .A2(G50), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT50), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(G68), .A2(G77), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n694), .A2(new_n1062), .A3(new_n301), .A4(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1060), .A2(new_n804), .A3(new_n1064), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(G107), .B2(new_n207), .C1(new_n694), .C2(new_n807), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n754), .B(new_n1058), .C1(new_n802), .C2(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1003), .A2(new_n749), .B1(new_n1041), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n745), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n1003), .A2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n696), .B1(new_n1003), .B2(new_n1069), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1068), .B1(new_n1070), .B2(new_n1071), .ZN(G393));
  NAND2_X1  g0872(.A1(new_n1070), .A2(new_n1001), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n688), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1076), .A2(KEYINPUT115), .A3(new_n1001), .ZN(new_n1077));
  OR3_X1    g0877(.A1(new_n1074), .A2(KEYINPUT115), .A3(new_n1075), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n696), .B(new_n1073), .C1(new_n1079), .C2(new_n1070), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n749), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n802), .B1(new_n212), .B2(new_n207), .C1(new_n247), .C2(new_n1036), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n750), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT116), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G150), .A2(new_n782), .B1(new_n758), .B2(G159), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT51), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(G87), .B2(new_n771), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n772), .A2(G68), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n444), .B1(G50), .B2(new_n778), .ZN(new_n1089));
  INV_X1    g0889(.A(G143), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n762), .A2(new_n418), .B1(new_n1090), .B2(new_n774), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(G77), .B2(new_n766), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .A4(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n792), .B1(new_n1045), .B2(new_n844), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(G116), .B2(new_n766), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n775), .A2(G322), .B1(new_n761), .B2(G294), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(G311), .A2(new_n758), .B1(new_n782), .B2(G317), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT52), .Z(new_n1098));
  NAND4_X1  g0898(.A1(new_n1095), .A2(new_n444), .A3(new_n1096), .A4(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n786), .A2(new_n1025), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1093), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1084), .B1(new_n1101), .B2(new_n755), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n974), .B2(new_n810), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1080), .A2(new_n1081), .A3(new_n1103), .ZN(G390));
  INV_X1    g0904(.A(KEYINPUT118), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n668), .A2(new_n955), .A3(new_n927), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n734), .A2(G330), .A3(new_n826), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n867), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n922), .A2(G330), .A3(new_n826), .A4(new_n923), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n945), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n634), .A2(new_n324), .A3(new_n597), .A4(new_n678), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1112), .A2(KEYINPUT31), .B1(new_n731), .B2(new_n677), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n726), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n826), .B(G330), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n867), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n734), .A2(G330), .A3(new_n826), .A4(new_n923), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n942), .B1(new_n742), .B2(new_n823), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT117), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n942), .B(KEYINPUT117), .C1(new_n742), .C2(new_n823), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n1116), .A2(new_n1117), .A3(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1107), .B1(new_n1111), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n860), .B1(new_n945), .B2(new_n867), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n948), .A2(new_n1125), .A3(new_n950), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1120), .A2(new_n923), .A3(new_n1121), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1127), .A2(new_n907), .A3(new_n860), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n1126), .A2(new_n1128), .A3(new_n1117), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1110), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1130));
  NOR3_X1   g0930(.A1(new_n1124), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1105), .B1(new_n1131), .B2(new_n697), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1110), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1126), .A2(new_n1128), .A3(new_n1117), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n1124), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1116), .A2(new_n1117), .A3(new_n1122), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(G330), .A2(new_n868), .B1(new_n1108), .B2(new_n867), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1139), .B1(new_n1140), .B2(new_n945), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1135), .A2(new_n1141), .A3(new_n1136), .A4(new_n1107), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1142), .A2(KEYINPUT118), .A3(new_n696), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1132), .A2(new_n1138), .A3(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1137), .A2(new_n748), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n948), .A2(new_n799), .A3(new_n950), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n772), .A2(G150), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n1147), .B(KEYINPUT53), .Z(new_n1148));
  INV_X1    g0948(.A(G128), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n767), .A2(new_n793), .B1(new_n1149), .B2(new_n783), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n444), .B(new_n1150), .C1(new_n771), .C2(G50), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(KEYINPUT54), .B(G143), .ZN(new_n1152));
  INV_X1    g0952(.A(G125), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n762), .A2(new_n1152), .B1(new_n1153), .B2(new_n774), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(new_n778), .B2(new_n1009), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1148), .A2(new_n1151), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(G132), .B2(new_n758), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n771), .A2(G68), .B1(G107), .B2(new_n778), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n1158), .B1(new_n212), .B2(new_n762), .C1(new_n1045), .C2(new_n783), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n774), .A2(new_n768), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n844), .A2(new_n219), .B1(new_n210), .B2(new_n767), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n444), .B1(new_n1024), .B2(new_n518), .ZN(new_n1162));
  NOR4_X1   g0962(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n755), .B1(new_n1157), .B2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1146), .A2(new_n750), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(new_n418), .B2(new_n848), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1145), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1144), .A2(new_n1167), .ZN(G378));
  INV_X1    g0968(.A(G124), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n259), .B1(new_n774), .B2(new_n1169), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G132), .A2(new_n778), .B1(new_n761), .B2(G137), .ZN(new_n1171));
  XOR2_X1   g0971(.A(new_n1171), .B(KEYINPUT120), .Z(new_n1172));
  OAI221_X1 g0972(.A(new_n1172), .B1(new_n1153), .B2(new_n783), .C1(new_n844), .C2(new_n1152), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G128), .B2(new_n758), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n417), .B2(new_n767), .ZN(new_n1175));
  AOI211_X1 g0975(.A(G41), .B(new_n1170), .C1(new_n1175), .C2(KEYINPUT59), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1176), .B1(KEYINPUT59), .B2(new_n1175), .C1(new_n793), .C2(new_n790), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n202), .B1(new_n264), .B2(G41), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1050), .B1(new_n552), .B2(new_n761), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n449), .B2(new_n790), .C1(new_n518), .C2(new_n783), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n373), .B1(new_n775), .B2(G283), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1181), .B(new_n1017), .C1(new_n1024), .C2(new_n285), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n786), .A2(new_n212), .ZN(new_n1183));
  NOR4_X1   g0983(.A1(new_n1180), .A2(G41), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1178), .B1(new_n1184), .B2(KEYINPUT58), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(KEYINPUT119), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1184), .A2(KEYINPUT58), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1177), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1185), .A2(KEYINPUT119), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n755), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n442), .A2(new_n428), .A3(new_n875), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n428), .A2(new_n875), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n438), .A2(new_n441), .A3(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n1191), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1194), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1190), .B(new_n750), .C1(new_n800), .C2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(new_n202), .B2(new_n848), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n947), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n952), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n951), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1198), .B1(new_n937), .B2(G330), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n682), .B(new_n1197), .C1(new_n935), .C2(new_n936), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1204), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n926), .A2(new_n1197), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n937), .A2(G330), .A3(new_n1198), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1208), .A2(new_n953), .A3(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1207), .A2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1200), .B1(new_n1211), .B2(new_n749), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1207), .A2(new_n1210), .B1(new_n1142), .B2(new_n1107), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n696), .B1(new_n1213), .B2(KEYINPUT57), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1142), .A2(new_n1107), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n1211), .A2(KEYINPUT57), .A3(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1212), .B1(new_n1214), .B2(new_n1216), .ZN(G375));
  OAI211_X1 g1017(.A(new_n1106), .B(new_n1139), .C1(new_n1140), .C2(new_n945), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1124), .A2(new_n1218), .A3(new_n1005), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1009), .A2(new_n758), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n1149), .B2(new_n774), .C1(new_n767), .C2(new_n202), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n373), .B1(new_n790), .B2(new_n449), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT121), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1222), .A2(new_n1223), .B1(G150), .B2(new_n761), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n782), .A2(G132), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1224), .B(new_n1225), .C1(new_n786), .C2(new_n1152), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1221), .B(new_n1226), .C1(G159), .C2(new_n772), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n1223), .B2(new_n1222), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n783), .A2(new_n768), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1011), .B1(new_n285), .B2(new_n762), .C1(new_n1025), .C2(new_n774), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n1229), .B(new_n1230), .C1(G97), .C2(new_n772), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n373), .B1(new_n758), .B2(G283), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n778), .A2(G116), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1231), .A2(new_n1051), .A3(new_n1232), .A4(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n756), .B1(new_n1228), .B2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n750), .B1(new_n923), .B2(new_n800), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n1235), .B(new_n1236), .C1(new_n222), .C2(new_n848), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n1141), .B2(new_n749), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1219), .A2(new_n1238), .ZN(G381));
  XOR2_X1   g1039(.A(G375), .B(KEYINPUT122), .Z(new_n1240));
  NOR2_X1   g1040(.A1(new_n1240), .A2(G378), .ZN(new_n1241));
  INV_X1    g1041(.A(G381), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(G390), .A2(G384), .A3(G387), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(G393), .A2(G396), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1241), .A2(new_n1242), .A3(new_n1243), .A4(new_n1244), .ZN(G407));
  INV_X1    g1045(.A(G213), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(new_n1241), .B2(new_n676), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(G407), .ZN(G409));
  NAND3_X1  g1048(.A1(G390), .A2(new_n1008), .A3(new_n1039), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(G387), .A2(new_n1080), .A3(new_n1081), .A4(new_n1103), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1249), .A2(KEYINPUT124), .A3(new_n1250), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(G393), .B(G396), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1251), .B(new_n1253), .C1(KEYINPUT124), .C2(new_n1249), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1249), .A2(new_n1250), .A3(new_n1252), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT125), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1249), .A2(KEYINPUT125), .A3(new_n1250), .A4(new_n1252), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1254), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1211), .A2(new_n1005), .A3(new_n1215), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1212), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1261), .A2(new_n1167), .A3(new_n1144), .ZN(new_n1262));
  INV_X1    g1062(.A(G378), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1262), .B1(G375), .B2(new_n1263), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1246), .A2(G343), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT60), .ZN(new_n1267));
  OR2_X1    g1067(.A1(new_n1218), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1218), .A2(new_n1267), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1268), .A2(new_n1269), .A3(new_n696), .A4(new_n1124), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1238), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1271), .A2(new_n829), .A3(new_n852), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1270), .A2(G384), .A3(new_n1238), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  XOR2_X1   g1075(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1276));
  NAND4_X1  g1076(.A1(new_n1264), .A2(new_n1266), .A3(new_n1275), .A4(new_n1276), .ZN(new_n1277));
  OAI211_X1 g1077(.A(G378), .B(new_n1212), .C1(new_n1216), .C2(new_n1214), .ZN(new_n1278));
  AOI211_X1 g1078(.A(new_n1265), .B(new_n1274), .C1(new_n1278), .C2(new_n1262), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1277), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT61), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1265), .A2(G2897), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1274), .B(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1265), .B1(new_n1278), .B2(new_n1262), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1282), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1259), .B1(new_n1281), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT123), .ZN(new_n1289));
  OAI21_X1  g1089(.A(KEYINPUT63), .B1(new_n1279), .B2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1254), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1274), .B(new_n1283), .ZN(new_n1293));
  AOI21_X1  g1093(.A(KEYINPUT61), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1264), .A2(new_n1266), .A3(new_n1275), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT63), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1295), .A2(KEYINPUT123), .A3(new_n1296), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1290), .A2(new_n1291), .A3(new_n1294), .A4(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1288), .A2(new_n1298), .ZN(G405));
  NAND2_X1  g1099(.A1(new_n1275), .A2(KEYINPUT127), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(G375), .A2(new_n1263), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT127), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1274), .A2(new_n1302), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1300), .A2(new_n1278), .A3(new_n1301), .A4(new_n1303), .ZN(new_n1304));
  AND2_X1   g1104(.A1(new_n1301), .A2(new_n1278), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1304), .B1(new_n1305), .B2(new_n1303), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(new_n1306), .B(new_n1291), .ZN(G402));
endmodule


