

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747;

  XOR2_X1 U374 ( .A(KEYINPUT69), .B(KEYINPUT68), .Z(n436) );
  INV_X2 U375 ( .A(G953), .ZN(n726) );
  NAND2_X1 U376 ( .A1(G234), .A2(n726), .ZN(n435) );
  XNOR2_X1 U377 ( .A(n436), .B(n435), .ZN(n438) );
  XNOR2_X1 U378 ( .A(n438), .B(n437), .ZN(n490) );
  AND2_X4 U379 ( .A1(n405), .A2(n622), .ZN(n717) );
  NAND2_X2 U380 ( .A1(n555), .A2(n590), .ZN(n613) );
  XNOR2_X2 U381 ( .A(n447), .B(n446), .ZN(n590) );
  XNOR2_X2 U382 ( .A(n472), .B(n450), .ZN(n732) );
  INV_X1 U383 ( .A(n618), .ZN(n721) );
  NAND2_X1 U384 ( .A1(n658), .A2(n654), .ZN(n532) );
  NAND2_X1 U385 ( .A1(n399), .A2(n398), .ZN(n405) );
  AND2_X1 U386 ( .A1(n395), .A2(n407), .ZN(n399) );
  OR2_X1 U387 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U388 ( .A(n619), .B(n434), .ZN(n433) );
  NAND2_X1 U389 ( .A1(n571), .A2(n570), .ZN(n619) );
  AND2_X1 U390 ( .A1(n557), .A2(n666), .ZN(n558) );
  NOR2_X1 U391 ( .A1(n401), .A2(n402), .ZN(n539) );
  XNOR2_X1 U392 ( .A(n521), .B(n354), .ZN(n389) );
  XNOR2_X2 U393 ( .A(n509), .B(n476), .ZN(n424) );
  XNOR2_X1 U394 ( .A(n510), .B(n430), .ZN(n733) );
  XNOR2_X1 U395 ( .A(n390), .B(G146), .ZN(n510) );
  XNOR2_X1 U396 ( .A(G104), .B(G101), .ZN(n452) );
  XNOR2_X1 U397 ( .A(G110), .B(G107), .ZN(n451) );
  XNOR2_X1 U398 ( .A(G128), .B(G119), .ZN(n372) );
  XNOR2_X1 U399 ( .A(G110), .B(KEYINPUT23), .ZN(n374) );
  NOR2_X1 U400 ( .A1(n365), .A2(n356), .ZN(n352) );
  NOR2_X1 U401 ( .A1(n365), .A2(n356), .ZN(n540) );
  XNOR2_X1 U402 ( .A(n588), .B(KEYINPUT6), .ZN(n607) );
  XNOR2_X2 U403 ( .A(n580), .B(n579), .ZN(n593) );
  XNOR2_X2 U404 ( .A(n424), .B(n493), .ZN(n472) );
  XNOR2_X1 U405 ( .A(n644), .B(KEYINPUT91), .ZN(n404) );
  INV_X1 U406 ( .A(G125), .ZN(n390) );
  INV_X1 U407 ( .A(KEYINPUT45), .ZN(n413) );
  NOR2_X1 U408 ( .A1(n415), .A2(n616), .ZN(n414) );
  NAND2_X1 U409 ( .A1(n682), .A2(n590), .ZN(n611) );
  AND2_X1 U410 ( .A1(n355), .A2(n363), .ZN(n362) );
  OR2_X1 U411 ( .A1(n536), .A2(n403), .ZN(n400) );
  INV_X1 U412 ( .A(KEYINPUT65), .ZN(n411) );
  INV_X1 U413 ( .A(KEYINPUT44), .ZN(n393) );
  XNOR2_X1 U414 ( .A(n532), .B(KEYINPUT105), .ZN(n697) );
  XNOR2_X1 U415 ( .A(n416), .B(KEYINPUT71), .ZN(n476) );
  INV_X1 U416 ( .A(G131), .ZN(n416) );
  XOR2_X1 U417 ( .A(G140), .B(KEYINPUT102), .Z(n483) );
  XNOR2_X1 U418 ( .A(n480), .B(G122), .ZN(n420) );
  XNOR2_X1 U419 ( .A(G143), .B(G104), .ZN(n478) );
  XOR2_X1 U420 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n479) );
  NOR2_X1 U421 ( .A1(n475), .A2(n367), .ZN(n366) );
  NOR2_X1 U422 ( .A1(n382), .A2(KEYINPUT83), .ZN(n367) );
  INV_X1 U423 ( .A(KEYINPUT112), .ZN(n383) );
  XNOR2_X1 U424 ( .A(n586), .B(n585), .ZN(n600) );
  XNOR2_X1 U425 ( .A(n584), .B(KEYINPUT77), .ZN(n585) );
  XNOR2_X1 U426 ( .A(n426), .B(n425), .ZN(n442) );
  XNOR2_X1 U427 ( .A(n441), .B(KEYINPUT99), .ZN(n425) );
  NOR2_X1 U428 ( .A1(G953), .A2(G237), .ZN(n481) );
  XNOR2_X1 U429 ( .A(n372), .B(n376), .ZN(n371) );
  XOR2_X1 U430 ( .A(KEYINPUT92), .B(KEYINPUT8), .Z(n437) );
  XNOR2_X1 U431 ( .A(KEYINPUT70), .B(KEYINPUT10), .ZN(n430) );
  NAND2_X1 U432 ( .A1(n410), .A2(n408), .ZN(n407) );
  NAND2_X1 U433 ( .A1(n431), .A2(n409), .ZN(n408) );
  NAND2_X1 U434 ( .A1(n397), .A2(n358), .ZN(n398) );
  NOR2_X1 U435 ( .A1(n611), .A2(n607), .ZN(n592) );
  NAND2_X1 U436 ( .A1(G234), .A2(G237), .ZN(n460) );
  XNOR2_X1 U437 ( .A(n489), .B(n488), .ZN(n544) );
  NAND2_X1 U438 ( .A1(n717), .A2(G472), .ZN(n422) );
  INV_X1 U439 ( .A(KEYINPUT46), .ZN(n384) );
  INV_X1 U440 ( .A(n747), .ZN(n415) );
  XOR2_X1 U441 ( .A(KEYINPUT94), .B(KEYINPUT48), .Z(n560) );
  OR2_X1 U442 ( .A1(G237), .A2(G902), .ZN(n518) );
  NAND2_X1 U443 ( .A1(KEYINPUT2), .A2(n411), .ZN(n409) );
  NAND2_X1 U444 ( .A1(n431), .A2(n411), .ZN(n406) );
  NAND2_X1 U445 ( .A1(n617), .A2(n411), .ZN(n410) );
  XNOR2_X1 U446 ( .A(n511), .B(n510), .ZN(n512) );
  XOR2_X1 U447 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n511) );
  XNOR2_X1 U448 ( .A(n567), .B(KEYINPUT38), .ZN(n693) );
  INV_X1 U449 ( .A(n525), .ZN(n382) );
  INV_X1 U450 ( .A(G902), .ZN(n499) );
  INV_X1 U451 ( .A(KEYINPUT28), .ZN(n380) );
  INV_X1 U452 ( .A(KEYINPUT66), .ZN(n446) );
  OR2_X1 U453 ( .A1(n623), .A2(G902), .ZN(n412) );
  XNOR2_X1 U454 ( .A(G101), .B(G146), .ZN(n467) );
  XOR2_X1 U455 ( .A(KEYINPUT5), .B(G137), .Z(n468) );
  XOR2_X1 U456 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n504) );
  XNOR2_X1 U457 ( .A(G122), .B(KEYINPUT16), .ZN(n503) );
  XNOR2_X1 U458 ( .A(KEYINPUT3), .B(G119), .ZN(n465) );
  XOR2_X1 U459 ( .A(G113), .B(G116), .Z(n466) );
  XOR2_X1 U460 ( .A(G116), .B(G122), .Z(n494) );
  XOR2_X1 U461 ( .A(G107), .B(KEYINPUT7), .Z(n492) );
  XNOR2_X1 U462 ( .A(n419), .B(n418), .ZN(n631) );
  XNOR2_X1 U463 ( .A(n477), .B(n484), .ZN(n418) );
  XNOR2_X1 U464 ( .A(n420), .B(n485), .ZN(n419) );
  XNOR2_X1 U465 ( .A(n378), .B(n377), .ZN(n530) );
  INV_X1 U466 ( .A(KEYINPUT114), .ZN(n377) );
  NAND2_X1 U467 ( .A1(n555), .A2(n379), .ZN(n378) );
  XNOR2_X1 U468 ( .A(n528), .B(n380), .ZN(n379) );
  XNOR2_X1 U469 ( .A(KEYINPUT95), .B(KEYINPUT0), .ZN(n579) );
  XNOR2_X1 U470 ( .A(n620), .B(n736), .ZN(n734) );
  XNOR2_X1 U471 ( .A(n375), .B(n733), .ZN(n429) );
  NAND2_X1 U472 ( .A1(n490), .A2(G221), .ZN(n428) );
  XNOR2_X1 U473 ( .A(KEYINPUT84), .B(G146), .ZN(n454) );
  INV_X1 U474 ( .A(n620), .ZN(n669) );
  XNOR2_X1 U475 ( .A(n386), .B(KEYINPUT35), .ZN(n744) );
  NAND2_X1 U476 ( .A1(n545), .A2(n417), .ZN(n658) );
  INV_X1 U477 ( .A(KEYINPUT113), .ZN(n360) );
  AND2_X1 U478 ( .A1(n382), .A2(KEYINPUT83), .ZN(n353) );
  NOR2_X1 U479 ( .A1(n520), .A2(n519), .ZN(n354) );
  XNOR2_X1 U480 ( .A(n440), .B(KEYINPUT20), .ZN(n444) );
  XNOR2_X1 U481 ( .A(n391), .B(n413), .ZN(n618) );
  OR2_X1 U482 ( .A1(n657), .A2(n538), .ZN(n355) );
  AND2_X1 U483 ( .A1(n370), .A2(n353), .ZN(n356) );
  XOR2_X1 U484 ( .A(n623), .B(KEYINPUT62), .Z(n357) );
  XNOR2_X1 U485 ( .A(n429), .B(n428), .ZN(n716) );
  AND2_X1 U486 ( .A1(n432), .A2(KEYINPUT65), .ZN(n358) );
  XNOR2_X2 U487 ( .A(n459), .B(n458), .ZN(n555) );
  XNOR2_X1 U488 ( .A(n359), .B(n560), .ZN(n571) );
  NAND2_X1 U489 ( .A1(n558), .A2(n559), .ZN(n359) );
  NAND2_X1 U490 ( .A1(n746), .A2(n745), .ZN(n385) );
  XNOR2_X2 U491 ( .A(n543), .B(KEYINPUT40), .ZN(n746) );
  INV_X1 U492 ( .A(KEYINPUT83), .ZN(n381) );
  XNOR2_X1 U493 ( .A(n732), .B(n456), .ZN(n638) );
  XNOR2_X1 U494 ( .A(n385), .B(n384), .ZN(n557) );
  NOR2_X1 U495 ( .A1(n598), .A2(n744), .ZN(n606) );
  XNOR2_X1 U496 ( .A(n394), .B(n393), .ZN(n392) );
  NAND2_X1 U497 ( .A1(n392), .A2(n414), .ZN(n391) );
  NOR2_X1 U498 ( .A1(n618), .A2(n406), .ZN(n396) );
  NOR2_X1 U499 ( .A1(n672), .A2(n594), .ZN(n388) );
  NAND2_X2 U500 ( .A1(n561), .A2(n660), .ZN(n543) );
  NOR2_X1 U501 ( .A1(n404), .A2(n400), .ZN(n402) );
  XNOR2_X2 U502 ( .A(n361), .B(n360), .ZN(n644) );
  NAND2_X1 U503 ( .A1(n352), .A2(n522), .ZN(n361) );
  NAND2_X1 U504 ( .A1(n536), .A2(n403), .ZN(n363) );
  NAND2_X1 U505 ( .A1(n364), .A2(n362), .ZN(n401) );
  NAND2_X1 U506 ( .A1(n534), .A2(n535), .ZN(n536) );
  NAND2_X1 U507 ( .A1(n404), .A2(n403), .ZN(n364) );
  NAND2_X1 U508 ( .A1(n368), .A2(n366), .ZN(n365) );
  NAND2_X1 U509 ( .A1(n369), .A2(n381), .ZN(n368) );
  INV_X1 U510 ( .A(n370), .ZN(n369) );
  XNOR2_X2 U511 ( .A(n613), .B(n383), .ZN(n370) );
  XNOR2_X1 U512 ( .A(n373), .B(n371), .ZN(n375) );
  XNOR2_X1 U513 ( .A(n449), .B(n374), .ZN(n373) );
  XNOR2_X2 U514 ( .A(G140), .B(G137), .ZN(n449) );
  INV_X1 U515 ( .A(KEYINPUT24), .ZN(n376) );
  NOR2_X1 U516 ( .A1(n524), .A2(n678), .ZN(n679) );
  NOR2_X1 U517 ( .A1(n524), .A2(n527), .ZN(n551) );
  AND2_X1 U518 ( .A1(n607), .A2(n524), .ZN(n608) );
  NOR2_X1 U519 ( .A1(n601), .A2(n524), .ZN(n602) );
  NOR2_X1 U520 ( .A1(n587), .A2(n524), .ZN(n589) );
  INV_X1 U521 ( .A(n530), .ZN(n547) );
  NAND2_X1 U522 ( .A1(n387), .A2(n597), .ZN(n386) );
  XNOR2_X1 U523 ( .A(n388), .B(n596), .ZN(n387) );
  INV_X1 U524 ( .A(n389), .ZN(n567) );
  NAND2_X1 U525 ( .A1(n389), .A2(n692), .ZN(n529) );
  AND2_X1 U526 ( .A1(n597), .A2(n389), .ZN(n522) );
  NAND2_X1 U527 ( .A1(n606), .A2(n743), .ZN(n394) );
  NAND2_X1 U528 ( .A1(n396), .A2(n433), .ZN(n395) );
  NAND2_X1 U529 ( .A1(n433), .A2(n721), .ZN(n397) );
  INV_X1 U530 ( .A(KEYINPUT89), .ZN(n403) );
  XNOR2_X1 U531 ( .A(n422), .B(n357), .ZN(n421) );
  NAND2_X1 U532 ( .A1(n421), .A2(n641), .ZN(n427) );
  INV_X1 U533 ( .A(n682), .ZN(n563) );
  XNOR2_X2 U534 ( .A(n412), .B(G472), .ZN(n588) );
  XNOR2_X2 U535 ( .A(n555), .B(KEYINPUT1), .ZN(n682) );
  XNOR2_X1 U536 ( .A(n509), .B(n512), .ZN(n516) );
  NOR2_X2 U537 ( .A1(n600), .A2(n682), .ZN(n609) );
  INV_X1 U538 ( .A(n654), .ZN(n662) );
  NAND2_X1 U539 ( .A1(n531), .A2(n544), .ZN(n654) );
  INV_X1 U540 ( .A(n544), .ZN(n417) );
  XNOR2_X2 U541 ( .A(n423), .B(n439), .ZN(n617) );
  XNOR2_X2 U542 ( .A(G902), .B(KEYINPUT97), .ZN(n423) );
  XNOR2_X2 U543 ( .A(n448), .B(KEYINPUT4), .ZN(n509) );
  NAND2_X1 U544 ( .A1(n444), .A2(G217), .ZN(n426) );
  XNOR2_X1 U545 ( .A(n427), .B(KEYINPUT63), .ZN(G57) );
  INV_X1 U546 ( .A(n617), .ZN(n431) );
  INV_X1 U547 ( .A(KEYINPUT2), .ZN(n432) );
  INV_X1 U548 ( .A(KEYINPUT82), .ZN(n434) );
  AND2_X1 U549 ( .A1(n709), .A2(G953), .ZN(n720) );
  NOR2_X1 U550 ( .A1(n716), .A2(G902), .ZN(n443) );
  INV_X1 U551 ( .A(KEYINPUT15), .ZN(n439) );
  NAND2_X1 U552 ( .A1(n617), .A2(G234), .ZN(n440) );
  XOR2_X1 U553 ( .A(KEYINPUT100), .B(KEYINPUT25), .Z(n441) );
  XNOR2_X1 U554 ( .A(n443), .B(n442), .ZN(n523) );
  NAND2_X1 U555 ( .A1(n444), .A2(G221), .ZN(n445) );
  XNOR2_X2 U556 ( .A(KEYINPUT21), .B(n445), .ZN(n677) );
  XNOR2_X1 U557 ( .A(KEYINPUT101), .B(n677), .ZN(n582) );
  NAND2_X1 U558 ( .A1(n523), .A2(n582), .ZN(n447) );
  XNOR2_X2 U559 ( .A(KEYINPUT64), .B(KEYINPUT67), .ZN(n448) );
  XNOR2_X1 U560 ( .A(G143), .B(G128), .ZN(n514) );
  XNOR2_X1 U561 ( .A(n514), .B(G134), .ZN(n493) );
  XNOR2_X1 U562 ( .A(n449), .B(KEYINPUT98), .ZN(n450) );
  XNOR2_X1 U563 ( .A(n452), .B(n451), .ZN(n502) );
  NAND2_X1 U564 ( .A1(n726), .A2(G227), .ZN(n453) );
  XNOR2_X1 U565 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U566 ( .A(n502), .B(n455), .ZN(n456) );
  OR2_X2 U567 ( .A1(n638), .A2(G902), .ZN(n459) );
  INV_X1 U568 ( .A(KEYINPUT73), .ZN(n457) );
  XNOR2_X1 U569 ( .A(n457), .B(G469), .ZN(n458) );
  XNOR2_X1 U570 ( .A(KEYINPUT14), .B(n460), .ZN(n706) );
  INV_X1 U571 ( .A(G952), .ZN(n709) );
  NOR2_X1 U572 ( .A1(G953), .A2(n709), .ZN(n574) );
  NAND2_X1 U573 ( .A1(n706), .A2(n574), .ZN(n464) );
  NAND2_X1 U574 ( .A1(G953), .A2(G902), .ZN(n572) );
  NOR2_X1 U575 ( .A1(G900), .A2(n572), .ZN(n461) );
  NAND2_X1 U576 ( .A1(n706), .A2(n461), .ZN(n462) );
  XNOR2_X1 U577 ( .A(n462), .B(KEYINPUT108), .ZN(n463) );
  AND2_X1 U578 ( .A1(n464), .A2(n463), .ZN(n525) );
  XNOR2_X1 U579 ( .A(n466), .B(n465), .ZN(n508) );
  XNOR2_X1 U580 ( .A(n468), .B(n467), .ZN(n470) );
  NAND2_X1 U581 ( .A1(n481), .A2(G210), .ZN(n469) );
  XOR2_X1 U582 ( .A(n470), .B(n469), .Z(n471) );
  XNOR2_X1 U583 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U584 ( .A(n508), .B(n473), .ZN(n623) );
  NAND2_X1 U585 ( .A1(G214), .A2(n518), .ZN(n692) );
  NAND2_X1 U586 ( .A1(n588), .A2(n692), .ZN(n474) );
  XNOR2_X1 U587 ( .A(n474), .B(KEYINPUT30), .ZN(n475) );
  XNOR2_X1 U588 ( .A(G113), .B(n476), .ZN(n477) );
  XNOR2_X1 U589 ( .A(n479), .B(n478), .ZN(n480) );
  NAND2_X1 U590 ( .A1(G214), .A2(n481), .ZN(n482) );
  XNOR2_X1 U591 ( .A(n483), .B(n482), .ZN(n484) );
  INV_X1 U592 ( .A(n733), .ZN(n485) );
  NAND2_X1 U593 ( .A1(n631), .A2(n499), .ZN(n489) );
  XOR2_X1 U594 ( .A(KEYINPUT104), .B(KEYINPUT13), .Z(n487) );
  XNOR2_X1 U595 ( .A(KEYINPUT103), .B(G475), .ZN(n486) );
  XNOR2_X1 U596 ( .A(n487), .B(n486), .ZN(n488) );
  NAND2_X1 U597 ( .A1(G217), .A2(n490), .ZN(n491) );
  XNOR2_X1 U598 ( .A(n492), .B(n491), .ZN(n498) );
  INV_X1 U599 ( .A(n493), .ZN(n496) );
  XNOR2_X1 U600 ( .A(KEYINPUT9), .B(n494), .ZN(n495) );
  XNOR2_X1 U601 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U602 ( .A(n498), .B(n497), .ZN(n714) );
  NAND2_X1 U603 ( .A1(n714), .A2(n499), .ZN(n501) );
  INV_X1 U604 ( .A(G478), .ZN(n500) );
  XNOR2_X1 U605 ( .A(n501), .B(n500), .ZN(n545) );
  NOR2_X1 U606 ( .A1(n544), .A2(n545), .ZN(n597) );
  INV_X1 U607 ( .A(n502), .ZN(n506) );
  XNOR2_X1 U608 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U609 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U610 ( .A(n508), .B(n507), .ZN(n728) );
  NAND2_X1 U611 ( .A1(G224), .A2(n726), .ZN(n513) );
  XNOR2_X1 U612 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U613 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U614 ( .A(n728), .B(n517), .ZN(n625) );
  NAND2_X1 U615 ( .A1(n625), .A2(n617), .ZN(n521) );
  INV_X1 U616 ( .A(n518), .ZN(n520) );
  INV_X1 U617 ( .A(G210), .ZN(n519) );
  BUF_X1 U618 ( .A(n523), .Z(n524) );
  NOR2_X1 U619 ( .A1(n677), .A2(n525), .ZN(n526) );
  XOR2_X1 U620 ( .A(KEYINPUT72), .B(n526), .Z(n527) );
  NAND2_X1 U621 ( .A1(n588), .A2(n551), .ZN(n528) );
  XNOR2_X1 U622 ( .A(n529), .B(KEYINPUT19), .ZN(n578) );
  NAND2_X1 U623 ( .A1(n530), .A2(n578), .ZN(n657) );
  NAND2_X1 U624 ( .A1(n657), .A2(KEYINPUT47), .ZN(n535) );
  INV_X1 U625 ( .A(n545), .ZN(n531) );
  NAND2_X1 U626 ( .A1(n697), .A2(KEYINPUT47), .ZN(n533) );
  XNOR2_X1 U627 ( .A(KEYINPUT90), .B(n533), .ZN(n534) );
  NOR2_X1 U628 ( .A1(KEYINPUT47), .A2(n697), .ZN(n537) );
  XNOR2_X1 U629 ( .A(KEYINPUT81), .B(n537), .ZN(n538) );
  XNOR2_X1 U630 ( .A(n539), .B(KEYINPUT80), .ZN(n559) );
  NAND2_X1 U631 ( .A1(n540), .A2(n693), .ZN(n542) );
  XOR2_X1 U632 ( .A(KEYINPUT75), .B(KEYINPUT39), .Z(n541) );
  XNOR2_X2 U633 ( .A(n542), .B(n541), .ZN(n561) );
  INV_X1 U634 ( .A(n658), .ZN(n660) );
  NAND2_X1 U635 ( .A1(n693), .A2(n692), .ZN(n696) );
  NAND2_X1 U636 ( .A1(n545), .A2(n544), .ZN(n695) );
  NOR2_X1 U637 ( .A1(n696), .A2(n695), .ZN(n546) );
  XNOR2_X1 U638 ( .A(n546), .B(KEYINPUT41), .ZN(n690) );
  NOR2_X1 U639 ( .A1(n547), .A2(n690), .ZN(n549) );
  XNOR2_X1 U640 ( .A(KEYINPUT115), .B(KEYINPUT42), .ZN(n548) );
  XNOR2_X1 U641 ( .A(n549), .B(n548), .ZN(n745) );
  NOR2_X1 U642 ( .A1(n607), .A2(n658), .ZN(n550) );
  NAND2_X1 U643 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U644 ( .A(n552), .B(KEYINPUT109), .ZN(n553) );
  NAND2_X1 U645 ( .A1(n553), .A2(n692), .ZN(n562) );
  NOR2_X1 U646 ( .A1(n562), .A2(n567), .ZN(n554) );
  XOR2_X1 U647 ( .A(KEYINPUT36), .B(n554), .Z(n556) );
  XNOR2_X1 U648 ( .A(n563), .B(KEYINPUT96), .ZN(n601) );
  OR2_X1 U649 ( .A1(n556), .A2(n601), .ZN(n666) );
  NAND2_X1 U650 ( .A1(n561), .A2(n662), .ZN(n667) );
  INV_X1 U651 ( .A(n667), .ZN(n569) );
  XNOR2_X1 U652 ( .A(KEYINPUT110), .B(n562), .ZN(n564) );
  NOR2_X1 U653 ( .A1(n564), .A2(n682), .ZN(n566) );
  XNOR2_X1 U654 ( .A(KEYINPUT111), .B(KEYINPUT43), .ZN(n565) );
  XNOR2_X1 U655 ( .A(n566), .B(n565), .ZN(n568) );
  AND2_X1 U656 ( .A1(n568), .A2(n567), .ZN(n668) );
  NOR2_X1 U657 ( .A1(n569), .A2(n668), .ZN(n570) );
  INV_X1 U658 ( .A(n706), .ZN(n576) );
  NOR2_X1 U659 ( .A1(G898), .A2(n572), .ZN(n573) );
  NOR2_X1 U660 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U661 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U662 ( .A1(n578), .A2(n577), .ZN(n580) );
  INV_X1 U663 ( .A(n695), .ZN(n581) );
  AND2_X1 U664 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U665 ( .A1(n593), .A2(n583), .ZN(n586) );
  INV_X1 U666 ( .A(KEYINPUT22), .ZN(n584) );
  XNOR2_X1 U667 ( .A(n609), .B(KEYINPUT107), .ZN(n587) );
  INV_X1 U668 ( .A(n588), .ZN(n681) );
  NAND2_X1 U669 ( .A1(n589), .A2(n681), .ZN(n652) );
  INV_X1 U670 ( .A(n652), .ZN(n598) );
  XNOR2_X1 U671 ( .A(KEYINPUT33), .B(KEYINPUT74), .ZN(n591) );
  XNOR2_X1 U672 ( .A(n592), .B(n591), .ZN(n672) );
  INV_X1 U673 ( .A(n593), .ZN(n594) );
  XOR2_X1 U674 ( .A(KEYINPUT34), .B(KEYINPUT85), .Z(n595) );
  XNOR2_X1 U675 ( .A(KEYINPUT76), .B(n595), .ZN(n596) );
  XNOR2_X1 U676 ( .A(KEYINPUT87), .B(n607), .ZN(n599) );
  NOR2_X1 U677 ( .A1(n600), .A2(n599), .ZN(n603) );
  NAND2_X1 U678 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U679 ( .A(n604), .B(KEYINPUT32), .ZN(n605) );
  XNOR2_X1 U680 ( .A(KEYINPUT86), .B(n605), .ZN(n743) );
  NAND2_X1 U681 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U682 ( .A(KEYINPUT106), .B(n610), .ZN(n747) );
  NOR2_X1 U683 ( .A1(n681), .A2(n611), .ZN(n687) );
  NAND2_X1 U684 ( .A1(n593), .A2(n687), .ZN(n612) );
  XNOR2_X1 U685 ( .A(n612), .B(KEYINPUT31), .ZN(n663) );
  NAND2_X1 U686 ( .A1(n681), .A2(n593), .ZN(n614) );
  NOR2_X1 U687 ( .A1(n614), .A2(n613), .ZN(n647) );
  NOR2_X1 U688 ( .A1(n663), .A2(n647), .ZN(n615) );
  NOR2_X1 U689 ( .A1(n615), .A2(n697), .ZN(n616) );
  NAND2_X1 U690 ( .A1(n721), .A2(KEYINPUT2), .ZN(n621) );
  BUF_X1 U691 ( .A(n619), .Z(n620) );
  NAND2_X1 U692 ( .A1(n717), .A2(G210), .ZN(n627) );
  XOR2_X1 U693 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n624) );
  XNOR2_X1 U694 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U695 ( .A(n627), .B(n626), .ZN(n628) );
  INV_X1 U696 ( .A(n720), .ZN(n641) );
  NAND2_X1 U697 ( .A1(n628), .A2(n641), .ZN(n630) );
  XNOR2_X1 U698 ( .A(KEYINPUT93), .B(KEYINPUT56), .ZN(n629) );
  XNOR2_X1 U699 ( .A(n630), .B(n629), .ZN(G51) );
  NAND2_X1 U700 ( .A1(n717), .A2(G475), .ZN(n633) );
  XOR2_X1 U701 ( .A(KEYINPUT59), .B(n631), .Z(n632) );
  XNOR2_X1 U702 ( .A(n633), .B(n632), .ZN(n634) );
  NAND2_X1 U703 ( .A1(n634), .A2(n641), .ZN(n636) );
  INV_X1 U704 ( .A(KEYINPUT60), .ZN(n635) );
  XNOR2_X1 U705 ( .A(n636), .B(n635), .ZN(G60) );
  NAND2_X1 U706 ( .A1(n717), .A2(G469), .ZN(n640) );
  XNOR2_X1 U707 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n637) );
  XNOR2_X1 U708 ( .A(n638), .B(n637), .ZN(n639) );
  XNOR2_X1 U709 ( .A(n640), .B(n639), .ZN(n642) );
  NAND2_X1 U710 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U711 ( .A(n643), .B(KEYINPUT123), .ZN(G54) );
  XNOR2_X1 U712 ( .A(n644), .B(G143), .ZN(G45) );
  NAND2_X1 U713 ( .A1(n647), .A2(n660), .ZN(n645) );
  XNOR2_X1 U714 ( .A(n645), .B(KEYINPUT116), .ZN(n646) );
  XNOR2_X1 U715 ( .A(G104), .B(n646), .ZN(G6) );
  XOR2_X1 U716 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n649) );
  NAND2_X1 U717 ( .A1(n647), .A2(n662), .ZN(n648) );
  XNOR2_X1 U718 ( .A(n649), .B(n648), .ZN(n651) );
  XOR2_X1 U719 ( .A(G107), .B(KEYINPUT117), .Z(n650) );
  XNOR2_X1 U720 ( .A(n651), .B(n650), .ZN(G9) );
  XNOR2_X1 U721 ( .A(G110), .B(KEYINPUT118), .ZN(n653) );
  XNOR2_X1 U722 ( .A(n653), .B(n652), .ZN(G12) );
  NOR2_X1 U723 ( .A1(n657), .A2(n654), .ZN(n656) );
  XNOR2_X1 U724 ( .A(G128), .B(KEYINPUT29), .ZN(n655) );
  XNOR2_X1 U725 ( .A(n656), .B(n655), .ZN(G30) );
  NOR2_X1 U726 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U727 ( .A(G146), .B(n659), .Z(G48) );
  NAND2_X1 U728 ( .A1(n663), .A2(n660), .ZN(n661) );
  XNOR2_X1 U729 ( .A(n661), .B(G113), .ZN(G15) );
  NAND2_X1 U730 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U731 ( .A(n664), .B(G116), .ZN(G18) );
  XOR2_X1 U732 ( .A(G125), .B(KEYINPUT37), .Z(n665) );
  XNOR2_X1 U733 ( .A(n666), .B(n665), .ZN(G27) );
  XNOR2_X1 U734 ( .A(G134), .B(n667), .ZN(G36) );
  XOR2_X1 U735 ( .A(G140), .B(n668), .Z(G42) );
  NAND2_X1 U736 ( .A1(n721), .A2(n669), .ZN(n670) );
  NAND2_X1 U737 ( .A1(n670), .A2(KEYINPUT88), .ZN(n671) );
  XOR2_X1 U738 ( .A(n671), .B(n432), .Z(n676) );
  NOR2_X1 U739 ( .A1(n672), .A2(n690), .ZN(n673) );
  XNOR2_X1 U740 ( .A(KEYINPUT122), .B(n673), .ZN(n674) );
  NOR2_X1 U741 ( .A1(G953), .A2(n674), .ZN(n675) );
  NAND2_X1 U742 ( .A1(n676), .A2(n675), .ZN(n711) );
  INV_X1 U743 ( .A(n677), .ZN(n678) );
  XNOR2_X1 U744 ( .A(n679), .B(KEYINPUT49), .ZN(n680) );
  NAND2_X1 U745 ( .A1(n681), .A2(n680), .ZN(n685) );
  NOR2_X1 U746 ( .A1(n590), .A2(n682), .ZN(n683) );
  XNOR2_X1 U747 ( .A(n683), .B(KEYINPUT50), .ZN(n684) );
  NOR2_X1 U748 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U749 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U750 ( .A(KEYINPUT51), .B(n688), .Z(n689) );
  NOR2_X1 U751 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U752 ( .A(KEYINPUT119), .B(n691), .ZN(n704) );
  NOR2_X1 U753 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U754 ( .A1(n695), .A2(n694), .ZN(n700) );
  NOR2_X1 U755 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U756 ( .A(n698), .B(KEYINPUT120), .ZN(n699) );
  NOR2_X1 U757 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U758 ( .A1(n672), .A2(n701), .ZN(n702) );
  XNOR2_X1 U759 ( .A(KEYINPUT121), .B(n702), .ZN(n703) );
  NAND2_X1 U760 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U761 ( .A(KEYINPUT52), .B(n705), .ZN(n707) );
  NAND2_X1 U762 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U763 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U764 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U765 ( .A(KEYINPUT53), .B(n712), .ZN(G75) );
  NAND2_X1 U766 ( .A1(n717), .A2(G478), .ZN(n713) );
  XOR2_X1 U767 ( .A(n714), .B(n713), .Z(n715) );
  NOR2_X1 U768 ( .A1(n720), .A2(n715), .ZN(G63) );
  NAND2_X1 U769 ( .A1(n717), .A2(G217), .ZN(n718) );
  XNOR2_X1 U770 ( .A(n716), .B(n718), .ZN(n719) );
  NOR2_X1 U771 ( .A1(n720), .A2(n719), .ZN(G66) );
  NAND2_X1 U772 ( .A1(n726), .A2(n721), .ZN(n725) );
  NAND2_X1 U773 ( .A1(G953), .A2(G224), .ZN(n722) );
  XNOR2_X1 U774 ( .A(KEYINPUT61), .B(n722), .ZN(n723) );
  NAND2_X1 U775 ( .A1(n723), .A2(G898), .ZN(n724) );
  NAND2_X1 U776 ( .A1(n725), .A2(n724), .ZN(n730) );
  NOR2_X1 U777 ( .A1(G898), .A2(n726), .ZN(n727) );
  NOR2_X1 U778 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U779 ( .A(n730), .B(n729), .ZN(n731) );
  XNOR2_X1 U780 ( .A(KEYINPUT124), .B(n731), .ZN(G69) );
  XNOR2_X1 U781 ( .A(n732), .B(n733), .ZN(n736) );
  NOR2_X1 U782 ( .A1(n734), .A2(G953), .ZN(n735) );
  XNOR2_X1 U783 ( .A(n735), .B(KEYINPUT125), .ZN(n741) );
  XOR2_X1 U784 ( .A(G227), .B(n736), .Z(n737) );
  XNOR2_X1 U785 ( .A(n737), .B(KEYINPUT126), .ZN(n738) );
  NAND2_X1 U786 ( .A1(n738), .A2(G900), .ZN(n739) );
  NAND2_X1 U787 ( .A1(G953), .A2(n739), .ZN(n740) );
  NAND2_X1 U788 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U789 ( .A(KEYINPUT127), .B(n742), .Z(G72) );
  XNOR2_X1 U790 ( .A(G119), .B(n743), .ZN(G21) );
  XOR2_X1 U791 ( .A(G122), .B(n744), .Z(G24) );
  XNOR2_X1 U792 ( .A(G137), .B(n745), .ZN(G39) );
  XNOR2_X1 U793 ( .A(n746), .B(G131), .ZN(G33) );
  XNOR2_X1 U794 ( .A(G101), .B(n747), .ZN(G3) );
endmodule

