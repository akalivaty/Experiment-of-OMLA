//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 0 1 1 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n796, new_n798, new_n799, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n986, new_n987, new_n988, new_n989, new_n990, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1030, new_n1031;
  INV_X1    g000(.A(KEYINPUT18), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT17), .ZN(new_n203));
  XOR2_X1   g002(.A(G43gat), .B(G50gat), .Z(new_n204));
  INV_X1    g003(.A(KEYINPUT15), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT93), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G43gat), .B(G50gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT15), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT91), .B(G29gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(KEYINPUT92), .B(G36gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(G29gat), .A2(G36gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT14), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n214));
  AOI22_X1  g013(.A1(new_n209), .A2(new_n210), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AND3_X1   g014(.A1(new_n206), .A2(new_n208), .A3(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n208), .B1(new_n206), .B2(new_n215), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n203), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n206), .A2(new_n215), .ZN(new_n219));
  INV_X1    g018(.A(new_n208), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n206), .A2(new_n215), .A3(new_n208), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(KEYINPUT17), .A3(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G15gat), .B(G22gat), .ZN(new_n224));
  INV_X1    g023(.A(G1gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT16), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(G1gat), .B2(new_n224), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G8gat), .ZN(new_n229));
  INV_X1    g028(.A(G8gat), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n227), .B(new_n230), .C1(G1gat), .C2(new_n224), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n218), .A2(new_n223), .A3(new_n232), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n221), .A2(new_n222), .B1(new_n229), .B2(new_n231), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G229gat), .A2(G233gat), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n202), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n221), .A2(new_n222), .A3(new_n229), .A4(new_n231), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT94), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT94), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n232), .A2(new_n242), .A3(new_n221), .A4(new_n222), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n241), .A2(new_n243), .A3(new_n235), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n237), .B(KEYINPUT13), .Z(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n233), .A2(new_n235), .A3(KEYINPUT18), .A4(new_n237), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n239), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G113gat), .B(G141gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(G197gat), .ZN(new_n250));
  XOR2_X1   g049(.A(KEYINPUT11), .B(G169gat), .Z(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(KEYINPUT12), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n248), .A2(KEYINPUT90), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n253), .B1(new_n248), .B2(KEYINPUT90), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G197gat), .B(G204gat), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT22), .ZN(new_n259));
  INV_X1    g058(.A(G211gat), .ZN(new_n260));
  INV_X1    g059(.A(G218gat), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G211gat), .B(G218gat), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(new_n258), .A3(new_n262), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G226gat), .A2(G233gat), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  AND2_X1   g070(.A1(G183gat), .A2(G190gat), .ZN(new_n272));
  NOR2_X1   g071(.A1(G183gat), .A2(G190gat), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT24), .ZN(new_n274));
  NOR3_X1   g073(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT23), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n276), .B1(G169gat), .B2(G176gat), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n274), .A2(G183gat), .A3(G190gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n275), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT65), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT64), .ZN(new_n283));
  INV_X1    g082(.A(G169gat), .ZN(new_n284));
  INV_X1    g083(.A(G176gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n286), .A2(KEYINPUT23), .A3(new_n287), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n281), .A2(new_n282), .A3(KEYINPUT25), .A4(new_n288), .ZN(new_n289));
  AOI22_X1  g088(.A1(new_n272), .A2(new_n274), .B1(G169gat), .B2(G176gat), .ZN(new_n290));
  INV_X1    g089(.A(G183gat), .ZN(new_n291));
  INV_X1    g090(.A(G190gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n293), .A2(KEYINPUT24), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n290), .A2(new_n295), .A3(new_n277), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n288), .A2(KEYINPUT25), .ZN(new_n297));
  OAI21_X1  g096(.A(KEYINPUT65), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n284), .A2(new_n285), .A3(KEYINPUT23), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n290), .A2(new_n295), .A3(new_n277), .A4(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT25), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n289), .A2(new_n298), .A3(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n286), .A2(new_n287), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n304), .B(new_n279), .C1(new_n305), .C2(KEYINPUT26), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT27), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT27), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G183gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n307), .A2(new_n309), .A3(new_n292), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT28), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n311), .A2(KEYINPUT66), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n272), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n307), .A2(new_n309), .ZN(new_n314));
  XNOR2_X1  g113(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n314), .A2(new_n315), .A3(new_n292), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n306), .A2(new_n313), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n303), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT29), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n271), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  AND3_X1   g119(.A1(new_n306), .A2(new_n313), .A3(new_n316), .ZN(new_n321));
  AND3_X1   g120(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n322), .A2(KEYINPUT25), .A3(new_n295), .A4(new_n288), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n323), .A2(KEYINPUT65), .B1(new_n301), .B2(new_n300), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n321), .B1(new_n324), .B2(new_n289), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n325), .A2(new_n270), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n269), .B1(new_n320), .B2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G8gat), .B(G36gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(KEYINPUT73), .ZN(new_n329));
  XNOR2_X1  g128(.A(G64gat), .B(G92gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n329), .B(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n270), .B1(new_n325), .B2(KEYINPUT29), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n318), .A2(new_n271), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(new_n333), .A3(new_n268), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n327), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT30), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n327), .A2(new_n334), .ZN(new_n338));
  INV_X1    g137(.A(new_n331), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n327), .A2(KEYINPUT30), .A3(new_n334), .A4(new_n331), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT89), .B(KEYINPUT35), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n337), .A2(new_n340), .A3(new_n341), .A4(new_n342), .ZN(new_n343));
  AND2_X1   g142(.A1(G113gat), .A2(G120gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(G113gat), .A2(G120gat), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT1), .ZN(new_n347));
  OR2_X1    g146(.A1(new_n347), .A2(KEYINPUT69), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(KEYINPUT69), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n346), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G127gat), .B(G134gat), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT68), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n352), .B1(new_n344), .B2(new_n345), .ZN(new_n353));
  INV_X1    g152(.A(G113gat), .ZN(new_n354));
  INV_X1    g153(.A(G120gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G113gat), .A2(G120gat), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n356), .A2(KEYINPUT68), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n353), .A2(new_n358), .A3(new_n347), .ZN(new_n359));
  INV_X1    g158(.A(G127gat), .ZN(new_n360));
  NOR3_X1   g159(.A1(new_n360), .A2(KEYINPUT67), .A3(G134gat), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n361), .B1(new_n351), .B2(KEYINPUT67), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n350), .A2(new_n351), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT75), .ZN(new_n364));
  AND2_X1   g163(.A1(G155gat), .A2(G162gat), .ZN(new_n365));
  NOR2_X1   g164(.A1(G155gat), .A2(G162gat), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(G155gat), .ZN(new_n368));
  INV_X1    g167(.A(G162gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(G155gat), .A2(G162gat), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n370), .A2(KEYINPUT75), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(KEYINPUT2), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT76), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT76), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n371), .A2(new_n376), .A3(KEYINPUT2), .ZN(new_n377));
  AND2_X1   g176(.A1(G141gat), .A2(G148gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(G141gat), .A2(G148gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n375), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n365), .A2(new_n366), .ZN(new_n382));
  XNOR2_X1  g181(.A(G141gat), .B(G148gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI22_X1  g183(.A1(new_n373), .A2(new_n381), .B1(new_n384), .B2(new_n374), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n363), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT4), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  XOR2_X1   g187(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n363), .A2(new_n385), .A3(new_n390), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT5), .ZN(new_n393));
  NAND2_X1  g192(.A1(G225gat), .A2(G233gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n359), .A2(new_n362), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n346), .A2(new_n351), .A3(new_n348), .A4(new_n349), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT77), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT77), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n395), .A2(new_n399), .A3(new_n396), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n376), .B1(new_n371), .B2(KEYINPUT2), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n383), .A2(new_n401), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n402), .A2(new_n377), .B1(new_n367), .B2(new_n372), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n380), .B(new_n374), .C1(new_n365), .C2(new_n366), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT3), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n381), .A2(new_n373), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT3), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n407), .A2(new_n408), .A3(new_n404), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n398), .A2(new_n400), .A3(new_n406), .A4(new_n409), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n392), .A2(new_n393), .A3(new_n394), .A4(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n385), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n398), .A2(new_n400), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n386), .ZN(new_n414));
  INV_X1    g213(.A(new_n394), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n393), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT79), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n363), .A2(KEYINPUT4), .A3(new_n385), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n386), .A2(new_n389), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n410), .A2(new_n394), .A3(new_n418), .A4(new_n419), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n416), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n417), .B1(new_n416), .B2(new_n420), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n411), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  XOR2_X1   g222(.A(G1gat), .B(G29gat), .Z(new_n424));
  XNOR2_X1  g223(.A(G57gat), .B(G85gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n423), .A2(new_n428), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n395), .A2(new_n399), .A3(new_n396), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n399), .B1(new_n395), .B2(new_n396), .ZN(new_n431));
  NOR3_X1   g230(.A1(new_n430), .A2(new_n431), .A3(new_n385), .ZN(new_n432));
  INV_X1    g231(.A(new_n386), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n415), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n434), .A2(new_n420), .A3(KEYINPUT5), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT79), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n416), .A2(new_n417), .A3(new_n420), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n428), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n411), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT6), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n429), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n439), .B1(new_n438), .B2(new_n411), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT6), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n343), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n268), .A2(new_n319), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n385), .B1(new_n446), .B2(new_n408), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(KEYINPUT85), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n268), .B1(new_n409), .B2(new_n319), .ZN(new_n449));
  NAND2_X1  g248(.A1(G228gat), .A2(G233gat), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT84), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n266), .A2(KEYINPUT82), .A3(new_n267), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT82), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n264), .A2(new_n258), .A3(new_n455), .A4(new_n262), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n456), .A2(new_n319), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT3), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  OAI22_X1  g257(.A1(new_n449), .A2(KEYINPUT83), .B1(new_n458), .B2(new_n385), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT29), .B1(new_n385), .B2(new_n408), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT83), .ZN(new_n461));
  NOR3_X1   g260(.A1(new_n460), .A2(new_n461), .A3(new_n268), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n453), .B(new_n450), .C1(new_n459), .C2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n461), .B1(new_n460), .B2(new_n268), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n454), .A2(new_n457), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n412), .B1(new_n466), .B2(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n449), .A2(KEYINPUT83), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n453), .B1(new_n469), .B2(new_n450), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n452), .B1(new_n464), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(G22gat), .ZN(new_n472));
  INV_X1    g271(.A(G22gat), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n473), .B(new_n452), .C1(new_n464), .C2(new_n470), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G78gat), .B(G106gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(KEYINPUT31), .B(G50gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n476), .B(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n472), .A2(new_n474), .A3(new_n478), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n318), .A2(new_n363), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n325), .A2(new_n397), .ZN(new_n484));
  NAND2_X1  g283(.A1(G227gat), .A2(G233gat), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n483), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT32), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT33), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  XOR2_X1   g289(.A(G71gat), .B(G99gat), .Z(new_n491));
  XNOR2_X1  g290(.A(G15gat), .B(G43gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n491), .B(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n488), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT70), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n489), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n496), .B1(new_n495), .B2(new_n493), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n487), .A2(KEYINPUT32), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n486), .B1(new_n483), .B2(new_n484), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT34), .B1(new_n486), .B2(KEYINPUT71), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n500), .B(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT72), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n500), .A2(new_n501), .ZN(new_n505));
  OR2_X1    g304(.A1(new_n500), .A2(new_n501), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n494), .A2(new_n505), .A3(new_n506), .A4(new_n498), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n503), .A2(new_n504), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n499), .A2(KEYINPUT72), .A3(new_n502), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n445), .A2(new_n482), .A3(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT6), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n429), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n440), .B1(new_n421), .B2(new_n422), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(new_n512), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT81), .B1(new_n515), .B2(new_n443), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT81), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n429), .A2(new_n441), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n513), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n503), .A2(new_n507), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n472), .A2(new_n474), .A3(new_n478), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n478), .B1(new_n472), .B2(new_n474), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n340), .A2(new_n341), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT74), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n340), .A2(KEYINPUT74), .A3(new_n341), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n526), .A2(new_n337), .A3(new_n527), .ZN(new_n528));
  NOR3_X1   g327(.A1(new_n519), .A2(new_n523), .A3(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT35), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n511), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n482), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n532), .B1(new_n519), .B2(new_n528), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT88), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n327), .A2(new_n534), .A3(new_n334), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT37), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n327), .A2(new_n534), .A3(new_n334), .A4(KEYINPUT37), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT38), .B1(new_n539), .B2(new_n331), .ZN(new_n540));
  INV_X1    g339(.A(new_n335), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n331), .B1(new_n537), .B2(new_n538), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT38), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n540), .A2(new_n544), .A3(new_n444), .A4(new_n442), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n413), .A2(new_n394), .A3(new_n386), .ZN(new_n546));
  AOI21_X1  g345(.A(KEYINPUT86), .B1(new_n546), .B2(KEYINPUT39), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n546), .A2(KEYINPUT86), .A3(KEYINPUT39), .ZN(new_n549));
  INV_X1    g348(.A(new_n410), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n388), .A2(new_n391), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n415), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n548), .A2(new_n549), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n394), .B1(new_n392), .B2(new_n410), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT39), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n428), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT40), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n337), .A2(new_n340), .A3(new_n341), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n553), .A2(new_n556), .A3(KEYINPUT40), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n429), .A2(new_n559), .A3(new_n560), .A4(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT87), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n439), .B1(new_n552), .B2(KEYINPUT39), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n554), .A2(new_n547), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n564), .B1(new_n565), .B2(new_n549), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n423), .A2(new_n428), .B1(new_n566), .B2(KEYINPUT40), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT87), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n567), .A2(new_n568), .A3(new_n560), .A4(new_n559), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n545), .A2(new_n482), .A3(new_n563), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n520), .A2(KEYINPUT36), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n571), .B1(new_n510), .B2(KEYINPUT36), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n533), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n257), .B1(new_n531), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT103), .ZN(new_n575));
  XNOR2_X1  g374(.A(G120gat), .B(G148gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(G176gat), .B(G204gat), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n576), .B(new_n577), .Z(new_n578));
  NOR2_X1   g377(.A1(G57gat), .A2(G64gat), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G57gat), .A2(G64gat), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n580), .A2(KEYINPUT95), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT95), .ZN(new_n583));
  INV_X1    g382(.A(new_n581), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n583), .B1(new_n584), .B2(new_n579), .ZN(new_n585));
  XNOR2_X1  g384(.A(G71gat), .B(G78gat), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n582), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT96), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n586), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n584), .A2(new_n579), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(KEYINPUT9), .ZN(new_n594));
  AOI22_X1  g393(.A1(new_n587), .A2(new_n591), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT99), .ZN(new_n596));
  OR2_X1    g395(.A1(G99gat), .A2(G106gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(G99gat), .A2(G106gat), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n597), .A2(new_n596), .A3(new_n598), .ZN(new_n600));
  INV_X1    g399(.A(G85gat), .ZN(new_n601));
  INV_X1    g400(.A(G92gat), .ZN(new_n602));
  AOI22_X1  g401(.A1(KEYINPUT8), .A2(new_n598), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(KEYINPUT98), .A2(G85gat), .A3(G92gat), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT7), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g406(.A1(KEYINPUT98), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n599), .B1(new_n604), .B2(new_n609), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n607), .A2(new_n608), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n597), .A2(new_n598), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT99), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n611), .A2(new_n613), .A3(new_n600), .A4(new_n603), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n595), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT10), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n594), .A2(new_n592), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n582), .A2(new_n585), .A3(new_n586), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n618), .B1(new_n619), .B2(new_n590), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n620), .A2(new_n610), .A3(new_n614), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n616), .A2(new_n617), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(KEYINPUT102), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT102), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n616), .A2(new_n621), .A3(new_n624), .A4(new_n617), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n610), .A2(new_n614), .ZN(new_n626));
  NOR3_X1   g425(.A1(new_n626), .A2(new_n617), .A3(new_n620), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n623), .A2(new_n625), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G230gat), .A2(G233gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n616), .A2(new_n621), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n632), .A2(new_n630), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n578), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n630), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n627), .B1(new_n622), .B2(KEYINPUT102), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n636), .B1(new_n637), .B2(new_n625), .ZN(new_n638));
  INV_X1    g437(.A(new_n578), .ZN(new_n639));
  NOR3_X1   g438(.A1(new_n638), .A2(new_n633), .A3(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n575), .B1(new_n635), .B2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n631), .A2(new_n634), .A3(new_n578), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n639), .B1(new_n638), .B2(new_n633), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n642), .A2(new_n643), .A3(KEYINPUT103), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n218), .A2(new_n223), .A3(new_n626), .ZN(new_n647));
  AOI22_X1  g446(.A1(new_n221), .A2(new_n222), .B1(new_n610), .B2(new_n614), .ZN(new_n648));
  NAND2_X1  g447(.A1(G232gat), .A2(G233gat), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT41), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n648), .A2(KEYINPUT100), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT100), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n615), .B1(new_n216), .B2(new_n217), .ZN(new_n654));
  INV_X1    g453(.A(new_n651), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n647), .B1(new_n652), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT97), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n659), .ZN(new_n661));
  OAI211_X1 g460(.A(new_n647), .B(new_n661), .C1(new_n652), .C2(new_n656), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(G190gat), .B(G218gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(G134gat), .B(G162gat), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n664), .B(new_n665), .Z(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n660), .A2(new_n662), .A3(new_n666), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n595), .A2(KEYINPUT21), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT21), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n620), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(G127gat), .B(G155gat), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  OAI211_X1 g476(.A(new_n232), .B(new_n671), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n677), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n232), .B1(new_n672), .B2(new_n620), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n679), .A2(new_n680), .A3(new_n675), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n682));
  NAND2_X1  g481(.A1(G231gat), .A2(G233gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(G183gat), .B(G211gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n678), .A2(new_n681), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n686), .B1(new_n678), .B2(new_n681), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(KEYINPUT101), .B1(new_n670), .B2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT101), .ZN(new_n692));
  AOI211_X1 g491(.A(new_n692), .B(new_n689), .C1(new_n668), .C2(new_n669), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n646), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n574), .A2(new_n694), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n515), .A2(new_n443), .A3(KEYINPUT81), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n517), .B1(new_n429), .B2(new_n441), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n444), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(new_n225), .ZN(G1324gat));
  INV_X1    g499(.A(new_n560), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n695), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g501(.A(KEYINPUT16), .B(G8gat), .Z(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n704), .B1(new_n230), .B2(new_n702), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT42), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT42), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(G1325gat));
  OAI21_X1  g508(.A(G15gat), .B1(new_n695), .B2(new_n572), .ZN(new_n710));
  INV_X1    g509(.A(new_n510), .ZN(new_n711));
  OR2_X1    g510(.A1(new_n711), .A2(G15gat), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n710), .B1(new_n695), .B2(new_n712), .ZN(G1326gat));
  NAND3_X1  g512(.A1(new_n574), .A2(new_n532), .A3(new_n694), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT104), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT43), .B(G22gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1327gat));
  NOR2_X1   g516(.A1(new_n646), .A2(new_n690), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n256), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT106), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n670), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n533), .A2(new_n570), .A3(new_n572), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n445), .A2(new_n482), .A3(new_n510), .ZN(new_n724));
  INV_X1    g523(.A(new_n528), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n503), .A2(new_n507), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n726), .B1(new_n480), .B2(new_n481), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n698), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n724), .B1(new_n728), .B2(KEYINPUT35), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n722), .B1(new_n723), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(KEYINPUT44), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n668), .A2(KEYINPUT107), .A3(new_n669), .ZN(new_n732));
  AOI21_X1  g531(.A(KEYINPUT107), .B1(new_n668), .B2(new_n669), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n736), .B1(new_n531), .B2(new_n573), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n721), .B1(new_n731), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n519), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n209), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n718), .A2(new_n722), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n742), .B(KEYINPUT105), .Z(new_n743));
  NOR2_X1   g542(.A1(new_n698), .A2(new_n209), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n574), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT45), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n741), .A2(new_n746), .ZN(G1328gat));
  NAND2_X1  g546(.A1(new_n739), .A2(new_n560), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n210), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n701), .A2(new_n210), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n574), .A2(new_n743), .A3(new_n750), .ZN(new_n751));
  XOR2_X1   g550(.A(new_n751), .B(KEYINPUT46), .Z(new_n752));
  NAND2_X1  g551(.A1(new_n749), .A2(new_n752), .ZN(G1329gat));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n754));
  XNOR2_X1  g553(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n755));
  INV_X1    g554(.A(G43gat), .ZN(new_n756));
  INV_X1    g555(.A(new_n572), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n756), .B1(new_n739), .B2(new_n757), .ZN(new_n758));
  AND4_X1   g557(.A1(new_n756), .A2(new_n574), .A3(new_n510), .A4(new_n743), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n754), .B(new_n755), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n755), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n531), .A2(new_n573), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n735), .B1(new_n762), .B2(new_n722), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n757), .B(new_n720), .C1(new_n763), .C2(new_n737), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n759), .B1(new_n764), .B2(G43gat), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n761), .B1(new_n765), .B2(KEYINPUT108), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n760), .A2(new_n766), .ZN(G1330gat));
  NAND2_X1  g566(.A1(new_n731), .A2(new_n738), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n768), .A2(G50gat), .A3(new_n532), .A4(new_n720), .ZN(new_n769));
  OR2_X1    g568(.A1(KEYINPUT110), .A2(KEYINPUT48), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n574), .A2(new_n532), .A3(new_n743), .ZN(new_n771));
  INV_X1    g570(.A(G50gat), .ZN(new_n772));
  AOI22_X1  g571(.A1(new_n771), .A2(new_n772), .B1(KEYINPUT110), .B2(KEYINPUT48), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n769), .A2(new_n770), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n770), .B1(new_n769), .B2(new_n773), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(G1331gat));
  NOR4_X1   g575(.A1(new_n691), .A2(new_n693), .A3(new_n645), .A4(new_n256), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n762), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n519), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT112), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n779), .B(new_n780), .ZN(new_n781));
  XNOR2_X1  g580(.A(KEYINPUT111), .B(G57gat), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n779), .B(KEYINPUT112), .ZN(new_n784));
  INV_X1    g583(.A(new_n782), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n783), .A2(new_n786), .ZN(G1332gat));
  NAND2_X1  g586(.A1(new_n762), .A2(new_n777), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(new_n701), .ZN(new_n789));
  NOR2_X1   g588(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n790));
  AND2_X1   g589(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n792), .B1(new_n789), .B2(new_n790), .ZN(G1333gat));
  OR3_X1    g592(.A1(new_n788), .A2(G71gat), .A3(new_n711), .ZN(new_n794));
  OAI21_X1  g593(.A(G71gat), .B1(new_n788), .B2(new_n572), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XOR2_X1   g595(.A(new_n796), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g596(.A1(new_n788), .A2(new_n482), .ZN(new_n798));
  XNOR2_X1  g597(.A(KEYINPUT113), .B(G78gat), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n798), .B(new_n799), .ZN(G1335gat));
  NOR3_X1   g599(.A1(new_n645), .A2(new_n256), .A3(new_n690), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n768), .A2(new_n519), .A3(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n256), .A2(new_n690), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n722), .B(new_n803), .C1(new_n723), .C2(new_n729), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n762), .A2(KEYINPUT51), .A3(new_n722), .A4(new_n803), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n519), .A2(new_n601), .A3(new_n646), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(KEYINPUT114), .ZN(new_n811));
  OAI22_X1  g610(.A1(new_n802), .A2(new_n601), .B1(new_n809), .B2(new_n811), .ZN(G1336gat));
  NOR3_X1   g611(.A1(new_n645), .A2(G92gat), .A3(new_n701), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(KEYINPUT115), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT52), .B1(new_n808), .B2(new_n814), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n560), .B(new_n801), .C1(new_n763), .C2(new_n737), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(G92gat), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n804), .A2(new_n819), .A3(KEYINPUT51), .ZN(new_n820));
  AOI21_X1  g619(.A(KEYINPUT51), .B1(new_n804), .B2(new_n819), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AOI22_X1  g621(.A1(new_n822), .A2(new_n814), .B1(G92gat), .B2(new_n816), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n818), .B1(new_n823), .B2(new_n824), .ZN(G1337gat));
  INV_X1    g624(.A(G99gat), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n808), .A2(new_n826), .A3(new_n510), .A4(new_n646), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n768), .A2(new_n757), .A3(new_n801), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n827), .B1(new_n828), .B2(new_n826), .ZN(G1338gat));
  OAI211_X1 g628(.A(new_n532), .B(new_n801), .C1(new_n763), .C2(new_n737), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n830), .A2(G106gat), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n482), .A2(G106gat), .A3(new_n645), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n820), .A2(new_n821), .A3(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT53), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT53), .B1(new_n830), .B2(G106gat), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n837), .B1(new_n808), .B2(new_n832), .ZN(new_n838));
  AOI211_X1 g637(.A(KEYINPUT117), .B(new_n833), .C1(new_n806), .C2(new_n807), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n835), .A2(new_n840), .ZN(G1339gat));
  AND3_X1   g640(.A1(new_n239), .A2(new_n247), .A3(new_n246), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT119), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n843), .B1(new_n244), .B2(new_n245), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n234), .B1(KEYINPUT94), .B2(new_n240), .ZN(new_n845));
  INV_X1    g644(.A(new_n245), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n845), .A2(KEYINPUT119), .A3(new_n846), .A4(new_n243), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n236), .A2(new_n238), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n844), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  AOI22_X1  g648(.A1(new_n842), .A2(new_n253), .B1(new_n849), .B2(new_n252), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n641), .A2(new_n850), .A3(new_n644), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n641), .A2(new_n850), .A3(KEYINPUT120), .A4(new_n644), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT118), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n637), .A2(new_n636), .A3(new_n625), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n631), .A2(KEYINPUT54), .A3(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n578), .B1(new_n638), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n858), .A2(new_n860), .A3(KEYINPUT55), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n642), .ZN(new_n862));
  AOI21_X1  g661(.A(KEYINPUT55), .B1(new_n858), .B2(new_n860), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n856), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n858), .A2(new_n860), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT55), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n867), .A2(KEYINPUT118), .A3(new_n642), .A4(new_n861), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n864), .A2(new_n256), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n734), .B1(new_n855), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n850), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n732), .A2(new_n871), .A3(new_n733), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n864), .A3(new_n868), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n689), .B1(new_n870), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n670), .A2(new_n690), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n692), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n670), .A2(new_n690), .A3(KEYINPUT101), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n877), .A2(new_n257), .A3(new_n645), .A4(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n532), .A2(new_n711), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n698), .A2(new_n560), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n882), .A2(new_n256), .A3(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT121), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n884), .A2(new_n885), .A3(G113gat), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n885), .B1(new_n884), .B2(G113gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n880), .A2(new_n519), .A3(new_n727), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n560), .B1(new_n888), .B2(KEYINPUT122), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n880), .A2(new_n890), .A3(new_n519), .A4(new_n727), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n256), .A2(new_n354), .ZN(new_n893));
  OAI22_X1  g692(.A1(new_n886), .A2(new_n887), .B1(new_n892), .B2(new_n893), .ZN(G1340gat));
  NAND2_X1  g693(.A1(new_n882), .A2(new_n883), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n895), .A2(new_n355), .A3(new_n645), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n889), .A2(new_n646), .A3(new_n891), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n896), .B1(new_n355), .B2(new_n897), .ZN(G1341gat));
  OAI21_X1  g697(.A(G127gat), .B1(new_n895), .B2(new_n689), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n690), .A2(new_n360), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n892), .B2(new_n900), .ZN(G1342gat));
  NOR2_X1   g700(.A1(new_n670), .A2(G134gat), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(KEYINPUT56), .B1(new_n892), .B2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT56), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n889), .A2(new_n905), .A3(new_n891), .A4(new_n902), .ZN(new_n906));
  OAI21_X1  g705(.A(G134gat), .B1(new_n895), .B2(new_n670), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n904), .A2(new_n906), .A3(new_n907), .ZN(G1343gat));
  INV_X1    g707(.A(G141gat), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n572), .A2(new_n532), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n701), .B1(new_n910), .B2(KEYINPUT123), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n911), .B1(KEYINPUT123), .B2(new_n910), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n912), .A2(new_n880), .A3(new_n519), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n909), .B1(new_n913), .B2(new_n257), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT57), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n482), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n867), .A2(new_n642), .A3(new_n861), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n851), .B1(new_n917), .B2(new_n257), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n670), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n690), .B1(new_n919), .B2(new_n873), .ZN(new_n920));
  INV_X1    g719(.A(new_n879), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n916), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n482), .B1(new_n875), .B2(new_n879), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n923), .B2(KEYINPUT57), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n757), .A2(new_n698), .A3(new_n560), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n256), .A2(G141gat), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n914), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT58), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI211_X1 g729(.A(KEYINPUT58), .B(new_n914), .C1(new_n926), .C2(new_n927), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(G1344gat));
  INV_X1    g731(.A(G148gat), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n933), .A2(KEYINPUT59), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n934), .B1(new_n926), .B2(new_n645), .ZN(new_n935));
  INV_X1    g734(.A(new_n916), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n936), .B1(new_n875), .B2(new_n879), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n879), .A2(KEYINPUT124), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n691), .A2(new_n693), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT124), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n939), .A2(new_n940), .A3(new_n257), .A4(new_n645), .ZN(new_n941));
  INV_X1    g740(.A(new_n917), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n871), .A2(new_n670), .ZN(new_n943));
  AOI22_X1  g742(.A1(new_n918), .A2(new_n670), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n938), .B(new_n941), .C1(new_n944), .C2(new_n690), .ZN(new_n945));
  AOI21_X1  g744(.A(KEYINPUT57), .B1(new_n945), .B2(new_n532), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n937), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n925), .A2(new_n646), .ZN(new_n948));
  OAI21_X1  g747(.A(G148gat), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(KEYINPUT59), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(new_n913), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n952), .A2(new_n933), .A3(new_n646), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n953), .ZN(G1345gat));
  OAI21_X1  g753(.A(G155gat), .B1(new_n926), .B2(new_n689), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n952), .A2(new_n368), .A3(new_n690), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(G1346gat));
  INV_X1    g756(.A(new_n734), .ZN(new_n958));
  OAI21_X1  g757(.A(KEYINPUT125), .B1(new_n926), .B2(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT125), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n924), .A2(new_n960), .A3(new_n734), .A4(new_n925), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n959), .A2(G162gat), .A3(new_n961), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n952), .A2(new_n369), .A3(new_n722), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(G1347gat));
  NOR2_X1   g763(.A1(new_n519), .A2(new_n701), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n966), .A2(new_n532), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n880), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n968), .A2(new_n726), .ZN(new_n969));
  AOI21_X1  g768(.A(G169gat), .B1(new_n969), .B2(new_n256), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n880), .A2(new_n881), .A3(new_n965), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n257), .A2(new_n284), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(G1348gat));
  AOI21_X1  g772(.A(G176gat), .B1(new_n969), .B2(new_n646), .ZN(new_n974));
  INV_X1    g773(.A(new_n968), .ZN(new_n975));
  NOR3_X1   g774(.A1(new_n711), .A2(new_n285), .A3(new_n645), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(G1349gat));
  NAND3_X1  g776(.A1(new_n969), .A2(new_n314), .A3(new_n690), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n880), .A2(new_n690), .A3(new_n881), .A4(new_n965), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(G183gat), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(KEYINPUT60), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT60), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n978), .A2(new_n983), .A3(new_n980), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n982), .A2(new_n984), .ZN(G1350gat));
  NAND3_X1  g784(.A1(new_n969), .A2(new_n292), .A3(new_n734), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT61), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n722), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n987), .B1(new_n988), .B2(G190gat), .ZN(new_n989));
  AOI211_X1 g788(.A(KEYINPUT61), .B(new_n292), .C1(new_n971), .C2(new_n722), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n986), .B1(new_n989), .B2(new_n990), .ZN(G1351gat));
  NOR2_X1   g790(.A1(new_n966), .A2(new_n757), .ZN(new_n992));
  AND2_X1   g791(.A1(new_n923), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g792(.A(G197gat), .B1(new_n993), .B2(new_n256), .ZN(new_n994));
  XNOR2_X1  g793(.A(new_n992), .B(KEYINPUT126), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n947), .A2(new_n995), .ZN(new_n996));
  AND2_X1   g795(.A1(new_n256), .A2(G197gat), .ZN(new_n997));
  AOI21_X1  g796(.A(new_n994), .B1(new_n996), .B2(new_n997), .ZN(G1352gat));
  INV_X1    g797(.A(G204gat), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n993), .A2(new_n999), .A3(new_n646), .ZN(new_n1000));
  OR2_X1    g799(.A1(new_n1000), .A2(KEYINPUT62), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1000), .A2(KEYINPUT62), .ZN(new_n1002));
  NOR3_X1   g801(.A1(new_n947), .A2(new_n645), .A3(new_n995), .ZN(new_n1003));
  OAI211_X1 g802(.A(new_n1001), .B(new_n1002), .C1(new_n999), .C2(new_n1003), .ZN(G1353gat));
  NAND2_X1  g803(.A1(new_n992), .A2(new_n690), .ZN(new_n1005));
  INV_X1    g804(.A(new_n1005), .ZN(new_n1006));
  NAND3_X1  g805(.A1(new_n923), .A2(new_n260), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g806(.A(KEYINPUT127), .ZN(new_n1008));
  OAI211_X1 g807(.A(new_n1008), .B(new_n1006), .C1(new_n937), .C2(new_n946), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1009), .A2(G211gat), .ZN(new_n1010));
  AND3_X1   g809(.A1(new_n864), .A2(new_n256), .A3(new_n868), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n853), .A2(new_n854), .ZN(new_n1012));
  OAI21_X1  g811(.A(new_n958), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g812(.A(new_n690), .B1(new_n1013), .B2(new_n873), .ZN(new_n1014));
  OAI21_X1  g813(.A(new_n916), .B1(new_n1014), .B2(new_n921), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n942), .A2(new_n943), .ZN(new_n1016));
  AOI21_X1  g815(.A(new_n690), .B1(new_n919), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n938), .A2(new_n941), .ZN(new_n1018));
  OAI21_X1  g817(.A(new_n532), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1019), .A2(new_n915), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1015), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g820(.A(new_n1008), .B1(new_n1021), .B2(new_n1006), .ZN(new_n1022));
  INV_X1    g821(.A(KEYINPUT63), .ZN(new_n1023));
  NOR3_X1   g822(.A1(new_n1010), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g823(.A(new_n1005), .B1(new_n1015), .B2(new_n1020), .ZN(new_n1025));
  AOI21_X1  g824(.A(new_n260), .B1(new_n1025), .B2(new_n1008), .ZN(new_n1026));
  OAI21_X1  g825(.A(KEYINPUT127), .B1(new_n947), .B2(new_n1005), .ZN(new_n1027));
  AOI21_X1  g826(.A(KEYINPUT63), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g827(.A(new_n1007), .B1(new_n1024), .B2(new_n1028), .ZN(G1354gat));
  NAND3_X1  g828(.A1(new_n993), .A2(new_n261), .A3(new_n734), .ZN(new_n1030));
  NOR3_X1   g829(.A1(new_n947), .A2(new_n670), .A3(new_n995), .ZN(new_n1031));
  OAI21_X1  g830(.A(new_n1030), .B1(new_n1031), .B2(new_n261), .ZN(G1355gat));
endmodule


