

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X2 U323 ( .A(n481), .B(KEYINPUT38), .ZN(n502) );
  XOR2_X2 U324 ( .A(n318), .B(n317), .Z(n558) );
  XNOR2_X1 U325 ( .A(n353), .B(n352), .ZN(n505) );
  XNOR2_X1 U326 ( .A(KEYINPUT37), .B(KEYINPUT103), .ZN(n479) );
  XOR2_X1 U327 ( .A(n446), .B(n445), .Z(n291) );
  XOR2_X1 U328 ( .A(KEYINPUT97), .B(n466), .Z(n292) );
  XOR2_X1 U329 ( .A(n475), .B(KEYINPUT101), .Z(n293) );
  XNOR2_X1 U330 ( .A(KEYINPUT114), .B(KEYINPUT46), .ZN(n368) );
  XNOR2_X1 U331 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U332 ( .A(n394), .B(n393), .ZN(n395) );
  INV_X1 U333 ( .A(KEYINPUT18), .ZN(n407) );
  XNOR2_X1 U334 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U335 ( .A(n420), .B(n351), .ZN(n352) );
  XNOR2_X1 U336 ( .A(n410), .B(n409), .ZN(n443) );
  XNOR2_X1 U337 ( .A(n436), .B(KEYINPUT55), .ZN(n437) );
  XNOR2_X1 U338 ( .A(KEYINPUT26), .B(n464), .ZN(n570) );
  XOR2_X1 U339 ( .A(n451), .B(n450), .Z(n463) );
  XNOR2_X1 U340 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U341 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U342 ( .A(n485), .B(n484), .ZN(G1330GAT) );
  XOR2_X1 U343 ( .A(KEYINPUT74), .B(KEYINPUT73), .Z(n295) );
  XNOR2_X1 U344 ( .A(G43GAT), .B(G92GAT), .ZN(n294) );
  XNOR2_X1 U345 ( .A(n295), .B(n294), .ZN(n318) );
  XOR2_X1 U346 ( .A(KEYINPUT10), .B(KEYINPUT75), .Z(n297) );
  XNOR2_X1 U347 ( .A(G36GAT), .B(G134GAT), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U349 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n299) );
  XNOR2_X1 U350 ( .A(G99GAT), .B(G162GAT), .ZN(n298) );
  XNOR2_X1 U351 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U352 ( .A(n301), .B(n300), .Z(n312) );
  INV_X1 U353 ( .A(G50GAT), .ZN(n302) );
  NAND2_X1 U354 ( .A1(G29GAT), .A2(n302), .ZN(n305) );
  INV_X1 U355 ( .A(G29GAT), .ZN(n303) );
  NAND2_X1 U356 ( .A1(n303), .A2(G50GAT), .ZN(n304) );
  NAND2_X1 U357 ( .A1(n305), .A2(n304), .ZN(n307) );
  XNOR2_X1 U358 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n306) );
  XNOR2_X1 U359 ( .A(n307), .B(n306), .ZN(n342) );
  XOR2_X1 U360 ( .A(KEYINPUT76), .B(G218GAT), .Z(n309) );
  NAND2_X1 U361 ( .A1(G232GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U362 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n342), .B(n310), .ZN(n311) );
  XNOR2_X1 U364 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U365 ( .A(n313), .B(KEYINPUT65), .Z(n316) );
  XNOR2_X1 U366 ( .A(G106GAT), .B(G85GAT), .ZN(n314) );
  XNOR2_X1 U367 ( .A(n314), .B(KEYINPUT72), .ZN(n358) );
  XNOR2_X1 U368 ( .A(G190GAT), .B(n358), .ZN(n315) );
  XNOR2_X1 U369 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U370 ( .A(KEYINPUT1), .B(KEYINPUT92), .Z(n320) );
  XNOR2_X1 U371 ( .A(G57GAT), .B(KEYINPUT6), .ZN(n319) );
  XNOR2_X1 U372 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U373 ( .A(KEYINPUT4), .B(n321), .Z(n323) );
  NAND2_X1 U374 ( .A1(G225GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U375 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U376 ( .A(n324), .B(KEYINPUT93), .Z(n329) );
  XOR2_X1 U377 ( .A(KEYINPUT2), .B(G162GAT), .Z(n326) );
  XNOR2_X1 U378 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n325) );
  XNOR2_X1 U379 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U380 ( .A(KEYINPUT89), .B(n327), .Z(n435) );
  XNOR2_X1 U381 ( .A(G1GAT), .B(n435), .ZN(n328) );
  XNOR2_X1 U382 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U383 ( .A(KEYINPUT75), .B(G85GAT), .Z(n331) );
  XNOR2_X1 U384 ( .A(G141GAT), .B(G29GAT), .ZN(n330) );
  XNOR2_X1 U385 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U386 ( .A(n333), .B(n332), .Z(n341) );
  XOR2_X1 U387 ( .A(KEYINPUT81), .B(G134GAT), .Z(n335) );
  XNOR2_X1 U388 ( .A(KEYINPUT80), .B(G127GAT), .ZN(n334) );
  XNOR2_X1 U389 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U390 ( .A(KEYINPUT0), .B(n336), .Z(n445) );
  XOR2_X1 U391 ( .A(KEYINPUT5), .B(G148GAT), .Z(n338) );
  XNOR2_X1 U392 ( .A(G113GAT), .B(G120GAT), .ZN(n337) );
  XNOR2_X1 U393 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U394 ( .A(n445), .B(n339), .ZN(n340) );
  XNOR2_X1 U395 ( .A(n341), .B(n340), .ZN(n519) );
  INV_X1 U396 ( .A(n558), .ZN(n486) );
  XNOR2_X1 U397 ( .A(n342), .B(KEYINPUT30), .ZN(n343) );
  XNOR2_X1 U398 ( .A(n343), .B(KEYINPUT68), .ZN(n346) );
  XOR2_X1 U399 ( .A(G1GAT), .B(KEYINPUT67), .Z(n385) );
  XNOR2_X1 U400 ( .A(G169GAT), .B(n385), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n344), .B(KEYINPUT29), .ZN(n345) );
  XNOR2_X1 U402 ( .A(n346), .B(n345), .ZN(n350) );
  XNOR2_X1 U403 ( .A(G43GAT), .B(G15GAT), .ZN(n347) );
  XNOR2_X1 U404 ( .A(n347), .B(G113GAT), .ZN(n444) );
  XNOR2_X1 U405 ( .A(G36GAT), .B(G197GAT), .ZN(n348) );
  XNOR2_X1 U406 ( .A(n348), .B(G8GAT), .ZN(n411) );
  XOR2_X1 U407 ( .A(n444), .B(n411), .Z(n349) );
  XNOR2_X1 U408 ( .A(n350), .B(n349), .ZN(n353) );
  XOR2_X1 U409 ( .A(G141GAT), .B(G22GAT), .Z(n420) );
  NAND2_X1 U410 ( .A1(G229GAT), .A2(G233GAT), .ZN(n351) );
  INV_X1 U411 ( .A(n505), .ZN(n547) );
  XNOR2_X1 U412 ( .A(G57GAT), .B(KEYINPUT70), .ZN(n354) );
  XNOR2_X1 U413 ( .A(n354), .B(KEYINPUT13), .ZN(n386) );
  XOR2_X1 U414 ( .A(G64GAT), .B(G92GAT), .Z(n356) );
  XNOR2_X1 U415 ( .A(G176GAT), .B(G204GAT), .ZN(n355) );
  XNOR2_X1 U416 ( .A(n356), .B(n355), .ZN(n404) );
  XOR2_X1 U417 ( .A(n386), .B(n404), .Z(n360) );
  XNOR2_X1 U418 ( .A(G99GAT), .B(G71GAT), .ZN(n357) );
  XNOR2_X1 U419 ( .A(n357), .B(G120GAT), .ZN(n446) );
  XNOR2_X1 U420 ( .A(n446), .B(n358), .ZN(n359) );
  XNOR2_X1 U421 ( .A(n360), .B(n359), .ZN(n367) );
  XOR2_X1 U422 ( .A(G148GAT), .B(G78GAT), .Z(n429) );
  XOR2_X1 U423 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n362) );
  XNOR2_X1 U424 ( .A(KEYINPUT71), .B(KEYINPUT31), .ZN(n361) );
  XNOR2_X1 U425 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U426 ( .A(n429), .B(n363), .Z(n365) );
  NAND2_X1 U427 ( .A1(G230GAT), .A2(G233GAT), .ZN(n364) );
  XOR2_X1 U428 ( .A(n365), .B(n364), .Z(n366) );
  XNOR2_X1 U429 ( .A(n367), .B(n366), .ZN(n575) );
  XOR2_X1 U430 ( .A(KEYINPUT41), .B(n575), .Z(n553) );
  NOR2_X1 U431 ( .A1(n547), .A2(n553), .ZN(n369) );
  NOR2_X1 U432 ( .A1(n486), .A2(n370), .ZN(n391) );
  XOR2_X1 U433 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n372) );
  XNOR2_X1 U434 ( .A(G8GAT), .B(G64GAT), .ZN(n371) );
  XNOR2_X1 U435 ( .A(n372), .B(n371), .ZN(n384) );
  XOR2_X1 U436 ( .A(G78GAT), .B(G211GAT), .Z(n374) );
  XNOR2_X1 U437 ( .A(G22GAT), .B(G155GAT), .ZN(n373) );
  XNOR2_X1 U438 ( .A(n374), .B(n373), .ZN(n382) );
  XOR2_X1 U439 ( .A(KEYINPUT79), .B(KEYINPUT78), .Z(n376) );
  XNOR2_X1 U440 ( .A(KEYINPUT15), .B(KEYINPUT77), .ZN(n375) );
  XNOR2_X1 U441 ( .A(n376), .B(n375), .ZN(n380) );
  XOR2_X1 U442 ( .A(G71GAT), .B(G127GAT), .Z(n378) );
  XNOR2_X1 U443 ( .A(G15GAT), .B(G183GAT), .ZN(n377) );
  XNOR2_X1 U444 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U445 ( .A(n380), .B(n379), .Z(n381) );
  XNOR2_X1 U446 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U447 ( .A(n384), .B(n383), .ZN(n390) );
  XOR2_X1 U448 ( .A(n386), .B(n385), .Z(n388) );
  NAND2_X1 U449 ( .A1(G231GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U450 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U451 ( .A(n390), .B(n389), .Z(n477) );
  INV_X1 U452 ( .A(n477), .ZN(n579) );
  NAND2_X1 U453 ( .A1(n391), .A2(n579), .ZN(n392) );
  XNOR2_X1 U454 ( .A(n392), .B(KEYINPUT47), .ZN(n398) );
  XOR2_X1 U455 ( .A(n505), .B(KEYINPUT69), .Z(n531) );
  XOR2_X1 U456 ( .A(KEYINPUT36), .B(n558), .Z(n581) );
  NAND2_X1 U457 ( .A1(n477), .A2(n581), .ZN(n394) );
  XOR2_X1 U458 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n393) );
  NAND2_X1 U459 ( .A1(n395), .A2(n575), .ZN(n396) );
  NOR2_X1 U460 ( .A1(n531), .A2(n396), .ZN(n397) );
  NOR2_X1 U461 ( .A1(n398), .A2(n397), .ZN(n399) );
  XNOR2_X1 U462 ( .A(n399), .B(KEYINPUT48), .ZN(n532) );
  XOR2_X1 U463 ( .A(G211GAT), .B(KEYINPUT88), .Z(n401) );
  XNOR2_X1 U464 ( .A(G218GAT), .B(KEYINPUT21), .ZN(n400) );
  XNOR2_X1 U465 ( .A(n401), .B(n400), .ZN(n421) );
  XOR2_X1 U466 ( .A(KEYINPUT94), .B(n421), .Z(n403) );
  NAND2_X1 U467 ( .A1(G226GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U468 ( .A(n403), .B(n402), .ZN(n405) );
  XOR2_X1 U469 ( .A(n405), .B(n404), .Z(n413) );
  XNOR2_X1 U470 ( .A(G183GAT), .B(KEYINPUT19), .ZN(n406) );
  XNOR2_X1 U471 ( .A(n406), .B(KEYINPUT17), .ZN(n410) );
  XNOR2_X1 U472 ( .A(G169GAT), .B(G190GAT), .ZN(n408) );
  XNOR2_X1 U473 ( .A(n411), .B(n443), .ZN(n412) );
  XOR2_X1 U474 ( .A(n413), .B(n412), .Z(n457) );
  BUF_X1 U475 ( .A(n457), .Z(n521) );
  XNOR2_X1 U476 ( .A(KEYINPUT119), .B(n521), .ZN(n414) );
  NOR2_X1 U477 ( .A1(n532), .A2(n414), .ZN(n415) );
  XOR2_X1 U478 ( .A(KEYINPUT54), .B(n415), .Z(n416) );
  NOR2_X1 U479 ( .A1(n519), .A2(n416), .ZN(n417) );
  XOR2_X1 U480 ( .A(KEYINPUT64), .B(n417), .Z(n571) );
  XOR2_X1 U481 ( .A(KEYINPUT23), .B(KEYINPUT90), .Z(n419) );
  XNOR2_X1 U482 ( .A(KEYINPUT22), .B(KEYINPUT87), .ZN(n418) );
  XNOR2_X1 U483 ( .A(n419), .B(n418), .ZN(n425) );
  XOR2_X1 U484 ( .A(n421), .B(n420), .Z(n423) );
  NAND2_X1 U485 ( .A1(G228GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U486 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U487 ( .A(n425), .B(n424), .ZN(n433) );
  XOR2_X1 U488 ( .A(KEYINPUT91), .B(KEYINPUT24), .Z(n427) );
  XNOR2_X1 U489 ( .A(G50GAT), .B(G106GAT), .ZN(n426) );
  XNOR2_X1 U490 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U491 ( .A(n428), .B(G204GAT), .Z(n431) );
  XNOR2_X1 U492 ( .A(G197GAT), .B(n429), .ZN(n430) );
  XNOR2_X1 U493 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U494 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U495 ( .A(n435), .B(n434), .ZN(n468) );
  NOR2_X1 U496 ( .A1(n571), .A2(n468), .ZN(n438) );
  XNOR2_X1 U497 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n436) );
  XNOR2_X1 U498 ( .A(n438), .B(n437), .ZN(n452) );
  XOR2_X1 U499 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n440) );
  XNOR2_X1 U500 ( .A(G176GAT), .B(KEYINPUT83), .ZN(n439) );
  XNOR2_X1 U501 ( .A(n440), .B(n439), .ZN(n442) );
  XOR2_X1 U502 ( .A(KEYINPUT82), .B(KEYINPUT85), .Z(n441) );
  XNOR2_X1 U503 ( .A(n442), .B(n441), .ZN(n449) );
  XNOR2_X1 U504 ( .A(n444), .B(n443), .ZN(n447) );
  XNOR2_X1 U505 ( .A(n447), .B(n291), .ZN(n448) );
  XNOR2_X1 U506 ( .A(n449), .B(n448), .ZN(n451) );
  NAND2_X1 U507 ( .A1(G227GAT), .A2(G233GAT), .ZN(n450) );
  INV_X1 U508 ( .A(n463), .ZN(n535) );
  NAND2_X1 U509 ( .A1(n452), .A2(n535), .ZN(n568) );
  NOR2_X1 U510 ( .A1(n558), .A2(n568), .ZN(n456) );
  XNOR2_X1 U511 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n454) );
  INV_X1 U512 ( .A(G190GAT), .ZN(n453) );
  XNOR2_X1 U513 ( .A(n456), .B(n455), .ZN(G1351GAT) );
  NAND2_X1 U514 ( .A1(n575), .A2(n531), .ZN(n491) );
  XOR2_X1 U515 ( .A(n457), .B(KEYINPUT95), .Z(n458) );
  XOR2_X1 U516 ( .A(n458), .B(KEYINPUT27), .Z(n465) );
  INV_X1 U517 ( .A(n465), .ZN(n459) );
  NAND2_X1 U518 ( .A1(n459), .A2(n519), .ZN(n460) );
  XOR2_X1 U519 ( .A(KEYINPUT96), .B(n460), .Z(n548) );
  XNOR2_X1 U520 ( .A(KEYINPUT28), .B(n468), .ZN(n525) );
  INV_X1 U521 ( .A(n525), .ZN(n461) );
  NAND2_X1 U522 ( .A1(n548), .A2(n461), .ZN(n533) );
  XOR2_X1 U523 ( .A(KEYINPUT86), .B(n463), .Z(n462) );
  NOR2_X1 U524 ( .A1(n533), .A2(n462), .ZN(n476) );
  NAND2_X1 U525 ( .A1(n463), .A2(n468), .ZN(n464) );
  NOR2_X1 U526 ( .A1(n570), .A2(n465), .ZN(n466) );
  AND2_X1 U527 ( .A1(n521), .A2(n535), .ZN(n467) );
  NOR2_X1 U528 ( .A1(n468), .A2(n467), .ZN(n471) );
  XNOR2_X1 U529 ( .A(KEYINPUT25), .B(KEYINPUT99), .ZN(n469) );
  XNOR2_X1 U530 ( .A(n469), .B(KEYINPUT98), .ZN(n470) );
  XNOR2_X1 U531 ( .A(n471), .B(n470), .ZN(n472) );
  NOR2_X1 U532 ( .A1(n292), .A2(n472), .ZN(n473) );
  XNOR2_X1 U533 ( .A(n473), .B(KEYINPUT100), .ZN(n474) );
  NOR2_X1 U534 ( .A1(n519), .A2(n474), .ZN(n475) );
  NOR2_X1 U535 ( .A1(n476), .A2(n293), .ZN(n489) );
  NOR2_X1 U536 ( .A1(n477), .A2(n489), .ZN(n478) );
  NAND2_X1 U537 ( .A1(n581), .A2(n478), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n480), .B(n479), .ZN(n517) );
  NOR2_X1 U539 ( .A1(n491), .A2(n517), .ZN(n481) );
  NAND2_X1 U540 ( .A1(n535), .A2(n502), .ZN(n485) );
  XOR2_X1 U541 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n483) );
  XNOR2_X1 U542 ( .A(G43GAT), .B(KEYINPUT105), .ZN(n482) );
  XNOR2_X1 U543 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n493) );
  NOR2_X1 U544 ( .A1(n486), .A2(n579), .ZN(n487) );
  XOR2_X1 U545 ( .A(KEYINPUT16), .B(n487), .Z(n488) );
  NOR2_X1 U546 ( .A1(n489), .A2(n488), .ZN(n490) );
  XOR2_X1 U547 ( .A(KEYINPUT102), .B(n490), .Z(n507) );
  NOR2_X1 U548 ( .A1(n507), .A2(n491), .ZN(n497) );
  NAND2_X1 U549 ( .A1(n519), .A2(n497), .ZN(n492) );
  XNOR2_X1 U550 ( .A(n493), .B(n492), .ZN(G1324GAT) );
  NAND2_X1 U551 ( .A1(n521), .A2(n497), .ZN(n494) );
  XNOR2_X1 U552 ( .A(n494), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U553 ( .A(G15GAT), .B(KEYINPUT35), .Z(n496) );
  NAND2_X1 U554 ( .A1(n497), .A2(n535), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n496), .B(n495), .ZN(G1326GAT) );
  NAND2_X1 U556 ( .A1(n497), .A2(n525), .ZN(n498) );
  XNOR2_X1 U557 ( .A(n498), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U558 ( .A(G29GAT), .B(KEYINPUT39), .Z(n500) );
  NAND2_X1 U559 ( .A1(n519), .A2(n502), .ZN(n499) );
  XNOR2_X1 U560 ( .A(n500), .B(n499), .ZN(G1328GAT) );
  NAND2_X1 U561 ( .A1(n502), .A2(n521), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n501), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U563 ( .A1(n502), .A2(n525), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n503), .B(KEYINPUT106), .ZN(n504) );
  XNOR2_X1 U565 ( .A(G50GAT), .B(n504), .ZN(G1331GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n509) );
  XOR2_X1 U567 ( .A(n553), .B(KEYINPUT107), .Z(n562) );
  NOR2_X1 U568 ( .A1(n562), .A2(n505), .ZN(n506) );
  XOR2_X1 U569 ( .A(KEYINPUT108), .B(n506), .Z(n518) );
  NOR2_X1 U570 ( .A1(n507), .A2(n518), .ZN(n514) );
  NAND2_X1 U571 ( .A1(n514), .A2(n519), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U573 ( .A(G57GAT), .B(n510), .ZN(G1332GAT) );
  NAND2_X1 U574 ( .A1(n521), .A2(n514), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n511), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U576 ( .A1(n514), .A2(n535), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n512), .B(KEYINPUT110), .ZN(n513) );
  XNOR2_X1 U578 ( .A(G71GAT), .B(n513), .ZN(G1334GAT) );
  XOR2_X1 U579 ( .A(G78GAT), .B(KEYINPUT43), .Z(n516) );
  NAND2_X1 U580 ( .A1(n514), .A2(n525), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  NOR2_X1 U582 ( .A1(n518), .A2(n517), .ZN(n526) );
  NAND2_X1 U583 ( .A1(n519), .A2(n526), .ZN(n520) );
  XNOR2_X1 U584 ( .A(G85GAT), .B(n520), .ZN(G1336GAT) );
  XOR2_X1 U585 ( .A(G92GAT), .B(KEYINPUT111), .Z(n523) );
  NAND2_X1 U586 ( .A1(n526), .A2(n521), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n523), .B(n522), .ZN(G1337GAT) );
  NAND2_X1 U588 ( .A1(n526), .A2(n535), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n524), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U590 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n530) );
  XOR2_X1 U591 ( .A(KEYINPUT113), .B(KEYINPUT112), .Z(n528) );
  NAND2_X1 U592 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n530), .B(n529), .ZN(G1339GAT) );
  INV_X1 U595 ( .A(n531), .ZN(n560) );
  NOR2_X1 U596 ( .A1(n532), .A2(n533), .ZN(n534) );
  NAND2_X1 U597 ( .A1(n535), .A2(n534), .ZN(n542) );
  NOR2_X1 U598 ( .A1(n560), .A2(n542), .ZN(n536) );
  XOR2_X1 U599 ( .A(G113GAT), .B(n536), .Z(G1340GAT) );
  NOR2_X1 U600 ( .A1(n562), .A2(n542), .ZN(n538) );
  XNOR2_X1 U601 ( .A(KEYINPUT115), .B(KEYINPUT49), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U603 ( .A(G120GAT), .B(n539), .Z(G1341GAT) );
  NOR2_X1 U604 ( .A1(n579), .A2(n542), .ZN(n540) );
  XOR2_X1 U605 ( .A(KEYINPUT50), .B(n540), .Z(n541) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n541), .ZN(G1342GAT) );
  NOR2_X1 U607 ( .A1(n542), .A2(n558), .ZN(n546) );
  XOR2_X1 U608 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n544) );
  XNOR2_X1 U609 ( .A(G134GAT), .B(KEYINPUT117), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n546), .B(n545), .ZN(G1343GAT) );
  NOR2_X1 U612 ( .A1(n570), .A2(n532), .ZN(n549) );
  NAND2_X1 U613 ( .A1(n549), .A2(n548), .ZN(n557) );
  NOR2_X1 U614 ( .A1(n547), .A2(n557), .ZN(n550) );
  XOR2_X1 U615 ( .A(G141GAT), .B(n550), .Z(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT52), .B(KEYINPUT53), .Z(n552) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(n555) );
  NOR2_X1 U619 ( .A1(n553), .A2(n557), .ZN(n554) );
  XOR2_X1 U620 ( .A(n555), .B(n554), .Z(G1345GAT) );
  NOR2_X1 U621 ( .A1(n579), .A2(n557), .ZN(n556) );
  XOR2_X1 U622 ( .A(G155GAT), .B(n556), .Z(G1346GAT) );
  NOR2_X1 U623 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U624 ( .A(G162GAT), .B(n559), .Z(G1347GAT) );
  NOR2_X1 U625 ( .A1(n560), .A2(n568), .ZN(n561) );
  XOR2_X1 U626 ( .A(G169GAT), .B(n561), .Z(G1348GAT) );
  NOR2_X1 U627 ( .A1(n562), .A2(n568), .ZN(n567) );
  XOR2_X1 U628 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n564) );
  XNOR2_X1 U629 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(KEYINPUT56), .B(n565), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(G1349GAT) );
  NOR2_X1 U633 ( .A1(n579), .A2(n568), .ZN(n569) );
  XOR2_X1 U634 ( .A(G183GAT), .B(n569), .Z(G1350GAT) );
  NOR2_X1 U635 ( .A1(n571), .A2(n570), .ZN(n582) );
  INV_X1 U636 ( .A(n582), .ZN(n578) );
  NOR2_X1 U637 ( .A1(n547), .A2(n578), .ZN(n573) );
  XNOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(n574), .ZN(G1352GAT) );
  NOR2_X1 U641 ( .A1(n575), .A2(n578), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U645 ( .A(G211GAT), .B(n580), .Z(G1354GAT) );
  NAND2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(n583), .B(KEYINPUT62), .ZN(n584) );
  XOR2_X1 U648 ( .A(n584), .B(KEYINPUT125), .Z(n586) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(G1355GAT) );
endmodule

