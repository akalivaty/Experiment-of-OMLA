

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U547 ( .A1(n537), .A2(n533), .ZN(n532) );
  NOR2_X1 U548 ( .A1(n715), .A2(n714), .ZN(n717) );
  AND2_X1 U549 ( .A1(n555), .A2(n554), .ZN(G164) );
  XNOR2_X1 U550 ( .A(n539), .B(KEYINPUT64), .ZN(n787) );
  OR2_X1 U551 ( .A1(G164), .A2(G1384), .ZN(n539) );
  AND2_X1 U552 ( .A1(n765), .A2(n540), .ZN(n755) );
  AND2_X1 U553 ( .A1(n544), .A2(n543), .ZN(n804) );
  NAND2_X1 U554 ( .A1(n525), .A2(n522), .ZN(n521) );
  NAND2_X1 U555 ( .A1(n835), .A2(n523), .ZN(n522) );
  NAND2_X1 U556 ( .A1(n527), .A2(n526), .ZN(n525) );
  NAND2_X1 U557 ( .A1(n524), .A2(n526), .ZN(n523) );
  XNOR2_X1 U558 ( .A(KEYINPUT30), .B(KEYINPUT100), .ZN(n708) );
  AND2_X1 U559 ( .A1(G286), .A2(KEYINPUT102), .ZN(n538) );
  NAND2_X1 U560 ( .A1(n535), .A2(n534), .ZN(n533) );
  NAND2_X1 U561 ( .A1(n749), .A2(n536), .ZN(n535) );
  OR2_X1 U562 ( .A1(n749), .A2(KEYINPUT102), .ZN(n534) );
  OR2_X1 U563 ( .A1(G286), .A2(KEYINPUT102), .ZN(n536) );
  AND2_X1 U564 ( .A1(n749), .A2(n530), .ZN(n529) );
  INV_X1 U565 ( .A(KEYINPUT102), .ZN(n530) );
  NAND2_X1 U566 ( .A1(n730), .A2(G8), .ZN(n703) );
  INV_X1 U567 ( .A(n821), .ZN(n524) );
  INV_X1 U568 ( .A(n835), .ZN(n527) );
  INV_X1 U569 ( .A(KEYINPUT40), .ZN(n526) );
  NAND2_X1 U570 ( .A1(n551), .A2(n542), .ZN(n541) );
  INV_X1 U571 ( .A(G2105), .ZN(n542) );
  INV_X1 U572 ( .A(n820), .ZN(n517) );
  OR2_X1 U573 ( .A1(n787), .A2(n786), .ZN(n730) );
  INV_X1 U574 ( .A(n730), .ZN(n720) );
  XNOR2_X1 U575 ( .A(n703), .B(KEYINPUT95), .ZN(n765) );
  NAND2_X1 U576 ( .A1(n821), .A2(KEYINPUT40), .ZN(n510) );
  AND2_X1 U577 ( .A1(n835), .A2(n526), .ZN(n511) );
  NAND2_X1 U578 ( .A1(n518), .A2(n512), .ZN(G329) );
  NAND2_X1 U579 ( .A1(n515), .A2(n513), .ZN(n512) );
  NAND2_X1 U580 ( .A1(n820), .A2(n514), .ZN(n513) );
  NAND2_X1 U581 ( .A1(n819), .A2(n511), .ZN(n514) );
  NAND2_X1 U582 ( .A1(n517), .A2(n516), .ZN(n515) );
  INV_X1 U583 ( .A(n520), .ZN(n516) );
  NAND2_X1 U584 ( .A1(n519), .A2(n520), .ZN(n518) );
  NAND2_X1 U585 ( .A1(n521), .A2(n510), .ZN(n520) );
  NAND2_X1 U586 ( .A1(n819), .A2(n521), .ZN(n519) );
  NAND2_X1 U587 ( .A1(n532), .A2(n528), .ZN(n750) );
  NAND2_X1 U588 ( .A1(n531), .A2(n529), .ZN(n528) );
  INV_X1 U589 ( .A(n756), .ZN(n531) );
  NAND2_X1 U590 ( .A1(n756), .A2(n538), .ZN(n537) );
  NAND2_X1 U591 ( .A1(n748), .A2(n747), .ZN(n756) );
  NOR2_X1 U592 ( .A1(n755), .A2(n752), .ZN(n707) );
  INV_X1 U593 ( .A(G1966), .ZN(n540) );
  NAND2_X1 U594 ( .A1(n884), .A2(G138), .ZN(n549) );
  XNOR2_X2 U595 ( .A(n541), .B(KEYINPUT17), .ZN(n884) );
  INV_X1 U596 ( .A(n982), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n546), .A2(n545), .ZN(n544) );
  INV_X1 U598 ( .A(KEYINPUT33), .ZN(n545) );
  NAND2_X1 U599 ( .A1(n547), .A2(n764), .ZN(n546) );
  XNOR2_X1 U600 ( .A(n763), .B(KEYINPUT104), .ZN(n547) );
  INV_X1 U601 ( .A(KEYINPUT31), .ZN(n716) );
  NOR2_X1 U602 ( .A1(G651), .A2(n660), .ZN(n666) );
  INV_X1 U603 ( .A(G2104), .ZN(n551) );
  NOR2_X2 U604 ( .A1(G2105), .A2(n551), .ZN(n886) );
  NAND2_X1 U605 ( .A1(G102), .A2(n886), .ZN(n548) );
  NAND2_X1 U606 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U607 ( .A(n550), .B(KEYINPUT87), .ZN(n555) );
  AND2_X1 U608 ( .A1(n551), .A2(G2105), .ZN(n880) );
  NAND2_X1 U609 ( .A1(G126), .A2(n880), .ZN(n553) );
  AND2_X1 U610 ( .A1(G2104), .A2(G2105), .ZN(n881) );
  NAND2_X1 U611 ( .A1(G114), .A2(n881), .ZN(n552) );
  AND2_X1 U612 ( .A1(n553), .A2(n552), .ZN(n554) );
  NAND2_X1 U613 ( .A1(G101), .A2(n886), .ZN(n556) );
  XOR2_X1 U614 ( .A(KEYINPUT23), .B(n556), .Z(n559) );
  NAND2_X1 U615 ( .A1(G125), .A2(n880), .ZN(n557) );
  XOR2_X1 U616 ( .A(KEYINPUT65), .B(n557), .Z(n558) );
  NAND2_X1 U617 ( .A1(n559), .A2(n558), .ZN(n563) );
  NAND2_X1 U618 ( .A1(n881), .A2(G113), .ZN(n561) );
  NAND2_X1 U619 ( .A1(n884), .A2(G137), .ZN(n560) );
  NAND2_X1 U620 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U621 ( .A1(n563), .A2(n562), .ZN(G160) );
  XOR2_X1 U622 ( .A(G543), .B(KEYINPUT0), .Z(n660) );
  NAND2_X1 U623 ( .A1(G52), .A2(n666), .ZN(n566) );
  XOR2_X1 U624 ( .A(KEYINPUT66), .B(G651), .Z(n567) );
  NOR2_X1 U625 ( .A1(G543), .A2(n567), .ZN(n564) );
  XOR2_X1 U626 ( .A(KEYINPUT1), .B(n564), .Z(n675) );
  NAND2_X1 U627 ( .A1(G64), .A2(n675), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n566), .A2(n565), .ZN(n575) );
  NOR2_X1 U629 ( .A1(n660), .A2(n567), .ZN(n670) );
  NAND2_X1 U630 ( .A1(G77), .A2(n670), .ZN(n568) );
  XNOR2_X1 U631 ( .A(KEYINPUT69), .B(n568), .ZN(n571) );
  NOR2_X1 U632 ( .A1(G543), .A2(G651), .ZN(n667) );
  NAND2_X1 U633 ( .A1(n667), .A2(G90), .ZN(n569) );
  XOR2_X1 U634 ( .A(n569), .B(KEYINPUT68), .Z(n570) );
  NOR2_X1 U635 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U636 ( .A(KEYINPUT70), .B(n572), .Z(n573) );
  XOR2_X1 U637 ( .A(KEYINPUT9), .B(n573), .Z(n574) );
  NOR2_X1 U638 ( .A1(n575), .A2(n574), .ZN(G171) );
  NAND2_X1 U639 ( .A1(G78), .A2(n670), .ZN(n583) );
  NAND2_X1 U640 ( .A1(G53), .A2(n666), .ZN(n577) );
  NAND2_X1 U641 ( .A1(G65), .A2(n675), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(KEYINPUT72), .B(n578), .ZN(n581) );
  NAND2_X1 U644 ( .A1(G91), .A2(n667), .ZN(n579) );
  XNOR2_X1 U645 ( .A(KEYINPUT71), .B(n579), .ZN(n580) );
  NOR2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(KEYINPUT73), .B(n584), .ZN(n725) );
  INV_X1 U649 ( .A(n725), .ZN(G299) );
  AND2_X1 U650 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U651 ( .A(G57), .ZN(G237) );
  INV_X1 U652 ( .A(G132), .ZN(G219) );
  NAND2_X1 U653 ( .A1(G50), .A2(n666), .ZN(n586) );
  NAND2_X1 U654 ( .A1(G62), .A2(n675), .ZN(n585) );
  NAND2_X1 U655 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U656 ( .A(KEYINPUT84), .B(n587), .Z(n591) );
  NAND2_X1 U657 ( .A1(n670), .A2(G75), .ZN(n589) );
  NAND2_X1 U658 ( .A1(n667), .A2(G88), .ZN(n588) );
  AND2_X1 U659 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U660 ( .A1(n591), .A2(n590), .ZN(G303) );
  NAND2_X1 U661 ( .A1(G7), .A2(G661), .ZN(n592) );
  XOR2_X1 U662 ( .A(n592), .B(KEYINPUT10), .Z(n836) );
  NAND2_X1 U663 ( .A1(n836), .A2(G567), .ZN(n593) );
  XOR2_X1 U664 ( .A(KEYINPUT11), .B(n593), .Z(G234) );
  NAND2_X1 U665 ( .A1(n675), .A2(G56), .ZN(n594) );
  XNOR2_X1 U666 ( .A(n594), .B(KEYINPUT14), .ZN(n595) );
  XNOR2_X1 U667 ( .A(KEYINPUT75), .B(n595), .ZN(n602) );
  NAND2_X1 U668 ( .A1(n667), .A2(G81), .ZN(n596) );
  XOR2_X1 U669 ( .A(KEYINPUT12), .B(n596), .Z(n599) );
  NAND2_X1 U670 ( .A1(G68), .A2(n670), .ZN(n597) );
  XOR2_X1 U671 ( .A(KEYINPUT76), .B(n597), .Z(n598) );
  NOR2_X1 U672 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U673 ( .A(KEYINPUT13), .B(n600), .ZN(n601) );
  NOR2_X1 U674 ( .A1(n602), .A2(n601), .ZN(n604) );
  NAND2_X1 U675 ( .A1(n666), .A2(G43), .ZN(n603) );
  NAND2_X1 U676 ( .A1(n604), .A2(n603), .ZN(n997) );
  INV_X1 U677 ( .A(G860), .ZN(n644) );
  OR2_X1 U678 ( .A1(n997), .A2(n644), .ZN(G153) );
  XNOR2_X1 U679 ( .A(G171), .B(KEYINPUT77), .ZN(G301) );
  NAND2_X1 U680 ( .A1(G868), .A2(G301), .ZN(n605) );
  XNOR2_X1 U681 ( .A(n605), .B(KEYINPUT78), .ZN(n615) );
  NAND2_X1 U682 ( .A1(G66), .A2(n675), .ZN(n612) );
  NAND2_X1 U683 ( .A1(G54), .A2(n666), .ZN(n607) );
  NAND2_X1 U684 ( .A1(G92), .A2(n667), .ZN(n606) );
  NAND2_X1 U685 ( .A1(n607), .A2(n606), .ZN(n610) );
  NAND2_X1 U686 ( .A1(G79), .A2(n670), .ZN(n608) );
  XNOR2_X1 U687 ( .A(KEYINPUT79), .B(n608), .ZN(n609) );
  NOR2_X1 U688 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U689 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U690 ( .A(KEYINPUT15), .B(n613), .ZN(n990) );
  OR2_X1 U691 ( .A1(G868), .A2(n990), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(G284) );
  NAND2_X1 U693 ( .A1(n667), .A2(G89), .ZN(n616) );
  XNOR2_X1 U694 ( .A(n616), .B(KEYINPUT4), .ZN(n618) );
  NAND2_X1 U695 ( .A1(G76), .A2(n670), .ZN(n617) );
  NAND2_X1 U696 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U697 ( .A(n619), .B(KEYINPUT5), .ZN(n624) );
  NAND2_X1 U698 ( .A1(G51), .A2(n666), .ZN(n621) );
  NAND2_X1 U699 ( .A1(G63), .A2(n675), .ZN(n620) );
  NAND2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X1 U701 ( .A(KEYINPUT6), .B(n622), .Z(n623) );
  NAND2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U703 ( .A(n625), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U704 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U705 ( .A(KEYINPUT80), .B(G868), .Z(n626) );
  NOR2_X1 U706 ( .A1(G286), .A2(n626), .ZN(n628) );
  NOR2_X1 U707 ( .A1(G868), .A2(G299), .ZN(n627) );
  NOR2_X1 U708 ( .A1(n628), .A2(n627), .ZN(G297) );
  NAND2_X1 U709 ( .A1(n644), .A2(G559), .ZN(n629) );
  NAND2_X1 U710 ( .A1(n629), .A2(n990), .ZN(n630) );
  XNOR2_X1 U711 ( .A(n630), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U712 ( .A1(G868), .A2(n997), .ZN(n633) );
  NAND2_X1 U713 ( .A1(G868), .A2(n990), .ZN(n631) );
  NOR2_X1 U714 ( .A1(G559), .A2(n631), .ZN(n632) );
  NOR2_X1 U715 ( .A1(n633), .A2(n632), .ZN(G282) );
  XNOR2_X1 U716 ( .A(G2100), .B(KEYINPUT81), .ZN(n642) );
  NAND2_X1 U717 ( .A1(n880), .A2(G123), .ZN(n634) );
  XNOR2_X1 U718 ( .A(n634), .B(KEYINPUT18), .ZN(n636) );
  NAND2_X1 U719 ( .A1(G99), .A2(n886), .ZN(n635) );
  NAND2_X1 U720 ( .A1(n636), .A2(n635), .ZN(n640) );
  NAND2_X1 U721 ( .A1(G135), .A2(n884), .ZN(n638) );
  NAND2_X1 U722 ( .A1(G111), .A2(n881), .ZN(n637) );
  NAND2_X1 U723 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U724 ( .A1(n640), .A2(n639), .ZN(n928) );
  XNOR2_X1 U725 ( .A(n928), .B(G2096), .ZN(n641) );
  NAND2_X1 U726 ( .A1(n642), .A2(n641), .ZN(G156) );
  NAND2_X1 U727 ( .A1(G559), .A2(n990), .ZN(n643) );
  XOR2_X1 U728 ( .A(n997), .B(n643), .Z(n683) );
  NAND2_X1 U729 ( .A1(n644), .A2(n683), .ZN(n652) );
  NAND2_X1 U730 ( .A1(G55), .A2(n666), .ZN(n646) );
  NAND2_X1 U731 ( .A1(G93), .A2(n667), .ZN(n645) );
  NAND2_X1 U732 ( .A1(n646), .A2(n645), .ZN(n651) );
  NAND2_X1 U733 ( .A1(G80), .A2(n670), .ZN(n647) );
  XNOR2_X1 U734 ( .A(n647), .B(KEYINPUT82), .ZN(n649) );
  NAND2_X1 U735 ( .A1(G67), .A2(n675), .ZN(n648) );
  NAND2_X1 U736 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U737 ( .A1(n651), .A2(n650), .ZN(n686) );
  XOR2_X1 U738 ( .A(n652), .B(n686), .Z(G145) );
  INV_X1 U739 ( .A(G303), .ZN(G166) );
  NAND2_X1 U740 ( .A1(G47), .A2(n666), .ZN(n654) );
  NAND2_X1 U741 ( .A1(G85), .A2(n667), .ZN(n653) );
  NAND2_X1 U742 ( .A1(n654), .A2(n653), .ZN(n657) );
  NAND2_X1 U743 ( .A1(G60), .A2(n675), .ZN(n655) );
  XNOR2_X1 U744 ( .A(KEYINPUT67), .B(n655), .ZN(n656) );
  NOR2_X1 U745 ( .A1(n657), .A2(n656), .ZN(n659) );
  NAND2_X1 U746 ( .A1(G72), .A2(n670), .ZN(n658) );
  NAND2_X1 U747 ( .A1(n659), .A2(n658), .ZN(G290) );
  NAND2_X1 U748 ( .A1(G87), .A2(n660), .ZN(n662) );
  NAND2_X1 U749 ( .A1(G74), .A2(G651), .ZN(n661) );
  NAND2_X1 U750 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U751 ( .A1(n675), .A2(n663), .ZN(n665) );
  NAND2_X1 U752 ( .A1(n666), .A2(G49), .ZN(n664) );
  NAND2_X1 U753 ( .A1(n665), .A2(n664), .ZN(G288) );
  NAND2_X1 U754 ( .A1(G48), .A2(n666), .ZN(n669) );
  NAND2_X1 U755 ( .A1(G86), .A2(n667), .ZN(n668) );
  NAND2_X1 U756 ( .A1(n669), .A2(n668), .ZN(n674) );
  NAND2_X1 U757 ( .A1(n670), .A2(G73), .ZN(n671) );
  XNOR2_X1 U758 ( .A(n671), .B(KEYINPUT83), .ZN(n672) );
  XNOR2_X1 U759 ( .A(n672), .B(KEYINPUT2), .ZN(n673) );
  NOR2_X1 U760 ( .A1(n674), .A2(n673), .ZN(n677) );
  NAND2_X1 U761 ( .A1(G61), .A2(n675), .ZN(n676) );
  NAND2_X1 U762 ( .A1(n677), .A2(n676), .ZN(G305) );
  XOR2_X1 U763 ( .A(G299), .B(G166), .Z(n682) );
  XNOR2_X1 U764 ( .A(n686), .B(G290), .ZN(n680) );
  XOR2_X1 U765 ( .A(KEYINPUT19), .B(G305), .Z(n678) );
  XNOR2_X1 U766 ( .A(G288), .B(n678), .ZN(n679) );
  XNOR2_X1 U767 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U768 ( .A(n682), .B(n681), .ZN(n905) );
  XNOR2_X1 U769 ( .A(n905), .B(n683), .ZN(n684) );
  NAND2_X1 U770 ( .A1(n684), .A2(G868), .ZN(n685) );
  XOR2_X1 U771 ( .A(KEYINPUT85), .B(n685), .Z(n688) );
  OR2_X1 U772 ( .A1(n686), .A2(G868), .ZN(n687) );
  NAND2_X1 U773 ( .A1(n688), .A2(n687), .ZN(G295) );
  NAND2_X1 U774 ( .A1(G2078), .A2(G2084), .ZN(n689) );
  XOR2_X1 U775 ( .A(KEYINPUT20), .B(n689), .Z(n690) );
  NAND2_X1 U776 ( .A1(G2090), .A2(n690), .ZN(n691) );
  XNOR2_X1 U777 ( .A(KEYINPUT21), .B(n691), .ZN(n692) );
  NAND2_X1 U778 ( .A1(n692), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U779 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U780 ( .A(KEYINPUT74), .B(G82), .Z(G220) );
  NAND2_X1 U781 ( .A1(G483), .A2(G661), .ZN(n700) );
  NOR2_X1 U782 ( .A1(G220), .A2(G219), .ZN(n693) );
  XOR2_X1 U783 ( .A(KEYINPUT22), .B(n693), .Z(n694) );
  NOR2_X1 U784 ( .A1(G218), .A2(n694), .ZN(n695) );
  NAND2_X1 U785 ( .A1(G96), .A2(n695), .ZN(n925) );
  NAND2_X1 U786 ( .A1(n925), .A2(G2106), .ZN(n699) );
  NAND2_X1 U787 ( .A1(G69), .A2(G120), .ZN(n696) );
  NOR2_X1 U788 ( .A1(G237), .A2(n696), .ZN(n697) );
  NAND2_X1 U789 ( .A1(G108), .A2(n697), .ZN(n926) );
  NAND2_X1 U790 ( .A1(n926), .A2(G567), .ZN(n698) );
  NAND2_X1 U791 ( .A1(n699), .A2(n698), .ZN(n840) );
  NOR2_X1 U792 ( .A1(n700), .A2(n840), .ZN(n701) );
  XNOR2_X1 U793 ( .A(n701), .B(KEYINPUT86), .ZN(n839) );
  NAND2_X1 U794 ( .A1(G36), .A2(n839), .ZN(G176) );
  XNOR2_X1 U795 ( .A(G1981), .B(G305), .ZN(n982) );
  NAND2_X1 U796 ( .A1(G160), .A2(G40), .ZN(n786) );
  INV_X1 U797 ( .A(n720), .ZN(n711) );
  NOR2_X1 U798 ( .A1(G2090), .A2(n711), .ZN(n702) );
  XOR2_X1 U799 ( .A(KEYINPUT101), .B(n702), .Z(n705) );
  INV_X1 U800 ( .A(n765), .ZN(n813) );
  NOR2_X1 U801 ( .A1(G1971), .A2(n813), .ZN(n704) );
  NOR2_X1 U802 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U803 ( .A1(n706), .A2(G303), .ZN(n749) );
  NOR2_X1 U804 ( .A1(G2084), .A2(n730), .ZN(n752) );
  NAND2_X1 U805 ( .A1(G8), .A2(n707), .ZN(n709) );
  XNOR2_X1 U806 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X1 U807 ( .A1(G168), .A2(n710), .ZN(n715) );
  XNOR2_X1 U808 ( .A(G2078), .B(KEYINPUT25), .ZN(n965) );
  NOR2_X1 U809 ( .A1(n711), .A2(n965), .ZN(n713) );
  XOR2_X1 U810 ( .A(G1961), .B(KEYINPUT98), .Z(n1004) );
  NOR2_X1 U811 ( .A1(n720), .A2(n1004), .ZN(n712) );
  NOR2_X1 U812 ( .A1(n713), .A2(n712), .ZN(n718) );
  NOR2_X1 U813 ( .A1(G171), .A2(n718), .ZN(n714) );
  XNOR2_X1 U814 ( .A(n717), .B(n716), .ZN(n748) );
  NAND2_X1 U815 ( .A1(n718), .A2(G171), .ZN(n746) );
  XNOR2_X1 U816 ( .A(KEYINPUT99), .B(KEYINPUT29), .ZN(n744) );
  NAND2_X1 U817 ( .A1(n720), .A2(G2072), .ZN(n719) );
  XNOR2_X1 U818 ( .A(n719), .B(KEYINPUT27), .ZN(n722) );
  INV_X1 U819 ( .A(G1956), .ZN(n846) );
  NOR2_X1 U820 ( .A1(n846), .A2(n720), .ZN(n721) );
  NOR2_X1 U821 ( .A1(n722), .A2(n721), .ZN(n724) );
  NOR2_X1 U822 ( .A1(n725), .A2(n724), .ZN(n723) );
  XOR2_X1 U823 ( .A(n723), .B(KEYINPUT28), .Z(n742) );
  NAND2_X1 U824 ( .A1(n725), .A2(n724), .ZN(n740) );
  INV_X1 U825 ( .A(G1996), .ZN(n956) );
  NOR2_X1 U826 ( .A1(n730), .A2(n956), .ZN(n726) );
  XOR2_X1 U827 ( .A(n726), .B(KEYINPUT26), .Z(n728) );
  NAND2_X1 U828 ( .A1(n730), .A2(G1341), .ZN(n727) );
  NAND2_X1 U829 ( .A1(n728), .A2(n727), .ZN(n729) );
  NOR2_X1 U830 ( .A1(n997), .A2(n729), .ZN(n734) );
  INV_X1 U831 ( .A(n990), .ZN(n736) );
  NAND2_X1 U832 ( .A1(G1348), .A2(n730), .ZN(n732) );
  NAND2_X1 U833 ( .A1(G2067), .A2(n720), .ZN(n731) );
  NAND2_X1 U834 ( .A1(n732), .A2(n731), .ZN(n735) );
  NOR2_X1 U835 ( .A1(n736), .A2(n735), .ZN(n733) );
  OR2_X1 U836 ( .A1(n734), .A2(n733), .ZN(n738) );
  NAND2_X1 U837 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U838 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U839 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U840 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U841 ( .A(n744), .B(n743), .ZN(n745) );
  NAND2_X1 U842 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U843 ( .A1(n750), .A2(G8), .ZN(n751) );
  XNOR2_X1 U844 ( .A(n751), .B(KEYINPUT32), .ZN(n759) );
  NAND2_X1 U845 ( .A1(G8), .A2(n752), .ZN(n753) );
  XNOR2_X1 U846 ( .A(KEYINPUT97), .B(n753), .ZN(n754) );
  NOR2_X1 U847 ( .A1(n755), .A2(n754), .ZN(n757) );
  NAND2_X1 U848 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U849 ( .A1(n759), .A2(n758), .ZN(n811) );
  NOR2_X1 U850 ( .A1(G1976), .A2(G288), .ZN(n985) );
  NOR2_X1 U851 ( .A1(G1971), .A2(G303), .ZN(n760) );
  XOR2_X1 U852 ( .A(n760), .B(KEYINPUT103), .Z(n761) );
  NOR2_X1 U853 ( .A1(n985), .A2(n761), .ZN(n762) );
  NAND2_X1 U854 ( .A1(n811), .A2(n762), .ZN(n763) );
  NAND2_X1 U855 ( .A1(G1976), .A2(G288), .ZN(n988) );
  AND2_X1 U856 ( .A1(n988), .A2(n765), .ZN(n764) );
  AND2_X1 U857 ( .A1(n985), .A2(KEYINPUT33), .ZN(n766) );
  NAND2_X1 U858 ( .A1(n766), .A2(n765), .ZN(n802) );
  NAND2_X1 U859 ( .A1(G119), .A2(n880), .ZN(n767) );
  XNOR2_X1 U860 ( .A(n767), .B(KEYINPUT90), .ZN(n774) );
  NAND2_X1 U861 ( .A1(G95), .A2(n886), .ZN(n769) );
  NAND2_X1 U862 ( .A1(G131), .A2(n884), .ZN(n768) );
  NAND2_X1 U863 ( .A1(n769), .A2(n768), .ZN(n772) );
  NAND2_X1 U864 ( .A1(G107), .A2(n881), .ZN(n770) );
  XNOR2_X1 U865 ( .A(KEYINPUT91), .B(n770), .ZN(n771) );
  NOR2_X1 U866 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U867 ( .A1(n774), .A2(n773), .ZN(n898) );
  AND2_X1 U868 ( .A1(n898), .A2(G1991), .ZN(n785) );
  NAND2_X1 U869 ( .A1(G129), .A2(n880), .ZN(n776) );
  NAND2_X1 U870 ( .A1(G117), .A2(n881), .ZN(n775) );
  NAND2_X1 U871 ( .A1(n776), .A2(n775), .ZN(n779) );
  NAND2_X1 U872 ( .A1(n886), .A2(G105), .ZN(n777) );
  XOR2_X1 U873 ( .A(KEYINPUT38), .B(n777), .Z(n778) );
  NOR2_X1 U874 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U875 ( .A(n780), .B(KEYINPUT92), .ZN(n782) );
  NAND2_X1 U876 ( .A1(G141), .A2(n884), .ZN(n781) );
  NAND2_X1 U877 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U878 ( .A(KEYINPUT93), .B(n783), .ZN(n877) );
  NOR2_X1 U879 ( .A1(n877), .A2(n956), .ZN(n784) );
  NOR2_X1 U880 ( .A1(n785), .A2(n784), .ZN(n944) );
  INV_X1 U881 ( .A(n786), .ZN(n788) );
  NAND2_X1 U882 ( .A1(n788), .A2(n787), .ZN(n789) );
  NOR2_X1 U883 ( .A1(n944), .A2(n789), .ZN(n825) );
  XOR2_X1 U884 ( .A(KEYINPUT94), .B(n825), .Z(n801) );
  INV_X1 U885 ( .A(n789), .ZN(n833) );
  XNOR2_X1 U886 ( .A(KEYINPUT88), .B(KEYINPUT34), .ZN(n793) );
  NAND2_X1 U887 ( .A1(G104), .A2(n886), .ZN(n791) );
  NAND2_X1 U888 ( .A1(G140), .A2(n884), .ZN(n790) );
  NAND2_X1 U889 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U890 ( .A(n793), .B(n792), .ZN(n799) );
  XNOR2_X1 U891 ( .A(KEYINPUT35), .B(KEYINPUT89), .ZN(n797) );
  NAND2_X1 U892 ( .A1(G128), .A2(n880), .ZN(n795) );
  NAND2_X1 U893 ( .A1(G116), .A2(n881), .ZN(n794) );
  NAND2_X1 U894 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U895 ( .A(n797), .B(n796), .ZN(n798) );
  NOR2_X1 U896 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U897 ( .A(n800), .B(KEYINPUT36), .ZN(n897) );
  XNOR2_X1 U898 ( .A(KEYINPUT37), .B(G2067), .ZN(n831) );
  NOR2_X1 U899 ( .A1(n897), .A2(n831), .ZN(n933) );
  NAND2_X1 U900 ( .A1(n833), .A2(n933), .ZN(n829) );
  AND2_X1 U901 ( .A1(n801), .A2(n829), .ZN(n805) );
  AND2_X1 U902 ( .A1(n802), .A2(n805), .ZN(n803) );
  NAND2_X1 U903 ( .A1(n804), .A2(n803), .ZN(n820) );
  INV_X1 U904 ( .A(n805), .ZN(n818) );
  NOR2_X1 U905 ( .A1(G1981), .A2(G305), .ZN(n806) );
  XNOR2_X1 U906 ( .A(n806), .B(KEYINPUT96), .ZN(n807) );
  XNOR2_X1 U907 ( .A(n807), .B(KEYINPUT24), .ZN(n808) );
  AND2_X1 U908 ( .A1(n808), .A2(n765), .ZN(n816) );
  NOR2_X1 U909 ( .A1(G2090), .A2(G303), .ZN(n809) );
  NAND2_X1 U910 ( .A1(G8), .A2(n809), .ZN(n810) );
  NAND2_X1 U911 ( .A1(n811), .A2(n810), .ZN(n812) );
  NAND2_X1 U912 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U913 ( .A(KEYINPUT105), .B(n814), .ZN(n815) );
  NOR2_X1 U914 ( .A1(n816), .A2(n815), .ZN(n817) );
  OR2_X1 U915 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U916 ( .A(G1986), .B(G290), .ZN(n987) );
  NAND2_X1 U917 ( .A1(n987), .A2(n833), .ZN(n821) );
  XOR2_X1 U918 ( .A(KEYINPUT107), .B(KEYINPUT39), .Z(n822) );
  XNOR2_X1 U919 ( .A(KEYINPUT106), .B(n822), .ZN(n828) );
  AND2_X1 U920 ( .A1(n956), .A2(n877), .ZN(n946) );
  NOR2_X1 U921 ( .A1(G1986), .A2(G290), .ZN(n823) );
  NOR2_X1 U922 ( .A1(G1991), .A2(n898), .ZN(n929) );
  NOR2_X1 U923 ( .A1(n823), .A2(n929), .ZN(n824) );
  NOR2_X1 U924 ( .A1(n825), .A2(n824), .ZN(n826) );
  NOR2_X1 U925 ( .A1(n946), .A2(n826), .ZN(n827) );
  XNOR2_X1 U926 ( .A(n828), .B(n827), .ZN(n830) );
  NAND2_X1 U927 ( .A1(n830), .A2(n829), .ZN(n832) );
  NAND2_X1 U928 ( .A1(n897), .A2(n831), .ZN(n934) );
  NAND2_X1 U929 ( .A1(n832), .A2(n934), .ZN(n834) );
  NAND2_X1 U930 ( .A1(n834), .A2(n833), .ZN(n835) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n836), .ZN(G217) );
  INV_X1 U932 ( .A(n836), .ZN(G223) );
  AND2_X1 U933 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U934 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U936 ( .A1(n839), .A2(n838), .ZN(G188) );
  INV_X1 U937 ( .A(n840), .ZN(G319) );
  XOR2_X1 U938 ( .A(KEYINPUT110), .B(G1986), .Z(n842) );
  XOR2_X1 U939 ( .A(n956), .B(G1991), .Z(n841) );
  XNOR2_X1 U940 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U941 ( .A(n843), .B(KEYINPUT109), .Z(n845) );
  XNOR2_X1 U942 ( .A(G1976), .B(G1966), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(n850) );
  XOR2_X1 U944 ( .A(G1971), .B(G1961), .Z(n848) );
  XOR2_X1 U945 ( .A(G1981), .B(n846), .Z(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U947 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U948 ( .A(G2474), .B(KEYINPUT41), .ZN(n851) );
  XNOR2_X1 U949 ( .A(n852), .B(n851), .ZN(G229) );
  XOR2_X1 U950 ( .A(G2100), .B(KEYINPUT43), .Z(n854) );
  XNOR2_X1 U951 ( .A(G2067), .B(KEYINPUT108), .ZN(n853) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U953 ( .A(n855), .B(G2678), .Z(n857) );
  XNOR2_X1 U954 ( .A(G2072), .B(G2090), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U956 ( .A(KEYINPUT42), .B(G2096), .Z(n859) );
  XNOR2_X1 U957 ( .A(G2078), .B(G2084), .ZN(n858) );
  XNOR2_X1 U958 ( .A(n859), .B(n858), .ZN(n860) );
  XNOR2_X1 U959 ( .A(n861), .B(n860), .ZN(G227) );
  NAND2_X1 U960 ( .A1(n880), .A2(G124), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n862), .B(KEYINPUT44), .ZN(n864) );
  NAND2_X1 U962 ( .A1(G100), .A2(n886), .ZN(n863) );
  NAND2_X1 U963 ( .A1(n864), .A2(n863), .ZN(n868) );
  NAND2_X1 U964 ( .A1(G136), .A2(n884), .ZN(n866) );
  NAND2_X1 U965 ( .A1(G112), .A2(n881), .ZN(n865) );
  NAND2_X1 U966 ( .A1(n866), .A2(n865), .ZN(n867) );
  NOR2_X1 U967 ( .A1(n868), .A2(n867), .ZN(G162) );
  NAND2_X1 U968 ( .A1(G127), .A2(n880), .ZN(n870) );
  NAND2_X1 U969 ( .A1(G115), .A2(n881), .ZN(n869) );
  NAND2_X1 U970 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n871), .B(KEYINPUT47), .ZN(n873) );
  NAND2_X1 U972 ( .A1(G139), .A2(n884), .ZN(n872) );
  NAND2_X1 U973 ( .A1(n873), .A2(n872), .ZN(n876) );
  NAND2_X1 U974 ( .A1(G103), .A2(n886), .ZN(n874) );
  XNOR2_X1 U975 ( .A(KEYINPUT113), .B(n874), .ZN(n875) );
  NOR2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n936) );
  XOR2_X1 U977 ( .A(n928), .B(n936), .Z(n879) );
  XNOR2_X1 U978 ( .A(G164), .B(n877), .ZN(n878) );
  XNOR2_X1 U979 ( .A(n879), .B(n878), .ZN(n894) );
  NAND2_X1 U980 ( .A1(G130), .A2(n880), .ZN(n883) );
  NAND2_X1 U981 ( .A1(G118), .A2(n881), .ZN(n882) );
  NAND2_X1 U982 ( .A1(n883), .A2(n882), .ZN(n892) );
  NAND2_X1 U983 ( .A1(n884), .A2(G142), .ZN(n885) );
  XNOR2_X1 U984 ( .A(KEYINPUT112), .B(n885), .ZN(n889) );
  NAND2_X1 U985 ( .A1(n886), .A2(G106), .ZN(n887) );
  XOR2_X1 U986 ( .A(KEYINPUT111), .B(n887), .Z(n888) );
  NAND2_X1 U987 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U988 ( .A(n890), .B(KEYINPUT45), .Z(n891) );
  NOR2_X1 U989 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U990 ( .A(n894), .B(n893), .Z(n903) );
  XOR2_X1 U991 ( .A(KEYINPUT48), .B(KEYINPUT114), .Z(n896) );
  XNOR2_X1 U992 ( .A(G162), .B(KEYINPUT46), .ZN(n895) );
  XNOR2_X1 U993 ( .A(n896), .B(n895), .ZN(n901) );
  XNOR2_X1 U994 ( .A(G160), .B(n897), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U996 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U997 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U998 ( .A1(G37), .A2(n904), .ZN(G395) );
  XNOR2_X1 U999 ( .A(G286), .B(n905), .ZN(n907) );
  XNOR2_X1 U1000 ( .A(n997), .B(G171), .ZN(n906) );
  XNOR2_X1 U1001 ( .A(n907), .B(n906), .ZN(n909) );
  XOR2_X1 U1002 ( .A(n990), .B(KEYINPUT115), .Z(n908) );
  XNOR2_X1 U1003 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n910), .ZN(G397) );
  XOR2_X1 U1005 ( .A(G2451), .B(G2430), .Z(n912) );
  XNOR2_X1 U1006 ( .A(G2438), .B(G2443), .ZN(n911) );
  XNOR2_X1 U1007 ( .A(n912), .B(n911), .ZN(n918) );
  XOR2_X1 U1008 ( .A(G2435), .B(G2454), .Z(n914) );
  XNOR2_X1 U1009 ( .A(G1341), .B(G1348), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(n914), .B(n913), .ZN(n916) );
  XOR2_X1 U1011 ( .A(G2446), .B(G2427), .Z(n915) );
  XNOR2_X1 U1012 ( .A(n916), .B(n915), .ZN(n917) );
  XOR2_X1 U1013 ( .A(n918), .B(n917), .Z(n919) );
  NAND2_X1 U1014 ( .A1(G14), .A2(n919), .ZN(n927) );
  NAND2_X1 U1015 ( .A1(G319), .A2(n927), .ZN(n922) );
  NOR2_X1 U1016 ( .A1(G229), .A2(G227), .ZN(n920) );
  XNOR2_X1 U1017 ( .A(KEYINPUT49), .B(n920), .ZN(n921) );
  NOR2_X1 U1018 ( .A1(n922), .A2(n921), .ZN(n924) );
  NOR2_X1 U1019 ( .A1(G395), .A2(G397), .ZN(n923) );
  NAND2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(G225) );
  XOR2_X1 U1021 ( .A(KEYINPUT116), .B(G225), .Z(G308) );
  INV_X1 U1023 ( .A(G120), .ZN(G236) );
  INV_X1 U1024 ( .A(G96), .ZN(G221) );
  INV_X1 U1025 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(G325) );
  INV_X1 U1027 ( .A(G325), .ZN(G261) );
  INV_X1 U1028 ( .A(G108), .ZN(G238) );
  INV_X1 U1029 ( .A(n927), .ZN(G401) );
  XNOR2_X1 U1030 ( .A(G160), .B(G2084), .ZN(n931) );
  NOR2_X1 U1031 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1032 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1033 ( .A1(n933), .A2(n932), .ZN(n935) );
  NAND2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n942) );
  XOR2_X1 U1035 ( .A(G2072), .B(n936), .Z(n938) );
  XOR2_X1 U1036 ( .A(G164), .B(G2078), .Z(n937) );
  NOR2_X1 U1037 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1038 ( .A(KEYINPUT50), .B(n939), .Z(n940) );
  XNOR2_X1 U1039 ( .A(KEYINPUT118), .B(n940), .ZN(n941) );
  NOR2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n950) );
  XOR2_X1 U1042 ( .A(G2090), .B(G162), .Z(n945) );
  NOR2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1044 ( .A(KEYINPUT117), .B(n947), .Z(n948) );
  XNOR2_X1 U1045 ( .A(KEYINPUT51), .B(n948), .ZN(n949) );
  NOR2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1047 ( .A(KEYINPUT52), .B(n951), .ZN(n952) );
  XNOR2_X1 U1048 ( .A(KEYINPUT55), .B(KEYINPUT119), .ZN(n954) );
  NAND2_X1 U1049 ( .A1(n952), .A2(n954), .ZN(n953) );
  NAND2_X1 U1050 ( .A1(n953), .A2(G29), .ZN(n1034) );
  XNOR2_X1 U1051 ( .A(G29), .B(KEYINPUT123), .ZN(n977) );
  XNOR2_X1 U1052 ( .A(n954), .B(KEYINPUT122), .ZN(n975) );
  XNOR2_X1 U1053 ( .A(G2090), .B(G35), .ZN(n970) );
  XNOR2_X1 U1054 ( .A(KEYINPUT121), .B(G2072), .ZN(n955) );
  XNOR2_X1 U1055 ( .A(n955), .B(G33), .ZN(n964) );
  XOR2_X1 U1056 ( .A(n956), .B(G32), .Z(n958) );
  XNOR2_X1 U1057 ( .A(G1991), .B(G25), .ZN(n957) );
  NOR2_X1 U1058 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1059 ( .A1(G28), .A2(n959), .ZN(n962) );
  XNOR2_X1 U1060 ( .A(KEYINPUT120), .B(G2067), .ZN(n960) );
  XNOR2_X1 U1061 ( .A(G26), .B(n960), .ZN(n961) );
  NOR2_X1 U1062 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1063 ( .A1(n964), .A2(n963), .ZN(n967) );
  XOR2_X1 U1064 ( .A(G27), .B(n965), .Z(n966) );
  NOR2_X1 U1065 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1066 ( .A(KEYINPUT53), .B(n968), .ZN(n969) );
  NOR2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n973) );
  XOR2_X1 U1068 ( .A(G2084), .B(G34), .Z(n971) );
  XNOR2_X1 U1069 ( .A(KEYINPUT54), .B(n971), .ZN(n972) );
  NAND2_X1 U1070 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1071 ( .A(n975), .B(n974), .ZN(n976) );
  NAND2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1073 ( .A1(n978), .A2(G11), .ZN(n1032) );
  INV_X1 U1074 ( .A(G16), .ZN(n1028) );
  XOR2_X1 U1075 ( .A(n1028), .B(KEYINPUT56), .Z(n1003) );
  XOR2_X1 U1076 ( .A(G171), .B(G1961), .Z(n980) );
  XNOR2_X1 U1077 ( .A(G299), .B(G1956), .ZN(n979) );
  NOR2_X1 U1078 ( .A1(n980), .A2(n979), .ZN(n1001) );
  XOR2_X1 U1079 ( .A(G1966), .B(G168), .Z(n981) );
  NOR2_X1 U1080 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1081 ( .A(KEYINPUT57), .B(n983), .Z(n984) );
  XNOR2_X1 U1082 ( .A(KEYINPUT124), .B(n984), .ZN(n996) );
  XOR2_X1 U1083 ( .A(n985), .B(KEYINPUT125), .Z(n986) );
  NOR2_X1 U1084 ( .A1(n987), .A2(n986), .ZN(n989) );
  NAND2_X1 U1085 ( .A1(n989), .A2(n988), .ZN(n994) );
  XNOR2_X1 U1086 ( .A(n990), .B(G1348), .ZN(n992) );
  XOR2_X1 U1087 ( .A(G303), .B(G1971), .Z(n991) );
  NAND2_X1 U1088 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1089 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1090 ( .A1(n996), .A2(n995), .ZN(n999) );
  XNOR2_X1 U1091 ( .A(G1341), .B(n997), .ZN(n998) );
  NOR2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1030) );
  XNOR2_X1 U1095 ( .A(n1004), .B(G5), .ZN(n1018) );
  XNOR2_X1 U1096 ( .A(KEYINPUT127), .B(G1341), .ZN(n1005) );
  XNOR2_X1 U1097 ( .A(n1005), .B(G19), .ZN(n1010) );
  XOR2_X1 U1098 ( .A(G1348), .B(KEYINPUT59), .Z(n1006) );
  XNOR2_X1 U1099 ( .A(G4), .B(n1006), .ZN(n1008) );
  XNOR2_X1 U1100 ( .A(G6), .B(G1981), .ZN(n1007) );
  NOR2_X1 U1101 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1102 ( .A1(n1010), .A2(n1009), .ZN(n1013) );
  XNOR2_X1 U1103 ( .A(G20), .B(G1956), .ZN(n1011) );
  XNOR2_X1 U1104 ( .A(KEYINPUT126), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1105 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1106 ( .A(KEYINPUT60), .B(n1014), .Z(n1016) );
  XNOR2_X1 U1107 ( .A(G1966), .B(G21), .ZN(n1015) );
  NOR2_X1 U1108 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1109 ( .A1(n1018), .A2(n1017), .ZN(n1025) );
  XNOR2_X1 U1110 ( .A(G1976), .B(G23), .ZN(n1020) );
  XNOR2_X1 U1111 ( .A(G1971), .B(G22), .ZN(n1019) );
  NOR2_X1 U1112 ( .A1(n1020), .A2(n1019), .ZN(n1022) );
  XOR2_X1 U1113 ( .A(G1986), .B(G24), .Z(n1021) );
  NAND2_X1 U1114 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1115 ( .A(KEYINPUT58), .B(n1023), .ZN(n1024) );
  NOR2_X1 U1116 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1117 ( .A(KEYINPUT61), .B(n1026), .ZN(n1027) );
  NAND2_X1 U1118 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1119 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NOR2_X1 U1120 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1121 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XNOR2_X1 U1122 ( .A(KEYINPUT62), .B(n1035), .ZN(G150) );
  INV_X1 U1123 ( .A(G150), .ZN(G311) );
endmodule

