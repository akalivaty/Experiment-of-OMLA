//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 1 0 1 1 0 1 0 1 0 1 0 1 0 1 0 1 1 1 0 1 0 0 1 1 1 0 1 0 1 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1275, new_n1276, new_n1277, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G50), .ZN(new_n205));
  INV_X1    g0005(.A(KEYINPUT64), .ZN(new_n206));
  AOI21_X1  g0006(.A(new_n205), .B1(new_n202), .B2(new_n206), .ZN(new_n207));
  OAI21_X1  g0007(.A(new_n207), .B1(new_n206), .B2(new_n202), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT65), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G1), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n211), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(G13), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT0), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT67), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT66), .Z(new_n226));
  OAI21_X1  g0026(.A(new_n216), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n213), .B(new_n219), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT68), .Z(G361));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT69), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n234), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  XOR2_X1   g0046(.A(KEYINPUT8), .B(G58), .Z(new_n247));
  NAND2_X1  g0047(.A1(new_n214), .A2(G20), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n210), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G13), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(G1), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G20), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  OAI22_X1  g0056(.A1(new_n249), .A2(new_n256), .B1(new_n255), .B2(new_n247), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G200), .ZN(new_n259));
  AND2_X1   g0059(.A1(G1), .A2(G13), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(G1698), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n264), .A2(new_n266), .A3(G223), .A4(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT81), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT3), .B(G33), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n271), .A2(KEYINPUT81), .A3(G223), .A4(new_n267), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n264), .A2(new_n266), .A3(G226), .A4(G1698), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G87), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n262), .B1(new_n273), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G274), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n279), .B1(new_n260), .B2(new_n261), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n214), .B1(G41), .B2(G45), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n262), .A2(new_n281), .ZN(new_n284));
  INV_X1    g0084(.A(G232), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n259), .B1(new_n278), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n286), .ZN(new_n288));
  INV_X1    g0088(.A(G190), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n276), .B1(new_n270), .B2(new_n272), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n288), .B(new_n289), .C1(new_n290), .C2(new_n262), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G58), .ZN(new_n293));
  INV_X1    g0093(.A(G68), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(G20), .B1(new_n295), .B2(new_n201), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G20), .A2(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G159), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n296), .A2(KEYINPUT16), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n264), .A2(new_n266), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n300), .A2(KEYINPUT79), .A3(KEYINPUT7), .A4(new_n211), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT7), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n302), .B1(new_n271), .B2(G20), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(G20), .B1(new_n264), .B2(new_n266), .ZN(new_n305));
  AOI21_X1  g0105(.A(KEYINPUT79), .B1(new_n305), .B2(KEYINPUT7), .ZN(new_n306));
  OAI21_X1  g0106(.A(G68), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT80), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT80), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n309), .B(G68), .C1(new_n304), .C2(new_n306), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n299), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n296), .A2(new_n298), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n265), .A2(G33), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n314));
  OAI211_X1 g0114(.A(KEYINPUT7), .B(new_n211), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n303), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n312), .B1(new_n316), .B2(G68), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n251), .B1(new_n317), .B2(KEYINPUT16), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n258), .B(new_n292), .C1(new_n311), .C2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT82), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n299), .ZN(new_n322));
  INV_X1    g0122(.A(new_n310), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT79), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n315), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n325), .A2(new_n301), .A3(new_n303), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n309), .B1(new_n326), .B2(G68), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n322), .B1(new_n323), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n318), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n330), .A2(KEYINPUT82), .A3(new_n258), .A4(new_n292), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n321), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT17), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n257), .B1(new_n328), .B2(new_n329), .ZN(new_n334));
  OAI21_X1  g0134(.A(G169), .B1(new_n278), .B2(new_n286), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n288), .B(G179), .C1(new_n290), .C2(new_n262), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NOR3_X1   g0138(.A1(new_n334), .A2(KEYINPUT18), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT18), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n258), .B1(new_n311), .B2(new_n318), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n340), .B1(new_n341), .B2(new_n337), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n319), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n344), .A2(KEYINPUT17), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n333), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT77), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n271), .A2(G226), .A3(new_n267), .ZN(new_n349));
  AND3_X1   g0149(.A1(KEYINPUT75), .A2(G33), .A3(G97), .ZN(new_n350));
  AOI21_X1  g0150(.A(KEYINPUT75), .B1(G33), .B2(G97), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n264), .A2(new_n266), .A3(G232), .A4(G1698), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n349), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n262), .A2(G238), .A3(new_n281), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n283), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n360), .A2(KEYINPUT76), .A3(KEYINPUT13), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT76), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n358), .B1(new_n354), .B2(new_n355), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT13), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(new_n364), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n361), .A2(new_n365), .A3(G190), .A4(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  AOI211_X1 g0168(.A(KEYINPUT13), .B(new_n358), .C1(new_n355), .C2(new_n354), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n364), .B1(new_n356), .B2(new_n359), .ZN(new_n370));
  OAI21_X1  g0170(.A(G200), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT72), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n252), .A2(new_n255), .A3(new_n372), .ZN(new_n373));
  NOR3_X1   g0173(.A1(new_n253), .A2(new_n211), .A3(G1), .ZN(new_n374));
  OAI21_X1  g0174(.A(KEYINPUT72), .B1(new_n374), .B2(new_n251), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n376), .A2(G68), .A3(new_n248), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n297), .A2(G50), .B1(G20), .B2(new_n294), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n263), .A2(G20), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(G77), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n378), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n251), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT11), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n374), .A2(new_n294), .ZN(new_n386));
  XNOR2_X1  g0186(.A(new_n386), .B(KEYINPUT12), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n382), .A2(KEYINPUT11), .A3(new_n251), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n377), .A2(new_n385), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n371), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n348), .B1(new_n368), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n370), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n366), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n389), .B1(new_n394), .B2(G200), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n395), .A2(KEYINPUT77), .A3(new_n367), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(G169), .B1(new_n369), .B2(new_n370), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n398), .A2(KEYINPUT78), .A3(KEYINPUT14), .ZN(new_n399));
  NAND2_X1  g0199(.A1(KEYINPUT78), .A2(KEYINPUT14), .ZN(new_n400));
  OAI211_X1 g0200(.A(G169), .B(new_n400), .C1(new_n369), .C2(new_n370), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n361), .A2(new_n365), .A3(G179), .A4(new_n366), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n399), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n389), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n397), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n248), .A2(G50), .ZN(new_n406));
  OAI22_X1  g0206(.A1(new_n256), .A2(new_n406), .B1(G50), .B2(new_n255), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n211), .B1(new_n201), .B2(new_n205), .ZN(new_n409));
  INV_X1    g0209(.A(new_n297), .ZN(new_n410));
  INV_X1    g0210(.A(G150), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI211_X1 g0212(.A(new_n409), .B(new_n412), .C1(new_n247), .C2(new_n379), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n408), .B1(new_n252), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g0214(.A(new_n414), .B(KEYINPUT9), .ZN(new_n415));
  INV_X1    g0215(.A(G226), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n283), .B1(new_n284), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n271), .A2(G223), .A3(G1698), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n271), .A2(new_n267), .ZN(new_n419));
  INV_X1    g0219(.A(G222), .ZN(new_n420));
  OAI221_X1 g0220(.A(new_n418), .B1(new_n381), .B2(new_n271), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n417), .B1(new_n421), .B2(new_n355), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n289), .ZN(new_n423));
  XOR2_X1   g0223(.A(KEYINPUT73), .B(G200), .Z(new_n424));
  OAI21_X1  g0224(.A(new_n423), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n415), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(KEYINPUT10), .B1(new_n425), .B2(KEYINPUT74), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n415), .B(new_n425), .C1(KEYINPUT74), .C2(KEYINPUT10), .ZN(new_n429));
  INV_X1    g0229(.A(G179), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n422), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n431), .B(new_n414), .C1(G169), .C2(new_n422), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n428), .A2(new_n429), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n271), .A2(G238), .A3(G1698), .ZN(new_n434));
  INV_X1    g0234(.A(G107), .ZN(new_n435));
  OAI221_X1 g0235(.A(new_n434), .B1(new_n435), .B2(new_n271), .C1(new_n419), .C2(new_n285), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n436), .A2(new_n355), .ZN(new_n437));
  INV_X1    g0237(.A(G244), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n283), .B1(new_n284), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n424), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n376), .A2(G77), .A3(new_n248), .ZN(new_n441));
  XNOR2_X1  g0241(.A(KEYINPUT15), .B(G87), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n443), .A2(new_n379), .B1(G20), .B2(G77), .ZN(new_n444));
  OR2_X1    g0244(.A1(new_n297), .A2(KEYINPUT70), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n297), .A2(KEYINPUT70), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n247), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n252), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n374), .A2(new_n381), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n449), .B(KEYINPUT71), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n439), .B1(new_n436), .B2(new_n355), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G190), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n440), .A2(new_n441), .A3(new_n451), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n451), .A2(new_n441), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n452), .A2(new_n430), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n455), .B(new_n456), .C1(G169), .C2(new_n452), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  NOR4_X1   g0258(.A1(new_n347), .A2(new_n405), .A3(new_n433), .A4(new_n458), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n264), .A2(new_n266), .A3(new_n211), .A4(G87), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT22), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT22), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n271), .A2(new_n462), .A3(new_n211), .A4(G87), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT24), .ZN(new_n465));
  INV_X1    g0265(.A(G116), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n263), .A2(new_n466), .A3(G20), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT23), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(new_n211), .B2(G107), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n435), .A2(KEYINPUT23), .A3(G20), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n467), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AND3_X1   g0271(.A1(new_n464), .A2(new_n465), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n465), .B1(new_n464), .B2(new_n471), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n251), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n256), .B1(new_n214), .B2(G33), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT25), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n476), .B1(new_n255), .B2(G107), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n374), .A2(KEYINPUT25), .A3(new_n435), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n475), .A2(G107), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(KEYINPUT90), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n264), .A2(new_n266), .A3(G257), .A4(G1698), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n264), .A2(new_n266), .A3(G250), .A4(new_n267), .ZN(new_n483));
  INV_X1    g0283(.A(G294), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n482), .B(new_n483), .C1(new_n263), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n355), .ZN(new_n486));
  INV_X1    g0286(.A(G45), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n487), .A2(G1), .ZN(new_n488));
  INV_X1    g0288(.A(G41), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n488), .B(KEYINPUT84), .C1(KEYINPUT5), .C2(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n214), .B(G45), .C1(new_n489), .C2(KEYINPUT5), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT84), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n489), .A2(KEYINPUT5), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n490), .A2(new_n493), .A3(new_n280), .A4(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n494), .ZN(new_n496));
  OAI211_X1 g0296(.A(G264), .B(new_n262), .C1(new_n496), .C2(new_n491), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n486), .A2(G179), .A3(new_n495), .A4(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n498), .A2(KEYINPUT91), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n498), .A2(KEYINPUT91), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n486), .A2(new_n495), .A3(new_n497), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G169), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n499), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT90), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n474), .A2(new_n504), .A3(new_n479), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n481), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n501), .A2(new_n289), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n501), .A2(G200), .ZN(new_n508));
  OR3_X1    g0308(.A1(new_n480), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n488), .A2(new_n279), .ZN(new_n510));
  INV_X1    g0310(.A(G250), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n487), .B2(G1), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n510), .A2(new_n262), .A3(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n264), .A2(new_n266), .A3(G238), .A4(new_n267), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(new_n263), .B2(new_n466), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n264), .A2(new_n266), .A3(G244), .A4(G1698), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT85), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT85), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n271), .A2(new_n520), .A3(G244), .A4(G1698), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n514), .B1(new_n523), .B2(new_n355), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(G190), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n516), .B1(new_n521), .B2(new_n519), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n513), .B1(new_n526), .B2(new_n262), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n424), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n475), .A2(G87), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT19), .ZN(new_n530));
  INV_X1    g0330(.A(G97), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n530), .B1(new_n380), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n271), .A2(new_n211), .A3(G68), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(KEYINPUT19), .B1(new_n350), .B2(new_n351), .ZN(new_n535));
  INV_X1    g0335(.A(G87), .ZN(new_n536));
  NOR2_X1   g0336(.A1(G97), .A2(G107), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n535), .A2(new_n211), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n251), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n442), .A2(new_n374), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n529), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n525), .A2(new_n528), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n475), .A2(new_n443), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n543), .A2(new_n539), .A3(new_n540), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT87), .ZN(new_n545));
  INV_X1    g0345(.A(G169), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n544), .A2(new_n545), .B1(new_n527), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT86), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n524), .A2(new_n548), .A3(new_n430), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n543), .A2(new_n539), .A3(KEYINPUT87), .A4(new_n540), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n430), .B(new_n513), .C1(new_n526), .C2(new_n262), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(KEYINPUT86), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n547), .A2(new_n549), .A3(new_n550), .A4(new_n552), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n506), .A2(new_n509), .A3(new_n542), .A4(new_n553), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n250), .A2(new_n210), .B1(G20), .B2(new_n466), .ZN(new_n555));
  AOI21_X1  g0355(.A(G20), .B1(G33), .B2(G283), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n263), .A2(G97), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT88), .ZN(new_n558));
  AND3_X1   g0358(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n558), .B1(new_n556), .B2(new_n557), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n555), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT20), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(KEYINPUT20), .B(new_n555), .C1(new_n559), .C2(new_n560), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n374), .A2(new_n466), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n214), .A2(G33), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n373), .A2(new_n375), .A3(G116), .A4(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n565), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(G270), .B(new_n262), .C1(new_n496), .C2(new_n491), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n495), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n271), .A2(G264), .A3(G1698), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n271), .A2(G257), .A3(new_n267), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n300), .A2(G303), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n355), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n546), .B1(new_n571), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n569), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT21), .ZN(new_n579));
  OAI21_X1  g0379(.A(KEYINPUT89), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT89), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n569), .A2(new_n577), .A3(new_n581), .A4(KEYINPUT21), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n571), .A2(new_n576), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n584), .A2(new_n430), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n578), .A2(new_n579), .B1(new_n585), .B2(new_n569), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n569), .B1(G200), .B2(new_n584), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(new_n289), .B2(new_n584), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n583), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT6), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n531), .A2(new_n435), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n590), .B1(new_n591), .B2(new_n537), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n435), .A2(KEYINPUT6), .A3(G97), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n594), .A2(G20), .B1(G77), .B2(new_n297), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n316), .A2(G107), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n252), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  XNOR2_X1  g0397(.A(new_n597), .B(KEYINPUT83), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n255), .A2(G97), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n475), .B2(G97), .ZN(new_n600));
  OAI211_X1 g0400(.A(G257), .B(new_n262), .C1(new_n496), .C2(new_n491), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n271), .A2(G244), .A3(new_n267), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT4), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n271), .A2(KEYINPUT4), .A3(G244), .A4(new_n267), .ZN(new_n606));
  NAND2_X1  g0406(.A1(G33), .A2(G283), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n271), .A2(G250), .A3(G1698), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n605), .A2(new_n606), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n602), .B1(new_n609), .B2(new_n355), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n610), .A2(G190), .A3(new_n495), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n495), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(G200), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n598), .A2(new_n600), .A3(new_n611), .A4(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n597), .A2(KEYINPUT83), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT83), .ZN(new_n616));
  AOI211_X1 g0416(.A(new_n616), .B(new_n252), .C1(new_n595), .C2(new_n596), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n600), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n610), .A2(new_n430), .A3(new_n495), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n612), .A2(new_n546), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n614), .A2(new_n621), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n554), .A2(new_n589), .A3(new_n622), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n459), .A2(new_n623), .ZN(G372));
  AOI21_X1  g0424(.A(KEYINPUT77), .B1(new_n395), .B2(new_n367), .ZN(new_n625));
  AND4_X1   g0425(.A1(KEYINPUT77), .A2(new_n367), .A3(new_n371), .A4(new_n390), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n404), .B1(new_n627), .B2(new_n457), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n345), .B1(KEYINPUT17), .B2(new_n332), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n343), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n429), .B(new_n428), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n632), .A2(new_n432), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n553), .A2(new_n542), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT26), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n634), .A2(new_n621), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n262), .B1(new_n517), .B2(new_n522), .ZN(new_n637));
  XNOR2_X1  g0437(.A(new_n513), .B(KEYINPUT92), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n424), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n525), .A2(new_n541), .A3(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n637), .A2(new_n638), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n544), .B(new_n551), .C1(new_n641), .C2(G169), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n635), .B1(new_n621), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n636), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n503), .A2(new_n480), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n583), .A2(new_n586), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n643), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n614), .A2(new_n650), .A3(new_n509), .A4(new_n621), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n642), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n459), .B1(new_n646), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n633), .A2(new_n653), .ZN(G369));
  NAND2_X1  g0454(.A1(new_n254), .A2(new_n211), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(new_n657), .A3(G213), .ZN(new_n658));
  INV_X1    g0458(.A(G343), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n506), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n481), .A2(KEYINPUT93), .A3(new_n505), .A4(new_n660), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n663), .A2(new_n506), .A3(new_n509), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n481), .A2(new_n505), .A3(new_n660), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT93), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n662), .B1(new_n664), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n569), .A2(new_n660), .ZN(new_n669));
  AND4_X1   g0469(.A1(new_n583), .A2(new_n586), .A3(new_n588), .A4(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n669), .B1(new_n583), .B2(new_n586), .ZN(new_n671));
  OAI21_X1  g0471(.A(G330), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(KEYINPUT94), .B1(new_n668), .B2(new_n672), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n480), .A2(new_n507), .A3(new_n508), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n474), .A2(new_n504), .A3(new_n479), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n504), .B1(new_n474), .B2(new_n479), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n674), .B1(new_n677), .B2(new_n503), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n678), .A2(new_n667), .A3(new_n663), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n506), .B2(new_n661), .ZN(new_n680));
  INV_X1    g0480(.A(G330), .ZN(new_n681));
  INV_X1    g0481(.A(new_n671), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n583), .A2(new_n586), .A3(new_n588), .A4(new_n669), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT94), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n680), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n673), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n503), .A2(new_n480), .A3(new_n661), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n660), .B1(new_n583), .B2(new_n586), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n689), .A2(new_n678), .A3(new_n667), .A4(new_n663), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n687), .A2(new_n688), .A3(new_n690), .ZN(G399));
  NAND2_X1  g0491(.A1(new_n217), .A2(new_n489), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT95), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n537), .A2(new_n536), .A3(new_n466), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n693), .A2(new_n214), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n695), .B1(new_n209), .B2(new_n693), .ZN(new_n696));
  XOR2_X1   g0496(.A(new_n696), .B(KEYINPUT28), .Z(new_n697));
  AND3_X1   g0497(.A1(new_n506), .A2(new_n583), .A3(new_n586), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n642), .B1(new_n698), .B2(new_n651), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n621), .A2(new_n635), .A3(new_n643), .ZN(new_n700));
  INV_X1    g0500(.A(new_n621), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n701), .A2(new_n542), .A3(new_n553), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n700), .B1(new_n702), .B2(new_n635), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n661), .B1(new_n699), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT29), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n589), .A2(new_n622), .ZN(new_n706));
  INV_X1    g0506(.A(new_n554), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(new_n707), .A3(new_n661), .ZN(new_n708));
  INV_X1    g0508(.A(new_n498), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n495), .A2(new_n570), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n710), .B1(new_n355), .B2(new_n575), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n709), .A2(new_n610), .A3(new_n524), .A4(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT30), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n527), .A2(new_n584), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n715), .A2(KEYINPUT30), .A3(new_n610), .A4(new_n709), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n711), .A2(G179), .ZN(new_n717));
  OR2_X1    g0517(.A1(new_n637), .A2(new_n638), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n717), .A2(new_n612), .A3(new_n718), .A4(new_n501), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n714), .A2(new_n716), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(new_n660), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT31), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT96), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n720), .A2(KEYINPUT31), .A3(new_n660), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n720), .A2(KEYINPUT31), .A3(new_n660), .ZN(new_n727));
  AOI21_X1  g0527(.A(KEYINPUT31), .B1(new_n720), .B2(new_n660), .ZN(new_n728));
  OAI21_X1  g0528(.A(KEYINPUT96), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n708), .A2(new_n726), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G330), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT29), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n732), .B(new_n661), .C1(new_n646), .C2(new_n652), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n705), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n697), .B1(new_n735), .B2(G1), .ZN(G364));
  NOR2_X1   g0536(.A1(G13), .A2(G33), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G20), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n682), .A2(new_n683), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n253), .A2(G20), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n214), .B1(new_n741), .B2(G45), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n693), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n217), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n300), .ZN(new_n746));
  NAND2_X1  g0546(.A1(G355), .A2(KEYINPUT97), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G355), .A2(KEYINPUT97), .ZN(new_n749));
  OAI22_X1  g0549(.A1(new_n748), .A2(new_n749), .B1(G116), .B2(new_n217), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n209), .A2(new_n487), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n745), .A2(new_n271), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n753), .B1(new_n245), .B2(G45), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n750), .B1(new_n751), .B2(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n210), .B1(G20), .B2(new_n546), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n739), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n744), .B1(new_n755), .B2(new_n758), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n759), .A2(KEYINPUT98), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G179), .A2(G200), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n211), .B1(new_n761), .B2(G190), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n531), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n211), .A2(new_n430), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G200), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n289), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n205), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT32), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n211), .A2(G190), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(new_n761), .ZN(new_n771));
  INV_X1    g0571(.A(G159), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n763), .B(new_n768), .C1(new_n769), .C2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n430), .A2(G200), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n770), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n271), .B1(new_n776), .B2(new_n381), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n764), .A2(new_n289), .A3(G200), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n773), .A2(new_n769), .B1(new_n294), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n775), .A2(G20), .A3(G190), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n777), .B(new_n779), .C1(G58), .C2(new_n781), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n424), .A2(G20), .A3(new_n430), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G190), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G107), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n783), .A2(new_n289), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G87), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n774), .A2(new_n782), .A3(new_n785), .A4(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n771), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n784), .A2(G283), .B1(G329), .B2(new_n789), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT100), .Z(new_n791));
  INV_X1    g0591(.A(G317), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n792), .A2(KEYINPUT33), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(KEYINPUT33), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n778), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(KEYINPUT99), .B(G326), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n767), .A2(new_n796), .B1(new_n484), .B2(new_n762), .ZN(new_n797));
  INV_X1    g0597(.A(G303), .ZN(new_n798));
  NOR3_X1   g0598(.A1(new_n783), .A2(new_n289), .A3(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G311), .ZN(new_n800));
  INV_X1    g0600(.A(G322), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n300), .B1(new_n776), .B2(new_n800), .C1(new_n801), .C2(new_n780), .ZN(new_n802));
  OR4_X1    g0602(.A1(new_n795), .A2(new_n797), .A3(new_n799), .A4(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n788), .B1(new_n791), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n760), .B1(new_n756), .B2(new_n804), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n740), .B(new_n805), .C1(KEYINPUT98), .C2(new_n759), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n682), .A2(new_n681), .A3(new_n683), .ZN(new_n807));
  INV_X1    g0607(.A(new_n744), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n672), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(G396));
  NAND2_X1  g0611(.A1(new_n455), .A2(new_n660), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n454), .A2(new_n457), .A3(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT102), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n454), .A2(new_n457), .A3(KEYINPUT102), .A4(new_n812), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n661), .B(new_n817), .C1(new_n646), .C2(new_n652), .ZN(new_n818));
  INV_X1    g0618(.A(new_n642), .ZN(new_n819));
  AND4_X1   g0619(.A1(new_n621), .A2(new_n650), .A3(new_n614), .A4(new_n509), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n819), .B1(new_n820), .B2(new_n648), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n644), .B1(new_n702), .B2(new_n635), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n660), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n457), .A2(new_n661), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n815), .A2(new_n824), .A3(new_n816), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n818), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n744), .B1(new_n826), .B2(new_n731), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n731), .B2(new_n826), .ZN(new_n828));
  INV_X1    g0628(.A(new_n756), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n738), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n744), .B1(G77), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n776), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n832), .A2(G116), .B1(new_n789), .B2(G311), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n833), .B(new_n300), .C1(new_n484), .C2(new_n780), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n763), .B(new_n834), .C1(G303), .C2(new_n766), .ZN(new_n835));
  AOI22_X1  g0635(.A1(G87), .A2(new_n784), .B1(new_n786), .B2(G107), .ZN(new_n836));
  INV_X1    g0636(.A(G283), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n778), .A2(KEYINPUT101), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n778), .A2(KEYINPUT101), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n835), .B(new_n836), .C1(new_n837), .C2(new_n840), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n781), .A2(G143), .B1(new_n832), .B2(G159), .ZN(new_n842));
  INV_X1    g0642(.A(G137), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n842), .B1(new_n411), .B2(new_n778), .C1(new_n843), .C2(new_n767), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT34), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n844), .A2(new_n845), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n784), .A2(G68), .ZN(new_n848));
  INV_X1    g0648(.A(G132), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n271), .B1(new_n762), .B2(new_n293), .C1(new_n849), .C2(new_n771), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(G50), .B2(new_n786), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n847), .A2(new_n848), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n841), .B1(new_n846), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n831), .B1(new_n853), .B2(new_n756), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n825), .B2(new_n738), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n828), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(G384));
  OR2_X1    g0657(.A1(new_n594), .A2(KEYINPUT35), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n594), .A2(KEYINPUT35), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n858), .A2(G116), .A3(new_n212), .A4(new_n859), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT36), .Z(new_n861));
  OAI211_X1 g0661(.A(new_n209), .B(G77), .C1(new_n293), .C2(new_n294), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(G50), .B2(new_n294), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n214), .A2(G13), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT38), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n321), .A2(new_n331), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n334), .B2(new_n338), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n334), .A2(new_n658), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n867), .A2(new_n871), .A3(KEYINPUT104), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n319), .B1(new_n334), .B2(new_n338), .ZN(new_n873));
  OAI21_X1  g0673(.A(KEYINPUT37), .B1(new_n873), .B2(new_n870), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT37), .B1(new_n341), .B2(new_n337), .ZN(new_n875));
  INV_X1    g0675(.A(new_n658), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n341), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n875), .A2(new_n321), .A3(new_n331), .A4(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT104), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n872), .A2(new_n874), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n877), .B1(new_n629), .B2(new_n343), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n866), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n312), .B1(new_n308), .B2(new_n310), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n328), .B(new_n251), .C1(new_n884), .C2(KEYINPUT16), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n658), .B1(new_n885), .B2(new_n258), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n347), .A2(new_n886), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n885), .A2(new_n258), .B1(new_n338), .B2(new_n658), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT37), .B1(new_n332), .B2(new_n888), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n889), .A2(KEYINPUT103), .A3(new_n878), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT103), .B1(new_n889), .B2(new_n878), .ZN(new_n891));
  OAI211_X1 g0691(.A(KEYINPUT38), .B(new_n887), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n883), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n825), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n389), .A2(new_n660), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n405), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n397), .A2(new_n404), .A3(new_n895), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n727), .A2(new_n728), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n708), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n893), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n887), .B1(new_n890), .B2(new_n891), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n866), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n892), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT105), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT40), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n899), .A2(new_n901), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT105), .B1(new_n899), .B2(new_n901), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI22_X1  g0713(.A1(new_n904), .A2(KEYINPUT40), .B1(new_n907), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n459), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n723), .A2(new_n725), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n623), .B2(new_n661), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n914), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n906), .A2(new_n892), .ZN(new_n919));
  INV_X1    g0719(.A(new_n898), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n895), .B1(new_n397), .B2(new_n404), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n825), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n908), .B1(new_n922), .B2(new_n917), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n899), .A2(new_n901), .A3(new_n910), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n902), .B1(new_n883), .B2(new_n892), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n919), .A2(new_n925), .B1(new_n909), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n927), .A2(new_n459), .A3(new_n901), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n918), .A2(new_n928), .A3(G330), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n929), .B(KEYINPUT106), .Z(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n457), .A2(new_n660), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n823), .B2(new_n817), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n897), .A2(new_n898), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n936), .A2(new_n907), .B1(new_n631), .B2(new_n658), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT39), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n893), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n906), .A2(KEYINPUT39), .A3(new_n892), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n404), .A2(new_n660), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n937), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n705), .A2(new_n733), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n459), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n633), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n943), .B(new_n946), .Z(new_n947));
  NOR2_X1   g0747(.A1(new_n931), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n947), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n930), .A2(new_n949), .B1(new_n214), .B2(new_n741), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n865), .B1(new_n948), .B2(new_n950), .ZN(G367));
  NOR2_X1   g0751(.A1(new_n541), .A2(new_n661), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n642), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n650), .B2(new_n952), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n954), .A2(KEYINPUT107), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(KEYINPUT107), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n739), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n762), .A2(new_n294), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n300), .B1(new_n789), .B2(G137), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n960), .B1(new_n205), .B2(new_n776), .C1(new_n411), .C2(new_n780), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n959), .B(new_n961), .C1(G143), .C2(new_n766), .ZN(new_n962));
  AOI22_X1  g0762(.A1(G58), .A2(new_n786), .B1(new_n784), .B2(G77), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n962), .B(new_n963), .C1(new_n772), .C2(new_n840), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n786), .A2(G116), .B1(KEYINPUT111), .B2(KEYINPUT46), .ZN(new_n965));
  NOR2_X1   g0765(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n965), .B(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n840), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(G294), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n780), .A2(new_n798), .B1(new_n776), .B2(new_n837), .ZN(new_n970));
  AOI211_X1 g0770(.A(new_n271), .B(new_n970), .C1(G317), .C2(new_n789), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n784), .A2(G97), .ZN(new_n972));
  INV_X1    g0772(.A(new_n762), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n766), .A2(G311), .B1(G107), .B2(new_n973), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n969), .A2(new_n971), .A3(new_n972), .A4(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n964), .B1(new_n967), .B2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT47), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n756), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n234), .A2(new_n753), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n758), .B1(new_n745), .B2(new_n443), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n808), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AND3_X1   g0782(.A1(new_n958), .A2(new_n978), .A3(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n689), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n679), .B(new_n985), .C1(new_n506), .C2(new_n661), .ZN(new_n986));
  AND3_X1   g0786(.A1(new_n986), .A2(new_n672), .A3(new_n690), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n672), .B1(new_n986), .B2(new_n690), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n734), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n618), .A2(new_n660), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n614), .A2(new_n621), .A3(new_n991), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n618), .A2(new_n619), .A3(new_n620), .A4(new_n660), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n690), .A2(new_n688), .A3(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT45), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n690), .A2(KEYINPUT45), .A3(new_n688), .A4(new_n994), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n690), .A2(new_n688), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n992), .A2(new_n993), .ZN(new_n1001));
  AOI21_X1  g0801(.A(KEYINPUT44), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  AND3_X1   g0802(.A1(new_n1000), .A2(KEYINPUT44), .A3(new_n1001), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n999), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AND2_X1   g0804(.A1(new_n673), .A2(new_n686), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n687), .B(new_n999), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n990), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n735), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n693), .B(KEYINPUT41), .Z(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n743), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n1013));
  NAND2_X1  g0813(.A1(new_n957), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT109), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n690), .B2(new_n1001), .ZN(new_n1016));
  AND3_X1   g0816(.A1(new_n678), .A2(new_n667), .A3(new_n663), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1017), .A2(KEYINPUT109), .A3(new_n689), .A4(new_n994), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(KEYINPUT42), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT42), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1016), .A2(new_n1018), .A3(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n621), .B1(new_n992), .B2(new_n506), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n661), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1020), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1005), .A2(new_n994), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n955), .A2(KEYINPUT43), .A3(new_n956), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT110), .ZN(new_n1028));
  AND3_X1   g0828(.A1(new_n1025), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1026), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1014), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1026), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1014), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1025), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1031), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n984), .B1(new_n1012), .B2(new_n1038), .ZN(G387));
  INV_X1    g0839(.A(new_n989), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n735), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n734), .A2(new_n989), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1041), .A2(new_n693), .A3(new_n1042), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n746), .A2(new_n694), .B1(new_n435), .B2(new_n745), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n238), .A2(new_n487), .ZN(new_n1045));
  AOI211_X1 g0845(.A(G45), .B(new_n694), .C1(G68), .C2(G77), .ZN(new_n1046));
  AOI21_X1  g0846(.A(KEYINPUT50), .B1(new_n247), .B2(new_n205), .ZN(new_n1047));
  AND3_X1   g0847(.A1(new_n247), .A2(KEYINPUT50), .A3(new_n205), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1046), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n752), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1044), .B1(new_n1045), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n808), .B1(new_n1051), .B2(new_n757), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n762), .A2(new_n442), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n778), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1053), .B1(new_n1054), .B2(new_n247), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n772), .B2(new_n767), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n300), .B1(new_n789), .B2(G150), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n781), .A2(G50), .B1(new_n832), .B2(G68), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n972), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1056), .B(new_n1059), .C1(G77), .C2(new_n786), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n300), .B1(new_n771), .B2(new_n796), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n781), .A2(G317), .B1(new_n832), .B2(G303), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(new_n801), .B2(new_n767), .C1(new_n840), .C2(new_n800), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT48), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n786), .A2(G294), .B1(G283), .B2(new_n973), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT49), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1061), .B(new_n1070), .C1(G116), .C2(new_n784), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1060), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1052), .B1(new_n1073), .B2(new_n829), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n668), .B2(new_n739), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n1040), .B2(new_n743), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1043), .A2(new_n1076), .ZN(G393));
  INV_X1    g0877(.A(KEYINPUT112), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1006), .A2(new_n1078), .A3(new_n1007), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n1007), .A2(new_n1078), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1079), .A2(new_n1080), .A3(new_n1041), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1081), .A2(new_n693), .A3(new_n1008), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n300), .B1(new_n832), .B2(new_n247), .ZN(new_n1083));
  INV_X1    g0883(.A(G143), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1083), .B1(new_n1084), .B2(new_n771), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(G77), .B2(new_n973), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(G68), .A2(new_n786), .B1(new_n784), .B2(G87), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1086), .B(new_n1087), .C1(new_n205), .C2(new_n840), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n766), .A2(G150), .B1(new_n781), .B2(G159), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT51), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n300), .B1(new_n771), .B2(new_n801), .C1(new_n484), .C2(new_n776), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(G116), .B2(new_n973), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G107), .A2(new_n784), .B1(new_n786), .B2(G283), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1092), .B(new_n1093), .C1(new_n798), .C2(new_n840), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n766), .A2(G317), .B1(new_n781), .B2(G311), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT52), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n1088), .A2(new_n1090), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n756), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n752), .A2(new_n242), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1099), .B(new_n757), .C1(new_n531), .C2(new_n217), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1098), .A2(new_n744), .A3(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n1001), .B2(new_n739), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1102), .B1(new_n1103), .B2(new_n743), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1082), .A2(new_n1104), .ZN(G390));
  INV_X1    g0905(.A(KEYINPUT116), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT114), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n917), .A2(new_n681), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n899), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n932), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n818), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n941), .B1(new_n1111), .B2(new_n934), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n906), .A2(KEYINPUT39), .A3(new_n892), .ZN(new_n1114));
  AOI21_X1  g0914(.A(KEYINPUT39), .B1(new_n883), .B2(new_n892), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n941), .B(KEYINPUT113), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n661), .B(new_n817), .C1(new_n699), .C2(new_n703), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n1110), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1117), .B1(new_n1119), .B2(new_n934), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n893), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1109), .B1(new_n1116), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1112), .B1(new_n939), .B2(new_n940), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n1120), .A2(new_n893), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n730), .A2(new_n934), .A3(G330), .A4(new_n825), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n1123), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1107), .B1(new_n1122), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n901), .A2(G330), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n935), .B1(new_n1129), .B2(new_n894), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1130), .A2(new_n1110), .A3(new_n1125), .A4(new_n1118), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n730), .A2(G330), .A3(new_n825), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n935), .A2(new_n1132), .B1(new_n1108), .B2(new_n899), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1131), .B1(new_n933), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1108), .A2(new_n459), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n945), .A2(new_n633), .A3(new_n1135), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n1134), .A2(new_n1136), .A3(KEYINPUT115), .ZN(new_n1137));
  AOI21_X1  g0937(.A(KEYINPUT115), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1116), .A2(new_n1125), .A3(new_n1121), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1109), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1140), .A2(new_n1142), .A3(KEYINPUT114), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1128), .A2(new_n1139), .A3(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n945), .A2(new_n633), .A3(new_n1135), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n1132), .A2(new_n935), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1111), .B1(new_n1141), .B2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1145), .B1(new_n1147), .B2(new_n1131), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1140), .A2(new_n1142), .A3(new_n1148), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n1149), .A2(new_n693), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1106), .B1(new_n1144), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1140), .A2(new_n1142), .A3(new_n743), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n737), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n744), .B1(new_n247), .B2(new_n830), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n780), .A2(new_n466), .B1(new_n762), .B2(new_n381), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT117), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n300), .B1(new_n771), .B2(new_n484), .C1(new_n531), .C2(new_n776), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(G283), .B2(new_n766), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1159), .A2(new_n787), .A3(new_n848), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1157), .B(new_n1160), .C1(G107), .C2(new_n968), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  OR2_X1    g0962(.A1(new_n1162), .A2(KEYINPUT118), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(KEYINPUT118), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n786), .A2(G150), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n968), .A2(G137), .B1(new_n1165), .B2(KEYINPUT53), .ZN(new_n1166));
  OR2_X1    g0966(.A1(new_n1165), .A2(KEYINPUT53), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n784), .A2(G50), .ZN(new_n1168));
  INV_X1    g0968(.A(G128), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n767), .A2(new_n1169), .B1(new_n762), .B2(new_n772), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(KEYINPUT54), .B(G143), .ZN(new_n1171));
  INV_X1    g0971(.A(G125), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n776), .A2(new_n1171), .B1(new_n771), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n271), .B1(new_n780), .B2(new_n849), .ZN(new_n1174));
  NOR3_X1   g0974(.A1(new_n1170), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .A4(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1163), .A2(new_n1164), .A3(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1155), .B1(new_n1177), .B2(new_n756), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1154), .A2(new_n1178), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n1153), .A2(KEYINPUT119), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(KEYINPUT119), .B1(new_n1153), .B2(new_n1179), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1144), .A2(new_n1150), .A3(new_n1106), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1152), .A2(new_n1183), .A3(new_n1184), .ZN(G378));
  INV_X1    g0985(.A(new_n943), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n414), .A2(new_n876), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT120), .Z(new_n1188));
  XNOR2_X1  g0988(.A(new_n433), .B(new_n1188), .ZN(new_n1189));
  XOR2_X1   g0989(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1190));
  XNOR2_X1  g0990(.A(new_n1189), .B(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n925), .B1(new_n892), .B2(new_n906), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n926), .A2(new_n909), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1192), .B(G330), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1192), .B1(new_n927), .B2(G330), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1186), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1191), .B1(new_n914), .B2(new_n681), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1199), .A2(new_n943), .A3(new_n1195), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1198), .A2(new_n743), .A3(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n744), .B1(G50), .B2(new_n830), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n205), .B1(G33), .B2(G41), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n300), .B2(new_n489), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n489), .B(new_n300), .C1(new_n771), .C2(new_n837), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n780), .A2(new_n435), .B1(new_n776), .B2(new_n442), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1205), .B(new_n1206), .C1(new_n786), .C2(G77), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n778), .A2(new_n531), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n959), .B(new_n1208), .C1(G116), .C2(new_n766), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n784), .A2(G58), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1207), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT58), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1204), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1171), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n786), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1054), .A2(G132), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n781), .A2(G128), .B1(new_n832), .B2(G137), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n766), .A2(G125), .B1(G150), .B2(new_n973), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(KEYINPUT59), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n784), .A2(G159), .ZN(new_n1221));
  AOI211_X1 g1021(.A(G33), .B(G41), .C1(new_n789), .C2(G124), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1219), .A2(KEYINPUT59), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1213), .B1(new_n1212), .B2(new_n1211), .C1(new_n1223), .C2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1202), .B1(new_n1225), .B2(new_n756), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n1191), .B2(new_n738), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1201), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1149), .A2(new_n1136), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1230), .A2(KEYINPUT57), .A3(new_n1200), .A4(new_n1198), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n693), .ZN(new_n1232));
  AND3_X1   g1032(.A1(new_n1199), .A2(new_n943), .A3(new_n1195), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n943), .B1(new_n1199), .B2(new_n1195), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT57), .B1(new_n1235), .B2(new_n1230), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1229), .B1(new_n1232), .B2(new_n1236), .ZN(G375));
  OAI211_X1 g1037(.A(new_n1139), .B(new_n1011), .C1(new_n1136), .C2(new_n1134), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n935), .A2(new_n737), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n744), .B1(G68), .B2(new_n830), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT121), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n271), .B1(new_n789), .B2(G303), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n1242), .B1(new_n435), .B2(new_n776), .C1(new_n837), .C2(new_n780), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n1053), .B(new_n1243), .C1(G294), .C2(new_n766), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(G77), .A2(new_n784), .B1(new_n786), .B2(G97), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1244), .B(new_n1245), .C1(new_n466), .C2(new_n840), .ZN(new_n1246));
  OR3_X1    g1046(.A1(new_n767), .A2(KEYINPUT122), .A3(new_n849), .ZN(new_n1247));
  OAI21_X1  g1047(.A(KEYINPUT122), .B1(new_n767), .B2(new_n849), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n1247), .A2(new_n1248), .B1(new_n968), .B2(new_n1214), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n271), .B1(new_n771), .B2(new_n1169), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n780), .A2(new_n843), .B1(new_n776), .B2(new_n411), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n1250), .B(new_n1251), .C1(G50), .C2(new_n973), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n786), .A2(G159), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1249), .A2(new_n1210), .A3(new_n1252), .A4(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1246), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1241), .B1(new_n1255), .B2(new_n756), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1134), .A2(new_n743), .B1(new_n1239), .B2(new_n1256), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1238), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(G381));
  NAND2_X1  g1059(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n742), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1031), .A2(new_n1037), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n983), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  NOR4_X1   g1063(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1258), .A2(new_n1263), .A3(new_n1264), .ZN(new_n1265));
  XOR2_X1   g1065(.A(new_n1265), .B(KEYINPUT123), .Z(new_n1266));
  AND2_X1   g1066(.A1(new_n1231), .A2(new_n693), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1235), .A2(new_n1230), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT57), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1228), .B1(new_n1267), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1153), .A2(new_n1179), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(new_n1144), .B2(new_n1150), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1266), .A2(new_n1271), .A3(new_n1273), .ZN(G407));
  NAND2_X1  g1074(.A1(new_n659), .A2(G213), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1271), .A2(new_n1273), .A3(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(G407), .A2(G213), .A3(new_n1277), .ZN(G409));
  NOR2_X1   g1078(.A1(G393), .A2(G396), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n810), .B1(new_n1043), .B2(new_n1076), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1263), .A2(G390), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1082), .A2(new_n1104), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(G387), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1282), .B1(new_n1283), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT125), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1010), .B1(new_n1008), .B2(new_n735), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1037), .B(new_n1031), .C1(new_n1288), .C2(new_n743), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT124), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(G390), .A2(new_n1289), .A3(new_n1290), .A4(new_n984), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1285), .A2(new_n1291), .A3(new_n1282), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1290), .B1(new_n1263), .B2(G390), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1287), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1281), .B1(G387), .B2(new_n1284), .ZN(new_n1295));
  OAI21_X1  g1095(.A(KEYINPUT124), .B1(G387), .B2(new_n1284), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1295), .A2(new_n1296), .A3(KEYINPUT125), .A4(new_n1291), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1286), .B1(new_n1294), .B2(new_n1297), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1299), .A2(KEYINPUT60), .A3(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n693), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1299), .B1(KEYINPUT60), .B2(new_n1300), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1257), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n856), .ZN(new_n1305));
  OAI211_X1 g1105(.A(G384), .B(new_n1257), .C1(new_n1302), .C2(new_n1303), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1276), .A2(G2897), .ZN(new_n1308));
  XNOR2_X1  g1108(.A(new_n1307), .B(new_n1308), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1230), .A2(new_n1011), .A3(new_n1200), .A4(new_n1198), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1310), .A2(new_n1201), .A3(new_n1227), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1311), .A2(new_n1273), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1312), .B1(new_n1271), .B2(G378), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1309), .B1(new_n1313), .B2(new_n1276), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT61), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1311), .A2(new_n1273), .ZN(new_n1316));
  AND3_X1   g1116(.A1(new_n1144), .A2(new_n1106), .A3(new_n1150), .ZN(new_n1317));
  NOR3_X1   g1117(.A1(new_n1317), .A2(new_n1151), .A3(new_n1182), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1316), .B1(new_n1318), .B2(G375), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT62), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1307), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1319), .A2(new_n1320), .A3(new_n1275), .A4(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1314), .A2(new_n1315), .A3(new_n1322), .ZN(new_n1323));
  XOR2_X1   g1123(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1324));
  NAND2_X1  g1124(.A1(new_n1271), .A2(G378), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1276), .B1(new_n1325), .B2(new_n1316), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1324), .B1(new_n1326), .B2(new_n1321), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1298), .B1(new_n1323), .B2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT63), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1319), .A2(new_n1275), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1329), .B1(new_n1330), .B2(new_n1307), .ZN(new_n1331));
  AOI21_X1  g1131(.A(KEYINPUT61), .B1(new_n1330), .B2(new_n1309), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1326), .A2(KEYINPUT63), .A3(new_n1321), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1294), .A2(new_n1297), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1286), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  NAND4_X1  g1136(.A1(new_n1331), .A2(new_n1332), .A3(new_n1333), .A4(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1328), .A2(new_n1337), .ZN(G405));
  INV_X1    g1138(.A(KEYINPUT127), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1336), .A2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1298), .A2(KEYINPUT127), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1340), .A2(new_n1307), .A3(new_n1341), .ZN(new_n1342));
  AOI21_X1  g1142(.A(KEYINPUT127), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1343));
  AOI211_X1 g1143(.A(new_n1339), .B(new_n1286), .C1(new_n1294), .C2(new_n1297), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1321), .B1(new_n1343), .B2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(G375), .A2(new_n1273), .ZN(new_n1346));
  AND2_X1   g1146(.A1(new_n1325), .A2(new_n1346), .ZN(new_n1347));
  AND3_X1   g1147(.A1(new_n1342), .A2(new_n1345), .A3(new_n1347), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1347), .B1(new_n1342), .B2(new_n1345), .ZN(new_n1349));
  NOR2_X1   g1149(.A1(new_n1348), .A2(new_n1349), .ZN(G402));
endmodule


