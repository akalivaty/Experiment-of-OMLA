//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 1 1 1 1 0 1 0 0 1 0 0 0 1 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT2), .B(G113), .Z(new_n188));
  XNOR2_X1  g002(.A(G116), .B(G119), .ZN(new_n189));
  AND2_X1   g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n188), .A2(new_n189), .ZN(new_n191));
  OR2_X1    g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT64), .ZN(new_n193));
  XNOR2_X1  g007(.A(G143), .B(G146), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT0), .B(G128), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n193), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G143), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT0), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT0), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G128), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n201), .A2(new_n206), .A3(KEYINPUT64), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n194), .A2(KEYINPUT0), .A3(G128), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n196), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G134), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT11), .B1(new_n211), .B2(G137), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT11), .ZN(new_n213));
  INV_X1    g027(.A(G137), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(G134), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n217), .B1(new_n214), .B2(G134), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n211), .A2(KEYINPUT66), .A3(G137), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n216), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G131), .ZN(new_n222));
  INV_X1    g036(.A(G131), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n216), .A2(new_n220), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n226));
  OR2_X1    g040(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n200), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(G128), .B1(new_n198), .B2(new_n200), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n226), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n197), .A2(G143), .ZN(new_n232));
  AND2_X1   g046(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n233));
  NOR2_X1   g047(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n235), .B(KEYINPUT68), .C1(G128), .C2(new_n194), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n194), .A2(G128), .A3(new_n227), .A4(new_n228), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n231), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n211), .A2(G137), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n214), .A2(G134), .ZN(new_n240));
  OAI21_X1  g054(.A(G131), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n224), .A2(new_n241), .ZN(new_n242));
  AOI22_X1  g056(.A1(new_n210), .A2(new_n225), .B1(new_n238), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT30), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n224), .A2(new_n241), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n198), .A2(new_n200), .A3(G128), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n227), .A2(new_n228), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n235), .B1(G128), .B2(new_n194), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n248), .B1(new_n249), .B2(new_n226), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n245), .B1(new_n250), .B2(new_n236), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT65), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n196), .A2(new_n207), .A3(new_n252), .A4(new_n208), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n225), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n209), .A2(KEYINPUT65), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n251), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n192), .B(new_n244), .C1(new_n256), .C2(KEYINPUT30), .ZN(new_n257));
  INV_X1    g071(.A(new_n192), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n243), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(G237), .A2(G953), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G210), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT27), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n261), .B(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n263), .B(KEYINPUT26), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G101), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT26), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n263), .B(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G101), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n257), .A2(new_n259), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT31), .ZN(new_n273));
  OR2_X1    g087(.A1(new_n256), .A2(new_n258), .ZN(new_n274));
  AOI21_X1  g088(.A(KEYINPUT28), .B1(new_n243), .B2(new_n258), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n238), .A2(new_n242), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n201), .A2(new_n206), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n198), .A2(new_n200), .A3(G128), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n277), .A2(new_n193), .B1(new_n278), .B2(KEYINPUT0), .ZN(new_n279));
  INV_X1    g093(.A(new_n224), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n223), .B1(new_n216), .B2(new_n220), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n279), .B(new_n207), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  AND4_X1   g096(.A1(KEYINPUT28), .A2(new_n276), .A3(new_n282), .A4(new_n258), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n275), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n274), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n270), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n273), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n259), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n255), .A2(new_n253), .A3(new_n225), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT30), .B1(new_n289), .B2(new_n276), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n276), .A2(new_n282), .A3(KEYINPUT30), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n288), .B1(new_n292), .B2(new_n192), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT70), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT69), .B(KEYINPUT31), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n293), .A2(new_n294), .A3(new_n295), .A4(new_n271), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n257), .A2(new_n295), .A3(new_n259), .A4(new_n271), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT70), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n287), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(G472), .A2(G902), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  OAI211_X1 g115(.A(KEYINPUT71), .B(new_n187), .C1(new_n299), .C2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT71), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n296), .A2(new_n298), .ZN(new_n304));
  AOI22_X1  g118(.A1(new_n272), .A2(KEYINPUT31), .B1(new_n285), .B2(new_n270), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n301), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n303), .B1(new_n306), .B2(KEYINPUT32), .ZN(new_n307));
  INV_X1    g121(.A(G472), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT29), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n270), .B1(new_n274), .B2(new_n284), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n270), .A2(new_n259), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n311), .B1(new_n292), .B2(new_n192), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n309), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  OR2_X1    g127(.A1(new_n243), .A2(new_n258), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n284), .A2(KEYINPUT29), .A3(new_n271), .A4(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G902), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n308), .B1(new_n313), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n318), .B1(new_n306), .B2(KEYINPUT32), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n302), .A2(new_n307), .A3(new_n319), .ZN(new_n320));
  XOR2_X1   g134(.A(KEYINPUT72), .B(G217), .Z(new_n321));
  AOI21_X1  g135(.A(new_n321), .B1(G234), .B2(new_n316), .ZN(new_n322));
  INV_X1    g136(.A(G140), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G125), .ZN(new_n324));
  INV_X1    g138(.A(G125), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G140), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(new_n326), .A3(KEYINPUT16), .ZN(new_n327));
  OR3_X1    g141(.A1(new_n325), .A2(KEYINPUT16), .A3(G140), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(new_n328), .A3(G146), .ZN(new_n329));
  XNOR2_X1  g143(.A(G125), .B(G140), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n197), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G119), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT74), .B1(new_n333), .B2(G128), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT23), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(G128), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT23), .ZN(new_n337));
  OAI211_X1 g151(.A(KEYINPUT74), .B(new_n337), .C1(new_n333), .C2(G128), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n335), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G110), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT73), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n342), .B1(new_n333), .B2(G128), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n202), .A2(KEYINPUT73), .A3(G119), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n336), .A3(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT24), .B(G110), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI22_X1  g161(.A1(new_n340), .A2(new_n341), .B1(new_n347), .B2(KEYINPUT75), .ZN(new_n348));
  OR2_X1    g162(.A1(new_n347), .A2(KEYINPUT75), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n332), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OAI22_X1  g164(.A1(new_n340), .A2(new_n341), .B1(new_n346), .B2(new_n345), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n327), .A2(new_n328), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n197), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n353), .A2(new_n329), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n350), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G953), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n357), .A2(G221), .A3(G234), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n358), .B(KEYINPUT22), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n359), .B(G137), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n360), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n362), .B1(new_n350), .B2(new_n355), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(new_n363), .A3(new_n316), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT25), .ZN(new_n365));
  AND3_X1   g179(.A1(new_n364), .A2(KEYINPUT76), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n365), .B1(new_n364), .B2(KEYINPUT76), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n322), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n322), .A2(G902), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n361), .A2(new_n363), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT84), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT3), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(KEYINPUT78), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT78), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT3), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G107), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G104), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G104), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n382), .A2(G107), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n379), .A2(G104), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n377), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(KEYINPUT80), .B(G101), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n381), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n382), .A2(G107), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n380), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G101), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n189), .A2(KEYINPUT5), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT5), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(new_n333), .A3(G116), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G113), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n190), .B1(new_n392), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n391), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n387), .A2(KEYINPUT4), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n381), .A2(new_n385), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT79), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n268), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n381), .A2(new_n385), .A3(KEYINPUT79), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n399), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n383), .B1(new_n375), .B2(new_n377), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n380), .A2(new_n388), .B1(new_n376), .B2(KEYINPUT3), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n401), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT4), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n407), .A2(new_n403), .A3(new_n408), .A4(G101), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n192), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n398), .B1(new_n404), .B2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(G110), .B(G122), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n412), .B(new_n398), .C1(new_n404), .C2(new_n410), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(KEYINPUT6), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n209), .A2(G125), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n417), .B1(new_n238), .B2(G125), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n357), .A2(G224), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(KEYINPUT82), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n418), .B(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT6), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n411), .A2(new_n422), .A3(new_n413), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n416), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT7), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n418), .B1(new_n425), .B2(new_n420), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n420), .A2(new_n425), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n417), .B(new_n427), .C1(new_n238), .C2(G125), .ZN(new_n428));
  OR2_X1    g242(.A1(new_n395), .A2(KEYINPUT83), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n395), .A2(KEYINPUT83), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n429), .A2(new_n392), .A3(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n391), .B1(new_n431), .B2(new_n190), .ZN(new_n432));
  XOR2_X1   g246(.A(new_n412), .B(KEYINPUT8), .Z(new_n433));
  NAND2_X1  g247(.A1(new_n387), .A2(new_n390), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n433), .B1(new_n397), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n426), .A2(new_n428), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(G902), .B1(new_n437), .B2(new_n415), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n424), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(G210), .B1(G237), .B2(G902), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n424), .A2(new_n440), .A3(new_n438), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(G214), .B1(G237), .B2(G902), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n373), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n424), .A2(new_n440), .A3(new_n438), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n440), .B1(new_n424), .B2(new_n438), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n373), .B(new_n445), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G469), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n407), .A2(new_n403), .A3(G101), .ZN(new_n453));
  AOI22_X1  g267(.A1(new_n380), .A2(new_n378), .B1(new_n389), .B2(new_n377), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n408), .B1(new_n454), .B2(new_n386), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n456), .A2(new_n210), .A3(new_n409), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n387), .A2(KEYINPUT10), .A3(new_n390), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n201), .A2(new_n202), .B1(KEYINPUT1), .B2(new_n232), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n237), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(new_n387), .A3(new_n390), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT10), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n238), .A2(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n225), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n457), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n461), .B1(new_n391), .B2(new_n238), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n466), .A2(KEYINPUT12), .A3(new_n225), .ZN(new_n467));
  AOI21_X1  g281(.A(KEYINPUT12), .B1(new_n466), .B2(new_n225), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(G110), .B(G140), .ZN(new_n470));
  INV_X1    g284(.A(G227), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n471), .A2(G953), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n470), .B(new_n472), .ZN(new_n473));
  XOR2_X1   g287(.A(new_n473), .B(KEYINPUT77), .Z(new_n474));
  NAND2_X1  g288(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n456), .A2(new_n210), .A3(new_n409), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n458), .A2(new_n238), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n461), .A2(new_n462), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n225), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n473), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(new_n465), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n475), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n452), .B1(new_n483), .B2(new_n316), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n465), .B(new_n481), .C1(new_n467), .C2(new_n468), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n481), .B1(new_n480), .B2(new_n465), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n452), .B(new_n316), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT81), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n465), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n464), .B1(new_n457), .B2(new_n463), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n473), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(G902), .B1(new_n493), .B2(new_n485), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(KEYINPUT81), .A3(new_n452), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n484), .B1(new_n490), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G122), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(G113), .ZN(new_n498));
  INV_X1    g312(.A(G113), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(G122), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n498), .A2(new_n500), .A3(G104), .ZN(new_n501));
  AOI21_X1  g315(.A(G104), .B1(new_n498), .B2(new_n500), .ZN(new_n502));
  NOR3_X1   g316(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT86), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT86), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n498), .A2(new_n500), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n382), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n498), .A2(new_n500), .A3(G104), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n504), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n330), .B(new_n197), .ZN(new_n510));
  INV_X1    g324(.A(G237), .ZN(new_n511));
  AND4_X1   g325(.A1(G143), .A2(new_n511), .A3(new_n357), .A4(G214), .ZN(new_n512));
  AOI21_X1  g326(.A(G143), .B1(new_n260), .B2(G214), .ZN(new_n513));
  OAI211_X1 g327(.A(KEYINPUT18), .B(G131), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n511), .A2(new_n357), .A3(G214), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n199), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n260), .A2(G143), .A3(G214), .ZN(new_n517));
  NAND2_X1  g331(.A1(KEYINPUT18), .A2(G131), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n510), .A2(new_n514), .A3(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(G131), .B1(new_n512), .B2(new_n513), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT17), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n516), .A2(new_n223), .A3(new_n517), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  OAI211_X1 g338(.A(KEYINPUT17), .B(G131), .C1(new_n512), .C2(new_n513), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n353), .A2(new_n329), .A3(new_n525), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n509), .B(new_n520), .C1(new_n524), .C2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n524), .A2(new_n526), .ZN(new_n528));
  INV_X1    g342(.A(new_n520), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n501), .A2(new_n502), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n527), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n316), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(G475), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NOR3_X1   g349(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT85), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT19), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n325), .A2(G140), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n323), .A2(G125), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n324), .A2(new_n326), .A3(KEYINPUT19), .ZN(new_n542));
  AOI21_X1  g356(.A(G146), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n327), .A2(G146), .A3(new_n328), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n537), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n521), .A2(new_n523), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n324), .A2(new_n326), .A3(KEYINPUT19), .ZN(new_n547));
  AOI21_X1  g361(.A(KEYINPUT19), .B1(new_n324), .B2(new_n326), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n197), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n549), .A2(KEYINPUT85), .A3(new_n329), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n545), .A2(new_n546), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n531), .B1(new_n551), .B2(new_n520), .ZN(new_n552));
  INV_X1    g366(.A(new_n527), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n536), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT88), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g370(.A(KEYINPUT88), .B(new_n536), .C1(new_n552), .C2(new_n553), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n550), .A2(new_n546), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n529), .B1(new_n559), .B2(new_n545), .ZN(new_n560));
  OAI211_X1 g374(.A(KEYINPUT87), .B(new_n527), .C1(new_n560), .C2(new_n531), .ZN(new_n561));
  NOR2_X1   g375(.A1(G475), .A2(G902), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT87), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n563), .B1(new_n552), .B2(new_n553), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT20), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n535), .B1(new_n558), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(G234), .A2(G237), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n568), .A2(G952), .A3(new_n357), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT21), .B(G898), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n568), .A2(G902), .A3(G953), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n569), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(G128), .B(G143), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT13), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n199), .A2(G128), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n575), .B(G134), .C1(KEYINPUT13), .C2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(G116), .B(G122), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(new_n379), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n574), .A2(new_n211), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT14), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  OR2_X1    g397(.A1(new_n497), .A2(G116), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n583), .B(G107), .C1(new_n582), .C2(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n574), .B(new_n211), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n578), .A2(new_n379), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n581), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT9), .B(G234), .ZN(new_n590));
  NOR3_X1   g404(.A1(new_n321), .A2(G953), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT89), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n581), .A2(new_n588), .A3(new_n591), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n589), .A2(KEYINPUT89), .A3(new_n592), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(new_n316), .A3(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(G478), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n599), .A2(KEYINPUT15), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n598), .B(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n567), .A2(new_n573), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(G221), .B1(new_n590), .B2(G902), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n496), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n320), .A2(new_n372), .A3(new_n451), .A4(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(KEYINPUT90), .ZN(new_n608));
  XOR2_X1   g422(.A(new_n608), .B(new_n386), .Z(G3));
  NOR3_X1   g423(.A1(new_n496), .A2(new_n371), .A3(new_n605), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n304), .A2(new_n305), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n308), .B1(new_n611), .B2(new_n316), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(new_n306), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n445), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n615), .B1(new_n442), .B2(new_n443), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n573), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n558), .A2(new_n566), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n534), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n598), .A2(new_n599), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n589), .A2(KEYINPUT91), .A3(new_n592), .ZN(new_n621));
  AOI21_X1  g435(.A(KEYINPUT91), .B1(new_n589), .B2(new_n592), .ZN(new_n622));
  OAI211_X1 g436(.A(KEYINPUT33), .B(new_n595), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT33), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n596), .A2(new_n624), .A3(new_n597), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n316), .A2(G478), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n620), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n619), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n617), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n614), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT34), .B(G104), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G6));
  XNOR2_X1  g447(.A(new_n565), .B(KEYINPUT20), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n634), .A2(new_n534), .A3(new_n601), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n617), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n614), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(new_n637), .B(KEYINPUT92), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT35), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G107), .ZN(G9));
  INV_X1    g454(.A(KEYINPUT93), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n356), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(KEYINPUT93), .B1(new_n350), .B2(new_n355), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n644), .B1(KEYINPUT36), .B2(new_n362), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n362), .A2(KEYINPUT36), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n642), .A2(new_n646), .A3(new_n643), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n645), .A2(new_n369), .A3(new_n647), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n368), .A2(new_n648), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n612), .A2(new_n306), .A3(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n650), .A2(new_n451), .A3(new_n606), .ZN(new_n651));
  XOR2_X1   g465(.A(new_n651), .B(KEYINPUT37), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT94), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G110), .ZN(G12));
  INV_X1    g468(.A(new_n484), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n488), .A2(new_n489), .ZN(new_n656));
  AOI21_X1  g470(.A(KEYINPUT81), .B1(new_n494), .B2(new_n452), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n604), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n368), .A2(new_n648), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n616), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n569), .B1(new_n572), .B2(G900), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n634), .A2(new_n534), .A3(new_n601), .A4(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n662), .A2(new_n320), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G128), .ZN(G30));
  NOR2_X1   g481(.A1(new_n496), .A2(new_n605), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n663), .B(KEYINPUT95), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT39), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n671), .B(KEYINPUT96), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(KEYINPUT40), .ZN(new_n673));
  INV_X1    g487(.A(new_n293), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n271), .ZN(new_n675));
  INV_X1    g489(.A(new_n311), .ZN(new_n676));
  AOI21_X1  g490(.A(G902), .B1(new_n676), .B2(new_n314), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n308), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n678), .B1(new_n306), .B2(KEYINPUT32), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n302), .A2(new_n307), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n681), .A2(new_n660), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT38), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n444), .B(new_n683), .ZN(new_n684));
  NOR4_X1   g498(.A1(new_n684), .A2(new_n615), .A3(new_n567), .A4(new_n602), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n673), .A2(new_n682), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G143), .ZN(G45));
  AND2_X1   g501(.A1(new_n619), .A2(new_n628), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n688), .A2(new_n663), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n662), .A2(new_n320), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT97), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G146), .ZN(G48));
  OAI21_X1  g506(.A(new_n316), .B1(new_n486), .B2(new_n487), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT98), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n494), .A2(KEYINPUT98), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n695), .A2(new_n696), .A3(G469), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n490), .A2(new_n495), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n697), .A2(new_n698), .A3(new_n604), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  AND4_X1   g514(.A1(new_n320), .A2(new_n372), .A3(new_n630), .A4(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT41), .B(G113), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G15));
  NAND2_X1  g517(.A1(new_n320), .A2(new_n372), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(new_n636), .A3(new_n700), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G116), .ZN(G18));
  NAND4_X1  g521(.A1(new_n616), .A2(new_n697), .A3(new_n698), .A4(new_n604), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n660), .A2(new_n567), .A3(new_n573), .A4(new_n602), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n320), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G119), .ZN(G21));
  AND4_X1   g526(.A1(new_n604), .A2(new_n697), .A3(new_n698), .A4(new_n573), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT100), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n714), .B1(new_n567), .B2(new_n602), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n556), .A2(new_n557), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n716), .B1(KEYINPUT20), .B2(new_n565), .ZN(new_n717));
  OAI211_X1 g531(.A(KEYINPUT100), .B(new_n601), .C1(new_n717), .C2(new_n535), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n715), .A2(new_n616), .A3(new_n718), .ZN(new_n719));
  XOR2_X1   g533(.A(new_n300), .B(KEYINPUT99), .Z(new_n720));
  AOI21_X1  g534(.A(new_n271), .B1(new_n284), .B2(new_n314), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n721), .B1(KEYINPUT31), .B2(new_n272), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n720), .B1(new_n304), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n611), .A2(new_n316), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n723), .B1(new_n724), .B2(G472), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n713), .A2(new_n719), .A3(new_n372), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G122), .ZN(G24));
  INV_X1    g541(.A(new_n708), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n728), .A2(new_n689), .A3(new_n660), .A4(new_n725), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G125), .ZN(G27));
  XOR2_X1   g544(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n731));
  NAND3_X1  g545(.A1(new_n442), .A2(new_n445), .A3(new_n443), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n732), .B1(new_n659), .B2(KEYINPUT101), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT101), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n658), .A2(new_n734), .A3(new_n604), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n733), .A2(new_n320), .A3(new_n372), .A4(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n689), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n731), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OR3_X1    g552(.A1(new_n306), .A2(KEYINPUT103), .A3(KEYINPUT32), .ZN(new_n739));
  OAI21_X1  g553(.A(KEYINPUT103), .B1(new_n306), .B2(KEYINPUT32), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n739), .A2(new_n319), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n372), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g557(.A(KEYINPUT101), .B1(new_n496), .B2(new_n605), .ZN(new_n744));
  INV_X1    g558(.A(new_n732), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n735), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n689), .A2(KEYINPUT42), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n743), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n738), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G131), .ZN(G33));
  NOR3_X1   g565(.A1(new_n704), .A2(new_n746), .A3(new_n664), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n211), .ZN(G36));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n452), .B1(new_n483), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n475), .A2(KEYINPUT45), .A3(new_n482), .ZN(new_n756));
  AOI22_X1  g570(.A1(new_n755), .A2(new_n756), .B1(G469), .B2(G902), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT104), .ZN(new_n758));
  OR3_X1    g572(.A1(new_n757), .A2(new_n758), .A3(KEYINPUT46), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n758), .B1(new_n757), .B2(KEYINPUT46), .ZN(new_n760));
  AOI22_X1  g574(.A1(new_n757), .A2(KEYINPUT46), .B1(new_n490), .B2(new_n495), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n759), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n762), .A2(new_n604), .A3(new_n670), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(KEYINPUT105), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n567), .A2(new_n628), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT43), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT43), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n567), .A2(new_n767), .A3(new_n628), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(new_n660), .A3(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n613), .A2(new_n769), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n770), .A2(KEYINPUT44), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(KEYINPUT44), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n732), .B(KEYINPUT106), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n764), .A2(new_n771), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G137), .ZN(G39));
  INV_X1    g589(.A(KEYINPUT47), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n776), .B1(new_n762), .B2(new_n604), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n762), .A2(new_n776), .A3(new_n604), .ZN(new_n779));
  NOR4_X1   g593(.A1(new_n737), .A2(new_n320), .A3(new_n372), .A4(new_n732), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G140), .ZN(G42));
  NAND3_X1  g596(.A1(new_n372), .A2(new_n445), .A3(new_n604), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n697), .A2(new_n698), .ZN(new_n784));
  AOI211_X1 g598(.A(new_n765), .B(new_n783), .C1(KEYINPUT49), .C2(new_n784), .ZN(new_n785));
  XOR2_X1   g599(.A(new_n785), .B(KEYINPUT107), .Z(new_n786));
  NOR2_X1   g600(.A1(new_n784), .A2(KEYINPUT49), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT108), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n786), .A2(new_n681), .A3(new_n684), .A4(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(KEYINPUT109), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n711), .A2(new_n651), .A3(new_n726), .ZN(new_n791));
  INV_X1    g605(.A(new_n701), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n610), .A2(new_n613), .A3(new_n573), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n445), .B1(new_n447), .B2(new_n448), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(KEYINPUT84), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n795), .A2(new_n449), .A3(new_n567), .A4(new_n601), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n706), .A2(new_n791), .A3(new_n792), .A4(new_n798), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n795), .A2(new_n688), .A3(new_n449), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n800), .A2(new_n573), .A3(new_n613), .A4(new_n610), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n607), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(KEYINPUT110), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT110), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n607), .A2(new_n801), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n799), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n689), .A2(new_n660), .A3(new_n725), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n302), .A2(new_n307), .A3(new_n319), .ZN(new_n809));
  AND4_X1   g623(.A1(new_n534), .A2(new_n634), .A3(new_n602), .A4(new_n663), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n668), .A2(new_n660), .A3(new_n745), .A4(new_n810), .ZN(new_n811));
  OAI22_X1  g625(.A1(new_n808), .A2(new_n746), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  AOI211_X1 g626(.A(new_n812), .B(new_n752), .C1(new_n738), .C2(new_n749), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n662), .B(new_n320), .C1(new_n665), .C2(new_n689), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n658), .A2(new_n604), .A3(new_n663), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n715), .A2(new_n616), .A3(new_n718), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n817), .A2(new_n649), .A3(new_n680), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n814), .A2(new_n818), .A3(new_n729), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT52), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n814), .A2(new_n818), .A3(new_n821), .A4(new_n729), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n807), .A2(new_n813), .A3(new_n823), .A4(KEYINPUT53), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(KEYINPUT111), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n752), .A2(new_n812), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n750), .A2(new_n820), .A3(new_n826), .A4(new_n822), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n711), .A2(new_n651), .A3(new_n726), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n828), .A2(new_n701), .A3(new_n797), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n829), .A2(new_n706), .A3(new_n803), .A4(new_n805), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT111), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n831), .A2(new_n832), .A3(KEYINPUT53), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n834), .B1(new_n827), .B2(new_n830), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n825), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n836), .A2(KEYINPUT112), .A3(KEYINPUT54), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT112), .B1(new_n836), .B2(KEYINPUT54), .ZN(new_n838));
  XNOR2_X1  g652(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n824), .A2(new_n835), .A3(new_n839), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n837), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT115), .ZN(new_n843));
  INV_X1    g657(.A(new_n779), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n843), .B1(new_n844), .B2(new_n777), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n778), .A2(KEYINPUT115), .A3(new_n779), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n784), .A2(new_n604), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n845), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n725), .A2(new_n372), .ZN(new_n850));
  INV_X1    g664(.A(new_n569), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n766), .A2(new_n851), .A3(new_n768), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(new_n773), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(KEYINPUT114), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n849), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n699), .A2(new_n732), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n725), .A2(new_n660), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n859), .A2(new_n860), .A3(new_n852), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n684), .A2(new_n700), .A3(new_n615), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n853), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT50), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n853), .A2(new_n862), .A3(KEYINPUT50), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n861), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n371), .A2(new_n569), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n619), .A2(new_n628), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n681), .A2(new_n858), .A3(new_n868), .A4(new_n869), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT116), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT51), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n867), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n847), .B1(new_n778), .B2(new_n779), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n867), .B(new_n871), .C1(new_n855), .C2(new_n874), .ZN(new_n875));
  AOI22_X1  g689(.A1(new_n857), .A2(new_n873), .B1(new_n875), .B2(KEYINPUT51), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n742), .A2(new_n852), .A3(new_n859), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n877), .B(KEYINPUT48), .Z(new_n878));
  NAND2_X1  g692(.A1(new_n853), .A2(new_n728), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(KEYINPUT117), .Z(new_n880));
  NAND2_X1  g694(.A1(new_n858), .A2(new_n868), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n881), .A2(new_n629), .A3(new_n680), .ZN(new_n882));
  INV_X1    g696(.A(G952), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n882), .A2(new_n883), .A3(G953), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n878), .A2(new_n880), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n842), .B1(new_n876), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n885), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n875), .A2(KEYINPUT51), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n867), .A2(new_n871), .A3(new_n872), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n889), .B1(new_n856), .B2(new_n849), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n887), .B(KEYINPUT118), .C1(new_n888), .C2(new_n890), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n886), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT119), .B1(new_n841), .B2(new_n892), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n827), .A2(new_n830), .A3(new_n834), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n835), .B1(new_n894), .B2(new_n832), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n824), .A2(KEYINPUT111), .ZN(new_n896));
  OAI21_X1  g710(.A(KEYINPUT54), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT112), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n840), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n836), .A2(KEYINPUT112), .A3(KEYINPUT54), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n899), .A2(KEYINPUT119), .A3(new_n900), .A4(new_n892), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n883), .A2(new_n357), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n790), .B1(new_n893), .B2(new_n903), .ZN(G75));
  NAND2_X1  g718(.A1(new_n416), .A2(new_n423), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(new_n421), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT55), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT56), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n316), .B1(new_n824), .B2(new_n835), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n910), .A2(G210), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n911), .A2(KEYINPUT120), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(KEYINPUT120), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n909), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n357), .A2(G952), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(KEYINPUT121), .Z(new_n916));
  NOR2_X1   g730(.A1(new_n911), .A2(KEYINPUT56), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n916), .B1(new_n917), .B2(new_n907), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n914), .A2(new_n918), .ZN(G51));
  NAND2_X1  g733(.A1(new_n824), .A2(new_n835), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(new_n839), .ZN(new_n921));
  NAND2_X1  g735(.A1(G469), .A2(G902), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT122), .Z(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT57), .ZN(new_n924));
  OAI22_X1  g738(.A1(new_n921), .A2(new_n924), .B1(new_n487), .B2(new_n486), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n910), .A2(new_n756), .A3(new_n755), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n915), .B1(new_n925), .B2(new_n926), .ZN(G54));
  NAND3_X1  g741(.A1(new_n910), .A2(KEYINPUT58), .A3(G475), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n561), .A2(new_n564), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n928), .A2(new_n929), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n930), .A2(new_n931), .A3(new_n915), .ZN(G60));
  NAND2_X1  g746(.A1(G478), .A2(G902), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT59), .Z(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n623), .A2(new_n625), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n916), .B1(new_n921), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n899), .A2(new_n900), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n935), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n937), .B1(new_n939), .B2(new_n626), .ZN(G63));
  NAND2_X1  g754(.A1(G217), .A2(G902), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT60), .Z(new_n942));
  NAND2_X1  g756(.A1(new_n920), .A2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n363), .ZN(new_n944));
  INV_X1    g758(.A(new_n361), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n645), .A2(new_n647), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n946), .B(new_n916), .C1(new_n947), .C2(new_n943), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT61), .Z(G66));
  AOI21_X1  g763(.A(new_n357), .B1(new_n571), .B2(G224), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT123), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n951), .B1(new_n807), .B2(G953), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n905), .B1(G898), .B2(new_n357), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(G69));
  NAND3_X1  g768(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n547), .A2(new_n548), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n292), .B(new_n956), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n814), .A2(new_n729), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n686), .A2(new_n958), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n960), .A2(new_n357), .A3(new_n781), .A4(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n567), .A2(new_n601), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n732), .B1(new_n629), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n672), .A2(new_n705), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n774), .A2(new_n965), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT124), .Z(new_n967));
  OAI211_X1 g781(.A(new_n955), .B(new_n957), .C1(new_n962), .C2(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n774), .A2(new_n781), .A3(new_n958), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n764), .A2(new_n719), .A3(new_n743), .ZN(new_n970));
  OR2_X1    g784(.A1(new_n970), .A2(KEYINPUT125), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(KEYINPUT125), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n752), .B1(new_n738), .B2(new_n749), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT126), .Z(new_n975));
  AOI21_X1  g789(.A(G953), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n471), .A2(G900), .A3(G953), .ZN(new_n977));
  OR2_X1    g791(.A1(new_n957), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n968), .B1(new_n976), .B2(new_n978), .ZN(G72));
  NAND2_X1  g793(.A1(G472), .A2(G902), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT63), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT127), .Z(new_n982));
  NAND4_X1  g796(.A1(new_n960), .A2(new_n781), .A3(new_n807), .A4(new_n961), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n982), .B1(new_n983), .B2(new_n967), .ZN(new_n984));
  INV_X1    g798(.A(new_n675), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n836), .ZN(new_n987));
  NOR4_X1   g801(.A1(new_n987), .A2(new_n312), .A3(new_n985), .A4(new_n981), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n676), .A2(new_n257), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n973), .A2(new_n807), .A3(new_n975), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n989), .B1(new_n990), .B2(new_n982), .ZN(new_n991));
  NOR4_X1   g805(.A1(new_n986), .A2(new_n915), .A3(new_n988), .A4(new_n991), .ZN(G57));
endmodule


