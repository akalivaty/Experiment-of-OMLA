//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1 1 0 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1221, new_n1222, new_n1223, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n207));
  INV_X1    g0007(.A(G58), .ZN(new_n208));
  INV_X1    g0008(.A(G232), .ZN(new_n209));
  INV_X1    g0009(.A(G97), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n206), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT1), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n206), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(new_n201), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G50), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(new_n220), .A2(new_n221), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n228), .B1(new_n220), .B2(new_n221), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n217), .A2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT65), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(KEYINPUT66), .Z(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n235), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT67), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(KEYINPUT68), .ZN(new_n249));
  NOR2_X1   g0049(.A1(G41), .A2(G45), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n249), .B1(new_n250), .B2(G1), .ZN(new_n251));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  OAI211_X1 g0052(.A(new_n252), .B(KEYINPUT68), .C1(G41), .C2(G45), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G274), .ZN(new_n255));
  AND2_X1   g0055(.A1(G1), .A2(G13), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  INV_X1    g0061(.A(G45), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n252), .A2(new_n263), .B1(new_n256), .B2(new_n257), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n260), .B1(G226), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  OR2_X1    g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AND2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NOR2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n269), .A2(G223), .B1(new_n272), .B2(G77), .ZN(new_n273));
  INV_X1    g0073(.A(G222), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n267), .A2(new_n268), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n266), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n273), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n256), .A2(new_n257), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n265), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT9), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n252), .A2(G13), .A3(G20), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(new_n222), .A3(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n223), .A2(G1), .ZN(new_n286));
  NOR3_X1   g0086(.A1(new_n285), .A2(new_n202), .A3(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n283), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n287), .B1(new_n202), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n203), .A2(G20), .ZN(new_n290));
  INV_X1    g0090(.A(G150), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G20), .A2(G33), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n223), .A2(G33), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT8), .B(G58), .ZN(new_n295));
  OAI221_X1 g0095(.A(new_n290), .B1(new_n291), .B2(new_n293), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n284), .A2(new_n222), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n289), .A2(new_n298), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n281), .A2(G200), .B1(new_n282), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G190), .ZN(new_n301));
  INV_X1    g0101(.A(new_n299), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT9), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n303), .A2(KEYINPUT72), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n303), .A2(KEYINPUT72), .ZN(new_n305));
  OAI221_X1 g0105(.A(new_n300), .B1(new_n301), .B2(new_n281), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n306), .B(KEYINPUT10), .ZN(new_n307));
  INV_X1    g0107(.A(G169), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n302), .B1(new_n281), .B2(new_n308), .ZN(new_n309));
  AND2_X1   g0109(.A1(KEYINPUT69), .A2(G179), .ZN(new_n310));
  NOR2_X1   g0110(.A1(KEYINPUT69), .A2(G179), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n265), .A2(new_n280), .A3(new_n312), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n307), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G77), .ZN(new_n317));
  OAI22_X1  g0117(.A1(new_n295), .A2(new_n293), .B1(new_n223), .B2(new_n317), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT15), .B(G87), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n319), .A2(new_n294), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n297), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n285), .ZN(new_n322));
  INV_X1    g0122(.A(new_n286), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n322), .A2(G77), .A3(new_n323), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n321), .B(new_n324), .C1(G77), .C2(new_n283), .ZN(new_n325));
  XOR2_X1   g0125(.A(new_n325), .B(KEYINPUT71), .Z(new_n326));
  INV_X1    g0126(.A(KEYINPUT70), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n260), .B1(G244), .B2(new_n264), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n269), .A2(G238), .B1(new_n272), .B2(G107), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n329), .B1(new_n209), .B2(new_n276), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n279), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n327), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n328), .A2(new_n331), .A3(new_n327), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n326), .B1(new_n335), .B2(new_n308), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n333), .A2(new_n334), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n312), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  OAI22_X1  g0139(.A1(new_n293), .A2(new_n202), .B1(new_n223), .B2(G68), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n294), .A2(new_n317), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n297), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT11), .ZN(new_n343));
  OR2_X1    g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n343), .ZN(new_n345));
  INV_X1    g0145(.A(G68), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n288), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n347), .B(KEYINPUT12), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n322), .A2(G68), .A3(new_n323), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n344), .A2(new_n345), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT14), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n209), .A2(G1698), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(G226), .B2(G1698), .ZN(new_n353));
  INV_X1    g0153(.A(G33), .ZN(new_n354));
  OAI22_X1  g0154(.A1(new_n353), .A2(new_n272), .B1(new_n354), .B2(new_n210), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n355), .A2(new_n279), .B1(G238), .B2(new_n264), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT13), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n259), .A2(KEYINPUT73), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n259), .A2(KEYINPUT73), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n356), .B(new_n357), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  XNOR2_X1  g0161(.A(new_n259), .B(KEYINPUT73), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n357), .B1(new_n362), .B2(new_n356), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n351), .B(G169), .C1(new_n361), .C2(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n356), .B1(new_n358), .B2(new_n359), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(KEYINPUT13), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n366), .A2(G179), .A3(new_n360), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(new_n360), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n351), .B1(new_n369), .B2(G169), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n350), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n369), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n350), .B1(new_n372), .B2(G190), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n369), .A2(G200), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n337), .A2(G190), .ZN(new_n376));
  INV_X1    g0176(.A(G200), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n376), .B(new_n326), .C1(new_n377), .C2(new_n337), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n339), .A2(new_n371), .A3(new_n375), .A4(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n295), .A2(new_n286), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n322), .A2(new_n380), .B1(new_n288), .B2(new_n295), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n297), .ZN(new_n383));
  AOI21_X1  g0183(.A(KEYINPUT7), .B1(new_n272), .B2(new_n223), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT7), .ZN(new_n385));
  NOR4_X1   g0185(.A1(new_n270), .A2(new_n271), .A3(new_n385), .A4(G20), .ZN(new_n386));
  OAI21_X1  g0186(.A(G68), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n208), .A2(new_n346), .ZN(new_n388));
  OAI21_X1  g0188(.A(G20), .B1(new_n388), .B2(new_n201), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n292), .A2(G159), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT16), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n383), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n387), .A2(KEYINPUT16), .A3(new_n392), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n382), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI211_X1 g0197(.A(G223), .B(new_n266), .C1(new_n270), .C2(new_n271), .ZN(new_n398));
  OAI211_X1 g0198(.A(G226), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n399));
  NAND2_X1  g0199(.A1(G33), .A2(G87), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n279), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n254), .A2(new_n258), .B1(new_n264), .B2(G232), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n312), .ZN(new_n405));
  AOI21_X1  g0205(.A(G169), .B1(new_n402), .B2(new_n403), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT18), .B1(new_n397), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n385), .B1(new_n275), .B2(G20), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n272), .A2(KEYINPUT7), .A3(new_n223), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n346), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n394), .B1(new_n412), .B2(new_n391), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n413), .A2(new_n297), .A3(new_n396), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n381), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT18), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n406), .B1(new_n312), .B2(new_n404), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT17), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n402), .A2(new_n403), .A3(new_n301), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n404), .B2(G200), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n419), .B1(new_n397), .B2(new_n421), .ZN(new_n422));
  XOR2_X1   g0222(.A(KEYINPUT74), .B(KEYINPUT17), .Z(new_n423));
  AND4_X1   g0223(.A1(new_n414), .A2(new_n421), .A3(new_n381), .A4(new_n423), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n409), .B(new_n418), .C1(new_n422), .C2(new_n424), .ZN(new_n425));
  NOR3_X1   g0225(.A1(new_n316), .A2(new_n379), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT77), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(new_n354), .B2(G1), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n252), .A2(KEYINPUT77), .A3(G33), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n322), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n432), .A2(new_n210), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n288), .A2(new_n210), .ZN(new_n434));
  XNOR2_X1  g0234(.A(new_n434), .B(KEYINPUT76), .ZN(new_n435));
  OR2_X1    g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(G107), .B1(new_n384), .B2(new_n386), .ZN(new_n437));
  XNOR2_X1  g0237(.A(G97), .B(G107), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT75), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n438), .B1(new_n439), .B2(KEYINPUT6), .ZN(new_n440));
  MUX2_X1   g0240(.A(new_n439), .B(G97), .S(KEYINPUT6), .Z(new_n441));
  OAI21_X1  g0241(.A(new_n440), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  OAI221_X1 g0242(.A(new_n437), .B1(new_n317), .B2(new_n293), .C1(new_n223), .C2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n436), .B1(new_n443), .B2(new_n297), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n252), .A2(G45), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT5), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n261), .ZN(new_n447));
  NAND2_X1  g0247(.A1(KEYINPUT5), .A2(G41), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n445), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NOR3_X1   g0249(.A1(new_n449), .A2(new_n279), .A3(new_n211), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n269), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n451));
  OAI211_X1 g0251(.A(G244), .B(new_n266), .C1(new_n270), .C2(new_n271), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT4), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n453), .A2(G1698), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n455), .B(G244), .C1(new_n271), .C2(new_n270), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT78), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT78), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n275), .A2(new_n458), .A3(G244), .A4(new_n455), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n451), .A2(new_n454), .A3(new_n457), .A4(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n450), .B1(new_n460), .B2(new_n279), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT79), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n449), .A2(new_n258), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n461), .A2(new_n462), .A3(G190), .A4(new_n463), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n444), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n377), .B1(new_n461), .B2(new_n463), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n461), .A2(new_n463), .ZN(new_n467));
  OAI22_X1  g0267(.A1(new_n466), .A2(KEYINPUT79), .B1(new_n467), .B2(new_n301), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n461), .A2(new_n312), .A3(new_n463), .ZN(new_n469));
  OAI22_X1  g0269(.A1(new_n442), .A2(new_n223), .B1(new_n317), .B2(new_n293), .ZN(new_n470));
  INV_X1    g0270(.A(new_n437), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n297), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n433), .A2(new_n435), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n467), .A2(new_n308), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n465), .A2(new_n468), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n275), .A2(G257), .A3(G1698), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G33), .A2(G294), .ZN(new_n477));
  OAI211_X1 g0277(.A(G250), .B(new_n266), .C1(new_n270), .C2(new_n271), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n279), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n262), .A2(G1), .ZN(new_n481));
  INV_X1    g0281(.A(new_n448), .ZN(new_n482));
  NOR2_X1   g0282(.A1(KEYINPUT5), .A2(G41), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n484), .A2(G264), .A3(new_n278), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n463), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(G179), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n480), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n486), .B1(new_n279), .B2(new_n479), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n489), .B1(new_n490), .B2(G169), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n223), .B(G87), .C1(new_n270), .C2(new_n271), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT22), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT22), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n275), .A2(new_n494), .A3(new_n223), .A4(G87), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT24), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G33), .A2(G116), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n498), .A2(G20), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT23), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(new_n223), .B2(G107), .ZN(new_n501));
  INV_X1    g0301(.A(G107), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n502), .A2(KEYINPUT23), .A3(G20), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n499), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n496), .A2(new_n497), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n497), .B1(new_n496), .B2(new_n504), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n297), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n285), .A2(new_n430), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT25), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n283), .B2(G107), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n288), .A2(KEYINPUT25), .A3(new_n502), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n508), .A2(G107), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n491), .B1(new_n507), .B2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT83), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n480), .A2(new_n487), .A3(new_n301), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(new_n490), .B2(G200), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n517), .A2(new_n507), .A3(new_n512), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n514), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n518), .ZN(new_n520));
  OAI21_X1  g0320(.A(KEYINPUT83), .B1(new_n520), .B2(new_n513), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n447), .A2(new_n448), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n523), .A2(new_n481), .B1(new_n256), .B2(new_n257), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n524), .A2(G270), .B1(new_n258), .B2(new_n449), .ZN(new_n525));
  OAI211_X1 g0325(.A(G264), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n526));
  OAI211_X1 g0326(.A(G257), .B(new_n266), .C1(new_n270), .C2(new_n271), .ZN(new_n527));
  INV_X1    g0327(.A(G303), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n526), .B(new_n527), .C1(new_n528), .C2(new_n275), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n279), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(G200), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n322), .A2(new_n431), .A3(G116), .ZN(new_n533));
  INV_X1    g0333(.A(G116), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n288), .A2(new_n534), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n284), .A2(new_n222), .B1(G20), .B2(new_n534), .ZN(new_n536));
  AOI21_X1  g0336(.A(G20), .B1(G33), .B2(G283), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(G33), .B2(new_n210), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n536), .A2(new_n538), .A3(KEYINPUT20), .ZN(new_n539));
  AOI21_X1  g0339(.A(KEYINPUT20), .B1(new_n536), .B2(new_n538), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n533), .B(new_n535), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n525), .A2(new_n530), .A3(G190), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n532), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  XNOR2_X1  g0344(.A(new_n544), .B(KEYINPUT82), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n531), .A2(new_n541), .A3(G169), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT21), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n541), .A2(G179), .A3(new_n530), .A4(new_n525), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n531), .A2(new_n541), .A3(KEYINPUT21), .A4(G169), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(G87), .A2(G97), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n502), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(KEYINPUT80), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT80), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n553), .A2(new_n556), .A3(new_n502), .ZN(new_n557));
  NAND3_X1  g0357(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n555), .A2(new_n557), .B1(new_n223), .B2(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n223), .B(G68), .C1(new_n270), .C2(new_n271), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT19), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n561), .B1(new_n294), .B2(new_n210), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n297), .B1(new_n559), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n319), .A2(new_n288), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n508), .A2(G87), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n275), .A2(G244), .A3(G1698), .ZN(new_n569));
  OAI211_X1 g0369(.A(G238), .B(new_n266), .C1(new_n270), .C2(new_n271), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(new_n498), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n279), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n258), .A2(new_n481), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n278), .A2(G250), .A3(new_n445), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(G200), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n568), .B(new_n578), .C1(new_n301), .C2(new_n577), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n558), .A2(new_n223), .ZN(new_n580));
  NOR4_X1   g0380(.A1(KEYINPUT80), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n556), .B1(new_n553), .B2(new_n502), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n583), .A2(new_n560), .A3(new_n562), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n584), .A2(new_n297), .B1(new_n288), .B2(new_n319), .ZN(new_n585));
  OAI21_X1  g0385(.A(KEYINPUT81), .B1(new_n432), .B2(new_n319), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT81), .ZN(new_n587));
  INV_X1    g0387(.A(new_n319), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n508), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n585), .A2(new_n586), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n577), .A2(new_n308), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n575), .B1(new_n571), .B2(new_n279), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n312), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n579), .A2(new_n594), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n545), .A2(new_n552), .A3(new_n595), .ZN(new_n596));
  AND4_X1   g0396(.A1(new_n426), .A2(new_n475), .A3(new_n522), .A4(new_n596), .ZN(G372));
  NAND2_X1  g0397(.A1(new_n575), .A2(KEYINPUT84), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT84), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n573), .A2(new_n599), .A3(new_n574), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n572), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n308), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n590), .A2(new_n602), .A3(new_n593), .ZN(new_n603));
  XNOR2_X1  g0403(.A(new_n603), .B(KEYINPUT86), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n513), .A2(new_n551), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n601), .A2(G200), .B1(G190), .B2(new_n592), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT85), .B1(new_n585), .B2(new_n566), .ZN(new_n607));
  AND4_X1   g0407(.A1(KEYINPUT85), .A2(new_n564), .A3(new_n565), .A4(new_n566), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n609), .A2(new_n518), .A3(new_n603), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n604), .B1(new_n611), .B2(new_n475), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n474), .A2(new_n469), .A3(new_n594), .A4(new_n579), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT26), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n467), .A2(new_n308), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n472), .A2(new_n473), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(new_n469), .A3(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT26), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT85), .ZN(new_n620));
  XNOR2_X1  g0420(.A(new_n567), .B(new_n620), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n586), .A2(new_n589), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n622), .A2(new_n585), .B1(new_n312), .B2(new_n592), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n621), .A2(new_n606), .B1(new_n623), .B2(new_n602), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n618), .A2(new_n619), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n612), .A2(new_n614), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n426), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n371), .ZN(new_n628));
  INV_X1    g0428(.A(new_n339), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n628), .B1(new_n629), .B2(new_n375), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n422), .A2(new_n424), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n409), .B(new_n418), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n314), .B1(new_n632), .B2(new_n307), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n627), .A2(new_n633), .ZN(G369));
  NAND3_X1  g0434(.A1(new_n252), .A2(new_n223), .A3(G13), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n635), .A2(KEYINPUT27), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(KEYINPUT27), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(new_n637), .A3(G213), .ZN(new_n638));
  INV_X1    g0438(.A(G343), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n551), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n519), .B2(new_n521), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n643), .B1(new_n513), .B2(new_n641), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n551), .A2(new_n542), .A3(new_n641), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n545), .A2(new_n552), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n646), .A2(KEYINPUT87), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n646), .A2(KEYINPUT87), .B1(new_n541), .B2(new_n640), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(G330), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n507), .A2(new_n512), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n522), .B1(new_n651), .B2(new_n641), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n513), .A2(new_n640), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n644), .B1(new_n650), .B2(new_n655), .ZN(G399));
  INV_X1    g0456(.A(new_n218), .ZN(new_n657));
  OAI21_X1  g0457(.A(KEYINPUT88), .B1(new_n657), .B2(G41), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n657), .A2(KEYINPUT88), .A3(G41), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G1), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n555), .A2(new_n534), .A3(new_n557), .ZN(new_n664));
  OAI22_X1  g0464(.A1(new_n663), .A2(new_n664), .B1(new_n226), .B2(new_n662), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n665), .B(KEYINPUT28), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n522), .A2(new_n596), .A3(new_n475), .A4(new_n641), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT90), .ZN(new_n668));
  INV_X1    g0468(.A(new_n312), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n669), .B1(new_n525), .B2(new_n530), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n601), .B2(KEYINPUT89), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT89), .ZN(new_n672));
  INV_X1    g0472(.A(new_n600), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n599), .B1(new_n573), .B2(new_n574), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n672), .B1(new_n675), .B2(new_n572), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n668), .B1(new_n671), .B2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n490), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n601), .A2(KEYINPUT89), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n675), .A2(new_n672), .A3(new_n572), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n679), .A2(new_n680), .A3(KEYINPUT90), .A4(new_n670), .ZN(new_n681));
  AND4_X1   g0481(.A1(new_n467), .A2(new_n677), .A3(new_n678), .A4(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n531), .A2(new_n488), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n683), .A2(new_n461), .A3(new_n490), .A4(new_n592), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT30), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n684), .B(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n640), .B1(new_n682), .B2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT31), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OAI211_X1 g0489(.A(KEYINPUT31), .B(new_n640), .C1(new_n682), .C2(new_n686), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n667), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G330), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT92), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n618), .A2(new_n624), .A3(KEYINPUT91), .A4(KEYINPUT26), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT91), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n696), .B1(new_n613), .B2(new_n619), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n609), .A2(new_n603), .ZN(new_n698));
  NOR3_X1   g0498(.A1(new_n698), .A2(new_n617), .A3(new_n619), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n695), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n612), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n694), .B1(new_n701), .B2(new_n641), .ZN(new_n702));
  AOI211_X1 g0502(.A(KEYINPUT92), .B(new_n640), .C1(new_n700), .C2(new_n612), .ZN(new_n703));
  OAI21_X1  g0503(.A(KEYINPUT29), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n626), .A2(new_n641), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT29), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n693), .B1(new_n704), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n666), .B1(new_n708), .B2(G1), .ZN(G364));
  AND2_X1   g0509(.A1(new_n223), .A2(G13), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n252), .B1(new_n710), .B2(G45), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n661), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n657), .A2(new_n272), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G355), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n715), .B1(G116), .B2(new_n218), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n244), .A2(G45), .ZN(new_n717));
  XOR2_X1   g0517(.A(new_n717), .B(KEYINPUT93), .Z(new_n718));
  NOR2_X1   g0518(.A1(new_n657), .A2(new_n275), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n720), .B1(new_n262), .B2(new_n227), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n716), .B1(new_n718), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(G13), .A2(G33), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(G20), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n222), .B1(G20), .B2(new_n308), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n713), .B1(new_n722), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n312), .A2(G200), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n223), .A2(G190), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(KEYINPUT95), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n732), .A2(KEYINPUT95), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n223), .A2(new_n377), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n669), .A2(G190), .A3(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AOI22_X1  g0540(.A1(new_n737), .A2(G77), .B1(G50), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n223), .A2(new_n301), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n730), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(KEYINPUT94), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n744), .A2(KEYINPUT94), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n741), .B1(new_n208), .B2(new_n748), .ZN(new_n749));
  XOR2_X1   g0549(.A(new_n749), .B(KEYINPUT96), .Z(new_n750));
  NOR2_X1   g0550(.A1(new_n377), .A2(G179), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n731), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT97), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G107), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n742), .A2(new_n751), .ZN(new_n755));
  INV_X1    g0555(.A(G87), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n275), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G179), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G190), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n757), .B1(G97), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n731), .A2(new_n758), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G159), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT32), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n669), .A2(new_n301), .A3(new_n738), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n765), .B1(G68), .B2(new_n767), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n750), .A2(new_n754), .A3(new_n761), .A4(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G326), .ZN(new_n770));
  INV_X1    g0570(.A(new_n760), .ZN(new_n771));
  INV_X1    g0571(.A(G294), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n739), .A2(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n773), .B1(new_n737), .B2(G311), .ZN(new_n774));
  XOR2_X1   g0574(.A(new_n774), .B(KEYINPUT98), .Z(new_n775));
  OAI21_X1  g0575(.A(new_n272), .B1(new_n755), .B2(new_n528), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n776), .B1(G329), .B2(new_n763), .ZN(new_n777));
  INV_X1    g0577(.A(new_n753), .ZN(new_n778));
  INV_X1    g0578(.A(G283), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g0580(.A(KEYINPUT33), .B(G317), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n780), .B1(new_n767), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G322), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n782), .B1(new_n783), .B2(new_n748), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n769), .B1(new_n775), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n729), .B1(new_n785), .B2(new_n726), .ZN(new_n786));
  INV_X1    g0586(.A(new_n725), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n786), .B1(new_n649), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n713), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n650), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n649), .A2(G330), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n788), .B1(new_n790), .B2(new_n791), .ZN(G396));
  NAND2_X1  g0592(.A1(new_n335), .A2(new_n308), .ZN(new_n793));
  INV_X1    g0593(.A(new_n326), .ZN(new_n794));
  AND4_X1   g0594(.A1(new_n338), .A2(new_n793), .A3(new_n794), .A4(new_n641), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n378), .B1(new_n326), .B2(new_n641), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n795), .B1(new_n796), .B2(new_n339), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n705), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n797), .A2(new_n626), .A3(new_n641), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n713), .B1(new_n801), .B2(new_n692), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n692), .B2(new_n801), .ZN(new_n803));
  INV_X1    g0603(.A(G311), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n272), .B1(new_n762), .B2(new_n804), .C1(new_n502), .C2(new_n755), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n753), .A2(G87), .ZN(new_n806));
  XOR2_X1   g0606(.A(KEYINPUT99), .B(G283), .Z(new_n807));
  OAI221_X1 g0607(.A(new_n806), .B1(new_n528), .B2(new_n739), .C1(new_n766), .C2(new_n807), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n805), .B(new_n808), .C1(G97), .C2(new_n760), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n809), .B1(new_n534), .B2(new_n736), .C1(new_n772), .C2(new_n748), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT100), .Z(new_n811));
  INV_X1    g0611(.A(G137), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n812), .A2(new_n739), .B1(new_n766), .B2(new_n291), .ZN(new_n813));
  INV_X1    g0613(.A(G159), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n736), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n748), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n813), .B(new_n815), .C1(G143), .C2(new_n816), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n817), .A2(KEYINPUT34), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n817), .A2(KEYINPUT34), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n755), .A2(new_n202), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n272), .B(new_n820), .C1(G132), .C2(new_n763), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n753), .A2(G68), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n821), .B(new_n822), .C1(new_n208), .C2(new_n771), .ZN(new_n823));
  NOR3_X1   g0623(.A1(new_n818), .A2(new_n819), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n726), .B1(new_n811), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n726), .A2(new_n723), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n789), .B1(new_n317), .B2(new_n826), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n825), .B(new_n827), .C1(new_n724), .C2(new_n797), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n803), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(G384));
  INV_X1    g0630(.A(KEYINPUT35), .ZN(new_n831));
  OAI211_X1 g0631(.A(G116), .B(new_n224), .C1(new_n442), .C2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(new_n831), .B2(new_n442), .ZN(new_n833));
  XNOR2_X1  g0633(.A(KEYINPUT101), .B(KEYINPUT36), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n833), .B(new_n834), .ZN(new_n835));
  OR3_X1    g0635(.A1(new_n226), .A2(new_n317), .A3(new_n388), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n202), .A2(G68), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n252), .B(G13), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n638), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n415), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n409), .A2(new_n418), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n842), .B1(new_n631), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(KEYINPUT103), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n397), .A2(new_n421), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n415), .A2(new_n417), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n846), .A2(new_n847), .A3(new_n841), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(KEYINPUT37), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT37), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n846), .A2(new_n847), .A3(new_n841), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT103), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n425), .A2(new_n853), .A3(new_n842), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n845), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT38), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT104), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n425), .A2(new_n853), .A3(new_n842), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n853), .B1(new_n425), .B2(new_n842), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n856), .B1(new_n849), .B2(new_n851), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n858), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n845), .A2(new_n858), .A3(new_n854), .A4(new_n862), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n857), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n371), .A2(KEYINPUT102), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT102), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n868), .B(new_n350), .C1(new_n368), .C2(new_n370), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n350), .A2(new_n640), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n373), .B2(new_n374), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n867), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n368), .A2(new_n370), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n375), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n870), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n691), .A2(new_n876), .A3(new_n797), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT40), .B1(new_n866), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT40), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n845), .A2(new_n854), .A3(new_n862), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n852), .A2(new_n844), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n856), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n879), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n878), .B1(new_n877), .B2(new_n883), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n426), .A2(new_n691), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n884), .A2(new_n885), .ZN(new_n887));
  INV_X1    g0687(.A(G330), .ZN(new_n888));
  NOR3_X1   g0688(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n843), .A2(new_n638), .ZN(new_n890));
  INV_X1    g0690(.A(new_n795), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n800), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n876), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n880), .A2(KEYINPUT104), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n894), .A2(new_n864), .B1(new_n856), .B2(new_n855), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n890), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n640), .B1(new_n867), .B2(new_n869), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n880), .A2(new_n882), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT39), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n895), .B2(new_n900), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n896), .B1(new_n897), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n704), .A2(new_n426), .A3(new_n707), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n633), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n903), .B(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n889), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n889), .A2(new_n906), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT105), .ZN(new_n909));
  OAI221_X1 g0709(.A(new_n907), .B1(new_n252), .B2(new_n710), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n908), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n911), .A2(KEYINPUT105), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n839), .B1(new_n910), .B2(new_n912), .ZN(G367));
  NOR2_X1   g0713(.A1(new_n621), .A2(new_n641), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n698), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n604), .B2(new_n914), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n725), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n234), .A2(new_n720), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n728), .B1(new_n657), .B2(new_n588), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n789), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n760), .A2(G68), .ZN(new_n921));
  AOI22_X1  g0721(.A1(G143), .A2(new_n740), .B1(new_n767), .B2(G159), .ZN(new_n922));
  INV_X1    g0722(.A(new_n755), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n272), .B1(new_n923), .B2(G58), .ZN(new_n924));
  INV_X1    g0724(.A(new_n752), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n925), .A2(G77), .B1(new_n763), .B2(G137), .ZN(new_n926));
  AND4_X1   g0726(.A1(new_n921), .A2(new_n922), .A3(new_n924), .A4(new_n926), .ZN(new_n927));
  OAI221_X1 g0727(.A(new_n927), .B1(new_n202), .B2(new_n736), .C1(new_n291), .C2(new_n748), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n748), .A2(new_n528), .B1(new_n804), .B2(new_n739), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n929), .B(KEYINPUT108), .Z(new_n930));
  INV_X1    g0730(.A(KEYINPUT109), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT46), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n755), .B2(new_n534), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n767), .A2(G294), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n931), .B2(new_n933), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n755), .A2(new_n932), .A3(new_n534), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(G107), .B2(new_n760), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n275), .B1(new_n763), .B2(G317), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n937), .B(new_n938), .C1(new_n210), .C2(new_n752), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n935), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n736), .B2(new_n807), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n928), .B1(new_n930), .B2(new_n941), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT47), .Z(new_n943));
  INV_X1    g0743(.A(new_n726), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n917), .B(new_n920), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n475), .B1(new_n444), .B2(new_n641), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT106), .Z(new_n947));
  NAND2_X1  g0747(.A1(new_n618), .A2(new_n640), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n949), .A2(new_n644), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT44), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n644), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT45), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n952), .B(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n650), .A2(new_n655), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n955), .B(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n643), .B1(new_n655), .B2(new_n642), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(new_n650), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n708), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n708), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n661), .B(KEYINPUT41), .Z(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n712), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n949), .A2(new_n643), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(KEYINPUT42), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n617), .B1(new_n947), .B2(new_n514), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n641), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n965), .A2(KEYINPUT42), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT43), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n969), .A2(new_n970), .B1(new_n971), .B2(new_n916), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n916), .A2(new_n971), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n972), .B(new_n973), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n949), .A2(new_n956), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n974), .B1(KEYINPUT107), .B2(new_n975), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n975), .B(KEYINPUT107), .Z(new_n977));
  OAI21_X1  g0777(.A(new_n976), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n945), .B1(new_n964), .B2(new_n978), .ZN(G387));
  OR2_X1    g0779(.A1(new_n239), .A2(new_n262), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n980), .A2(new_n719), .B1(new_n664), .B2(new_n714), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n295), .A2(G50), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT50), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n262), .B1(new_n346), .B2(new_n317), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n664), .B(new_n984), .C1(new_n983), .C2(new_n982), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n981), .A2(new_n985), .B1(G107), .B2(new_n218), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n789), .B1(new_n986), .B2(new_n727), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n654), .B2(new_n787), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n816), .A2(G50), .B1(G68), .B2(new_n737), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n275), .B1(new_n762), .B2(new_n291), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n771), .A2(new_n319), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n990), .B(new_n991), .C1(G77), .C2(new_n923), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n778), .A2(new_n210), .B1(new_n295), .B2(new_n766), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(G159), .B2(new_n740), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n989), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  AOI22_X1  g0795(.A1(G311), .A2(new_n767), .B1(new_n740), .B2(G322), .ZN(new_n996));
  INV_X1    g0796(.A(G317), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n996), .B1(new_n736), .B2(new_n528), .C1(new_n748), .C2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT48), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n998), .A2(new_n999), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n771), .A2(new_n807), .B1(new_n755), .B2(new_n772), .ZN(new_n1002));
  NOR3_X1   g0802(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(KEYINPUT49), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n275), .B1(new_n763), .B2(G326), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1004), .B(new_n1005), .C1(new_n534), .C2(new_n752), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1003), .A2(KEYINPUT49), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n995), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT110), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n988), .B1(new_n1009), .B2(new_n726), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(new_n959), .B2(new_n712), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n960), .A2(new_n661), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n959), .A2(new_n708), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1011), .B1(new_n1012), .B2(new_n1013), .ZN(G393));
  AND2_X1   g0814(.A1(new_n957), .A2(new_n960), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n661), .B1(new_n957), .B2(new_n960), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n957), .A2(new_n711), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n947), .A2(new_n725), .A3(new_n948), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n727), .B1(new_n210), .B2(new_n218), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(new_n247), .B2(new_n719), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n748), .A2(new_n814), .B1(new_n291), .B2(new_n739), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT51), .Z(new_n1023));
  NOR2_X1   g0823(.A1(new_n778), .A2(new_n756), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n771), .A2(new_n317), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n272), .B1(new_n763), .B2(G143), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n346), .B2(new_n755), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n766), .A2(new_n202), .ZN(new_n1028));
  NOR4_X1   g0828(.A1(new_n1024), .A2(new_n1025), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n295), .B2(new_n736), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n748), .A2(new_n804), .B1(new_n997), .B2(new_n739), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT52), .Z(new_n1032));
  AOI21_X1  g0832(.A(new_n275), .B1(new_n763), .B2(G322), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n754), .B(new_n1033), .C1(new_n755), .C2(new_n807), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT111), .Z(new_n1035));
  AOI22_X1  g0835(.A1(new_n767), .A2(G303), .B1(G116), .B2(new_n760), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1035), .B(new_n1036), .C1(new_n772), .C2(new_n736), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n1023), .A2(new_n1030), .B1(new_n1032), .B2(new_n1037), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n789), .B(new_n1021), .C1(new_n1038), .C2(new_n726), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1018), .B1(new_n1019), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1017), .A2(new_n1040), .ZN(G390));
  NAND3_X1  g0841(.A1(new_n693), .A2(new_n797), .A3(new_n876), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT112), .ZN(new_n1043));
  NOR3_X1   g0843(.A1(new_n702), .A2(new_n703), .A3(new_n795), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n796), .A2(new_n339), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1043), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n702), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n701), .A2(new_n694), .A3(new_n641), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1048), .A2(new_n1049), .A3(new_n891), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1050), .A2(KEYINPUT112), .A3(new_n1045), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1047), .A2(new_n1051), .A3(new_n876), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n899), .A2(new_n897), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n897), .B1(new_n892), .B2(new_n876), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n902), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1042), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1042), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1059), .B(new_n1056), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n712), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n822), .B1(new_n502), .B2(new_n766), .C1(new_n779), .C2(new_n739), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n272), .B1(new_n762), .B2(new_n772), .C1(new_n756), .C2(new_n755), .ZN(new_n1064));
  NOR3_X1   g0864(.A1(new_n1063), .A2(new_n1025), .A3(new_n1064), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(new_n210), .B2(new_n736), .C1(new_n534), .C2(new_n748), .ZN(new_n1066));
  OR3_X1    g0866(.A1(new_n755), .A2(KEYINPUT53), .A3(new_n291), .ZN(new_n1067));
  OAI21_X1  g0867(.A(KEYINPUT53), .B1(new_n755), .B2(new_n291), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1067), .B(new_n1068), .C1(new_n814), .C2(new_n771), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n272), .B1(new_n925), .B2(G50), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n763), .A2(G125), .ZN(new_n1071));
  INV_X1    g0871(.A(G128), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1070), .B(new_n1071), .C1(new_n1072), .C2(new_n739), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1069), .B(new_n1073), .C1(new_n816), .C2(G132), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT115), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(KEYINPUT54), .B(G143), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n737), .A2(new_n1077), .B1(G137), .B2(new_n767), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1074), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1078), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1080), .A2(KEYINPUT115), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1066), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n726), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n789), .B1(new_n295), .B2(new_n826), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1083), .B(new_n1084), .C1(new_n902), .C2(new_n724), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1062), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT113), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n876), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n692), .B2(new_n798), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n1042), .A2(new_n1089), .B1(new_n891), .B2(new_n800), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1042), .A2(new_n1089), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1090), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n426), .A2(new_n693), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n904), .A2(new_n633), .A3(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1087), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1096), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1092), .B1(new_n1047), .B2(new_n1051), .ZN(new_n1099));
  OAI211_X1 g0899(.A(KEYINPUT113), .B(new_n1098), .C1(new_n1099), .C2(new_n1090), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1101), .A2(KEYINPUT114), .ZN(new_n1102));
  OR2_X1    g0902(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n662), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1061), .B1(new_n1101), .B2(KEYINPUT114), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1086), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(G378));
  INV_X1    g0907(.A(KEYINPUT57), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1096), .B1(new_n1061), .B2(new_n1101), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n903), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n302), .A2(new_n638), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n316), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n316), .A2(new_n1113), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1112), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1116), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1118), .A2(new_n1114), .A3(new_n1111), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n883), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n691), .A2(new_n876), .A3(new_n797), .ZN(new_n1122));
  OAI21_X1  g0922(.A(G330), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(KEYINPUT120), .B1(new_n878), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n879), .B1(new_n895), .B2(new_n1122), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n888), .B1(new_n877), .B2(new_n883), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT120), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1120), .B1(new_n1124), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1127), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1110), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n1125), .A2(new_n1127), .A3(new_n1126), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1131), .B1(new_n1134), .B2(new_n1130), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1124), .A2(new_n1120), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1135), .A2(new_n903), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1133), .A2(new_n1137), .A3(KEYINPUT121), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT121), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1139), .B(new_n1110), .C1(new_n1129), .C2(new_n1132), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1108), .B1(new_n1109), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT123), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g0944(.A(KEYINPUT123), .B(new_n1108), .C1(new_n1109), .C2(new_n1141), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1109), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n1133), .A2(new_n1137), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1147), .A2(new_n1108), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n662), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1144), .A2(new_n1145), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n789), .B1(new_n202), .B2(new_n826), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n275), .A2(G41), .ZN(new_n1152));
  AOI211_X1 g0952(.A(G50), .B(new_n1152), .C1(new_n354), .C2(new_n261), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n748), .A2(new_n502), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT116), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(G77), .A2(new_n923), .B1(new_n763), .B2(G283), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n925), .A2(G58), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1156), .A2(new_n921), .A3(new_n1152), .A4(new_n1157), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n210), .A2(new_n766), .B1(new_n739), .B2(new_n534), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1158), .B(new_n1159), .C1(new_n737), .C2(new_n588), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1155), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT58), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1153), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT117), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n740), .A2(G125), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1165), .B1(new_n291), .B2(new_n771), .C1(new_n755), .C2(new_n1076), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(G132), .B2(new_n767), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n1167), .B1(new_n748), .B2(new_n1072), .C1(new_n812), .C2(new_n736), .ZN(new_n1168));
  XOR2_X1   g0968(.A(new_n1168), .B(KEYINPUT118), .Z(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(KEYINPUT59), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n925), .A2(G159), .ZN(new_n1172));
  AOI211_X1 g0972(.A(G33), .B(G41), .C1(new_n763), .C2(G124), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1170), .A2(KEYINPUT59), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1164), .B1(new_n1162), .B2(new_n1161), .C1(new_n1174), .C2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(KEYINPUT119), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n726), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1176), .A2(KEYINPUT119), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1151), .B1(new_n724), .B2(new_n1120), .C1(new_n1178), .C2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n1141), .B2(new_n711), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT122), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  OAI211_X1 g0983(.A(KEYINPUT122), .B(new_n1180), .C1(new_n1141), .C2(new_n711), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1150), .A2(new_n1185), .ZN(G375));
  INV_X1    g0986(.A(new_n1101), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n963), .A3(new_n1188), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n1189), .B(KEYINPUT124), .Z(new_n1190));
  INV_X1    g0990(.A(new_n1094), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1088), .A2(new_n723), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n736), .A2(new_n502), .B1(new_n534), .B2(new_n766), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT125), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n816), .A2(G283), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n778), .A2(new_n317), .B1(new_n772), .B2(new_n739), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n272), .B1(new_n762), .B2(new_n528), .C1(new_n210), .C2(new_n755), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n1198), .A2(new_n991), .A3(new_n1199), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .A4(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT126), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n755), .A2(new_n814), .B1(new_n762), .B2(new_n1072), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1157), .A2(new_n275), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1204), .B(new_n1205), .C1(G50), .C2(new_n760), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G132), .A2(new_n740), .B1(new_n767), .B2(new_n1077), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1208), .B1(new_n812), .B2(new_n748), .C1(new_n291), .C2(new_n736), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1203), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n1211), .A2(new_n726), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n789), .B(new_n1212), .C1(new_n346), .C2(new_n826), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1191), .A2(new_n712), .B1(new_n1192), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1190), .A2(new_n1214), .ZN(G381));
  AND2_X1   g1015(.A1(new_n1017), .A2(new_n1040), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(G393), .A2(G396), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1216), .A2(new_n829), .A3(new_n1217), .ZN(new_n1218));
  OR3_X1    g1018(.A1(new_n1218), .A2(G387), .A3(G378), .ZN(new_n1219));
  OR3_X1    g1019(.A1(new_n1219), .A2(G381), .A3(G375), .ZN(G407));
  NAND2_X1  g1020(.A1(new_n639), .A2(G213), .ZN(new_n1221));
  XOR2_X1   g1021(.A(new_n1221), .B(KEYINPUT127), .Z(new_n1222));
  NAND2_X1  g1022(.A1(new_n1106), .A2(new_n1222), .ZN(new_n1223));
  OAI211_X1 g1023(.A(G407), .B(G213), .C1(G375), .C2(new_n1223), .ZN(G409));
  NAND3_X1  g1024(.A1(new_n1150), .A2(G378), .A3(new_n1185), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1109), .A2(new_n1141), .A3(new_n962), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1180), .B1(new_n1147), .B2(new_n711), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1106), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1225), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT60), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1188), .A2(new_n1230), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n661), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1214), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n829), .ZN(new_n1235));
  OAI211_X1 g1035(.A(G384), .B(new_n1214), .C1(new_n1231), .C2(new_n1233), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1229), .A2(new_n1221), .A3(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT63), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(G390), .B(new_n945), .C1(new_n964), .C2(new_n978), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1216), .A2(G387), .ZN(new_n1243));
  XOR2_X1   g1043(.A(G393), .B(G396), .Z(new_n1244));
  AND3_X1   g1044(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1244), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(new_n1245), .A2(new_n1246), .A3(KEYINPUT61), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1229), .A2(new_n1221), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n639), .A2(G213), .A3(G2897), .ZN(new_n1249));
  AND3_X1   g1049(.A1(new_n1235), .A2(new_n1236), .A3(new_n1249), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1235), .A2(new_n1236), .B1(G2897), .B2(new_n1222), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1248), .A2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1222), .B1(new_n1225), .B2(new_n1228), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1255), .A2(KEYINPUT63), .A3(new_n1238), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1241), .A2(new_n1247), .A3(new_n1254), .A4(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT61), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(new_n1255), .B2(new_n1252), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT62), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1239), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1255), .A2(KEYINPUT62), .A3(new_n1238), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1259), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1257), .B1(new_n1263), .B2(new_n1264), .ZN(G405));
  INV_X1    g1065(.A(new_n1225), .ZN(new_n1266));
  AOI21_X1  g1066(.A(G378), .B1(new_n1150), .B2(new_n1185), .ZN(new_n1267));
  OR3_X1    g1067(.A1(new_n1266), .A2(new_n1238), .A3(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1238), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1264), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1268), .A2(new_n1264), .A3(new_n1269), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(G402));
endmodule


