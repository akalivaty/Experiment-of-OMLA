//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 0 1 1 1 0 0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1333,
    new_n1334, new_n1335, new_n1336, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1395,
    new_n1396, new_n1397, new_n1398, new_n1399, new_n1400, new_n1401,
    new_n1402, new_n1403, new_n1404, new_n1405, new_n1406, new_n1407;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n202), .A2(new_n203), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n208), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT64), .Z(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n210), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n213), .B(new_n219), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G226), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XOR2_X1   g0038(.A(G50), .B(G58), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  XNOR2_X1  g0044(.A(KEYINPUT3), .B(G33), .ZN(new_n245));
  INV_X1    g0045(.A(G1698), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G222), .ZN(new_n247));
  NAND2_X1  g0047(.A1(G223), .A2(G1698), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n245), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g0049(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n250));
  OAI211_X1 g0050(.A(new_n249), .B(new_n250), .C1(G77), .C2(new_n245), .ZN(new_n251));
  INV_X1    g0051(.A(G226), .ZN(new_n252));
  INV_X1    g0052(.A(G41), .ZN(new_n253));
  INV_X1    g0053(.A(G45), .ZN(new_n254));
  AOI21_X1  g0054(.A(G1), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n251), .B1(new_n252), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G1), .A3(G13), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G274), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n262));
  NOR3_X1   g0062(.A1(new_n261), .A2(KEYINPUT66), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT66), .ZN(new_n264));
  INV_X1    g0064(.A(G274), .ZN(new_n265));
  AND2_X1   g0065(.A1(G1), .A2(G13), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n265), .B1(new_n266), .B2(new_n259), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n264), .B1(new_n267), .B2(new_n255), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n263), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n258), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(KEYINPUT10), .B1(new_n270), .B2(G190), .ZN(new_n271));
  INV_X1    g0071(.A(G13), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G1), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G20), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n201), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  AND2_X1   g0077(.A1(new_n277), .A2(new_n217), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(G1), .B2(new_n208), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT8), .B(G58), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n208), .A2(G33), .ZN(new_n281));
  INV_X1    g0081(.A(G150), .ZN(new_n282));
  INV_X1    g0082(.A(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n208), .A2(new_n283), .ZN(new_n284));
  OAI22_X1  g0084(.A1(new_n280), .A2(new_n281), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n285), .B1(G20), .B2(new_n204), .ZN(new_n286));
  OAI221_X1 g0086(.A(new_n276), .B1(new_n201), .B2(new_n279), .C1(new_n286), .C2(new_n278), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n287), .A2(KEYINPUT9), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(KEYINPUT9), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n271), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n270), .ZN(new_n292));
  AOI21_X1  g0092(.A(KEYINPUT69), .B1(new_n292), .B2(G200), .ZN(new_n293));
  AND3_X1   g0093(.A1(new_n292), .A2(KEYINPUT69), .A3(G200), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n291), .B(KEYINPUT70), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT70), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n294), .A2(new_n293), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n296), .B1(new_n297), .B2(new_n290), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n270), .A2(G190), .ZN(new_n299));
  INV_X1    g0099(.A(G200), .ZN(new_n300));
  OAI221_X1 g0100(.A(new_n299), .B1(new_n300), .B2(new_n270), .C1(new_n288), .C2(new_n289), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n295), .A2(new_n298), .B1(KEYINPUT10), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G179), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n270), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n304), .B(new_n287), .C1(G169), .C2(new_n270), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  OR2_X1    g0107(.A1(KEYINPUT3), .A2(G33), .ZN(new_n308));
  NAND2_X1  g0108(.A1(KEYINPUT3), .A2(G33), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n308), .A2(new_n208), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT7), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n308), .A2(KEYINPUT7), .A3(new_n208), .A4(new_n309), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G68), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT72), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G58), .A2(G68), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n208), .B1(new_n214), .B2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(G20), .A2(G33), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G159), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n316), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n317), .ZN(new_n323));
  NOR2_X1   g0123(.A1(G58), .A2(G68), .ZN(new_n324));
  OAI21_X1  g0124(.A(G20), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n325), .A2(KEYINPUT72), .A3(new_n320), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n315), .A2(new_n327), .A3(KEYINPUT16), .ZN(new_n328));
  INV_X1    g0128(.A(new_n278), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT16), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n203), .B1(new_n312), .B2(new_n313), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n325), .A2(new_n320), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n328), .A2(new_n329), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n280), .B1(new_n207), .B2(G20), .ZN(new_n335));
  AOI211_X1 g0135(.A(new_n275), .B(new_n329), .C1(new_n335), .C2(KEYINPUT73), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n335), .A2(KEYINPUT73), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n336), .A2(new_n338), .B1(new_n275), .B2(new_n280), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  AND3_X1   g0140(.A1(new_n260), .A2(G232), .A3(new_n262), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n252), .A2(G1698), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(G223), .B2(G1698), .ZN(new_n343));
  AND2_X1   g0143(.A1(KEYINPUT3), .A2(G33), .ZN(new_n344));
  NOR2_X1   g0144(.A1(KEYINPUT3), .A2(G33), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G87), .ZN(new_n347));
  OAI22_X1  g0147(.A1(new_n343), .A2(new_n346), .B1(new_n283), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n341), .B1(new_n348), .B2(new_n250), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT66), .B1(new_n261), .B2(new_n262), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n267), .A2(new_n264), .A3(new_n255), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AND3_X1   g0152(.A1(new_n349), .A2(G179), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G169), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n354), .B1(new_n349), .B2(new_n352), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT74), .ZN(new_n356));
  NOR3_X1   g0156(.A1(new_n353), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n341), .ZN(new_n358));
  NOR2_X1   g0158(.A1(G223), .A2(G1698), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n359), .B1(new_n252), .B2(G1698), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n360), .A2(new_n245), .B1(G33), .B2(G87), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n358), .B1(new_n361), .B2(new_n260), .ZN(new_n362));
  OAI21_X1  g0162(.A(G169), .B1(new_n362), .B2(new_n269), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n349), .A2(G179), .A3(new_n352), .ZN(new_n364));
  AOI21_X1  g0164(.A(KEYINPUT74), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n340), .B1(new_n357), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT18), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n356), .B1(new_n353), .B2(new_n355), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n363), .A2(KEYINPUT74), .A3(new_n364), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n371), .A2(KEYINPUT18), .A3(new_n340), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n335), .A2(KEYINPUT73), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n373), .A2(new_n274), .A3(new_n278), .ZN(new_n374));
  INV_X1    g0174(.A(new_n280), .ZN(new_n375));
  OAI22_X1  g0175(.A1(new_n374), .A2(new_n337), .B1(new_n274), .B2(new_n375), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n314), .A2(G68), .B1(new_n322), .B2(new_n326), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n278), .B1(new_n377), .B2(KEYINPUT16), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n376), .B1(new_n378), .B2(new_n333), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT75), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT17), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n300), .B1(new_n362), .B2(new_n269), .ZN(new_n382));
  INV_X1    g0182(.A(G190), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n349), .A2(new_n383), .A3(new_n352), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n379), .A2(new_n380), .A3(new_n381), .A4(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n385), .A2(new_n380), .A3(new_n334), .A4(new_n339), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT17), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n368), .A2(new_n372), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n319), .A2(G50), .ZN(new_n390));
  XNOR2_X1  g0190(.A(new_n390), .B(KEYINPUT71), .ZN(new_n391));
  INV_X1    g0191(.A(G77), .ZN(new_n392));
  OAI22_X1  g0192(.A1(new_n281), .A2(new_n392), .B1(new_n208), .B2(G68), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n329), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT11), .ZN(new_n395));
  OR2_X1    g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n394), .A2(new_n395), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n203), .B1(new_n279), .B2(KEYINPUT12), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n275), .A2(KEYINPUT12), .ZN(new_n399));
  AND4_X1   g0199(.A1(KEYINPUT12), .A2(new_n273), .A3(G20), .A4(new_n203), .ZN(new_n400));
  NOR3_X1   g0200(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n396), .A2(new_n397), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(G232), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(G1698), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(G226), .B2(G1698), .ZN(new_n405));
  INV_X1    g0205(.A(G97), .ZN(new_n406));
  OAI22_X1  g0206(.A1(new_n405), .A2(new_n346), .B1(new_n283), .B2(new_n406), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n407), .A2(new_n250), .B1(G238), .B2(new_n256), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n352), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(KEYINPUT13), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT13), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n408), .A2(new_n411), .A3(new_n352), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT14), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(new_n414), .A3(G169), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n303), .B2(new_n413), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n414), .B1(new_n413), .B2(G169), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n402), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n402), .B1(new_n413), .B2(G200), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n383), .B2(new_n413), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(G238), .A2(G1698), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n245), .B(new_n422), .C1(new_n403), .C2(G1698), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n423), .B(new_n250), .C1(G107), .C2(new_n245), .ZN(new_n424));
  INV_X1    g0224(.A(G244), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n424), .B1(new_n425), .B2(new_n257), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n426), .A2(new_n269), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n303), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n428), .B1(G169), .B2(new_n427), .ZN(new_n429));
  XNOR2_X1  g0229(.A(KEYINPUT15), .B(G87), .ZN(new_n430));
  OAI22_X1  g0230(.A1(new_n430), .A2(new_n281), .B1(new_n208), .B2(new_n392), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n280), .A2(new_n284), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n329), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  XNOR2_X1  g0233(.A(new_n433), .B(KEYINPUT67), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n275), .A2(new_n392), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(new_n279), .B2(new_n392), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  OR2_X1    g0237(.A1(new_n429), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(G200), .B1(new_n426), .B2(new_n269), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n437), .A2(KEYINPUT68), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n427), .A2(G190), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(KEYINPUT68), .B1(new_n437), .B2(new_n440), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n439), .A2(new_n445), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n421), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n307), .A2(new_n389), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT76), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n307), .A2(new_n447), .A3(KEYINPUT76), .A4(new_n389), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(G107), .ZN(new_n454));
  AND3_X1   g0254(.A1(new_n454), .A2(KEYINPUT23), .A3(G20), .ZN(new_n455));
  AOI21_X1  g0255(.A(KEYINPUT23), .B1(new_n454), .B2(G20), .ZN(new_n456));
  INV_X1    g0256(.A(G116), .ZN(new_n457));
  OAI22_X1  g0257(.A1(new_n455), .A2(new_n456), .B1(new_n457), .B2(new_n281), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n208), .B(G87), .C1(new_n344), .C2(new_n345), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT22), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT22), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n245), .A2(new_n461), .A3(new_n208), .A4(G87), .ZN(new_n462));
  AOI211_X1 g0262(.A(KEYINPUT24), .B(new_n458), .C1(new_n460), .C2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT24), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n460), .A2(new_n462), .ZN(new_n465));
  INV_X1    g0265(.A(new_n458), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n329), .B1(new_n463), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT82), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g0270(.A(KEYINPUT82), .B(new_n329), .C1(new_n463), .C2(new_n467), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n275), .A2(KEYINPUT25), .A3(new_n454), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT25), .B1(new_n275), .B2(new_n454), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n207), .A2(G33), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n278), .A2(new_n274), .A3(new_n476), .ZN(new_n477));
  OAI22_X1  g0277(.A1(new_n474), .A2(new_n475), .B1(new_n477), .B2(new_n454), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT83), .ZN(new_n480));
  INV_X1    g0280(.A(G250), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n481), .B1(new_n308), .B2(new_n309), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n482), .A2(new_n246), .B1(G33), .B2(G294), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n245), .A2(G257), .A3(G1698), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n260), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT5), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G41), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n253), .A2(KEYINPUT5), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n254), .A2(G1), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n267), .A2(new_n487), .A3(new_n488), .A4(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n489), .A2(new_n487), .A3(new_n488), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(G264), .A3(new_n260), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n480), .B1(new_n485), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n245), .A2(G250), .A3(new_n246), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G33), .A2(G294), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n484), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n250), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n498), .A2(KEYINPUT83), .A3(new_n490), .A4(new_n492), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n494), .A2(new_n499), .A3(new_n383), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n492), .A2(KEYINPUT84), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT84), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n491), .A2(new_n502), .A3(G264), .A4(new_n260), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n504), .A2(new_n498), .A3(new_n490), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n300), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n472), .A2(new_n479), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n494), .A2(new_n499), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G169), .ZN(new_n510));
  OR2_X1    g0310(.A1(new_n505), .A2(new_n303), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n472), .A2(new_n479), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n277), .A2(new_n217), .B1(G20), .B2(new_n457), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G283), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n515), .B(new_n208), .C1(G33), .C2(new_n406), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n514), .A2(KEYINPUT20), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT20), .B1(new_n514), .B2(new_n516), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n275), .A2(new_n457), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(new_n477), .B2(new_n457), .ZN(new_n521));
  OAI21_X1  g0321(.A(G169), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT79), .ZN(new_n524));
  AND2_X1   g0324(.A1(G264), .A2(G1698), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n524), .B1(new_n245), .B2(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n524), .B(new_n525), .C1(new_n344), .C2(new_n345), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n245), .A2(G257), .ZN(new_n530));
  INV_X1    g0330(.A(G303), .ZN(new_n531));
  OAI22_X1  g0331(.A1(new_n530), .A2(G1698), .B1(new_n531), .B2(new_n245), .ZN(new_n532));
  OAI21_X1  g0332(.A(KEYINPUT80), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n525), .B1(new_n344), .B2(new_n345), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT79), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n527), .ZN(new_n536));
  INV_X1    g0336(.A(G257), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n537), .B1(new_n308), .B2(new_n309), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n538), .A2(new_n246), .B1(new_n346), .B2(G303), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT80), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n536), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n260), .B1(new_n533), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n491), .A2(G270), .A3(new_n260), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n490), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n523), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT21), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n536), .A2(new_n539), .A3(new_n540), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n540), .B1(new_n536), .B2(new_n539), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n250), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n544), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT21), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n551), .A2(new_n552), .A3(new_n523), .ZN(new_n553));
  INV_X1    g0353(.A(new_n551), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n519), .A2(new_n521), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n555), .A2(new_n303), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n546), .A2(new_n553), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(G200), .B1(new_n542), .B2(new_n544), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n549), .A2(G190), .A3(new_n550), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n558), .A2(new_n555), .A3(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT81), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n555), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n563), .B1(new_n551), .B2(G200), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n564), .A2(KEYINPUT81), .A3(new_n559), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n454), .A2(KEYINPUT6), .A3(G97), .ZN(new_n567));
  XNOR2_X1  g0367(.A(G97), .B(G107), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT6), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI22_X1  g0370(.A1(new_n570), .A2(new_n208), .B1(new_n392), .B2(new_n284), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n454), .B1(new_n312), .B2(new_n313), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n329), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n274), .A2(G97), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n477), .B2(new_n406), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT4), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n579), .A2(G1698), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n580), .B(G244), .C1(new_n345), .C2(new_n344), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n425), .B1(new_n308), .B2(new_n309), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n581), .B(new_n515), .C1(new_n582), .C2(KEYINPUT4), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n245), .A2(G250), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n246), .B1(new_n584), .B2(KEYINPUT4), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n250), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n491), .A2(G257), .A3(new_n260), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n490), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n586), .A2(new_n303), .A3(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(G1698), .B1(new_n482), .B2(new_n579), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n579), .B1(new_n346), .B2(new_n425), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n591), .A2(new_n515), .A3(new_n592), .A4(new_n581), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n588), .B1(new_n593), .B2(new_n250), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n578), .B(new_n590), .C1(G169), .C2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT78), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n283), .A2(new_n457), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  OR2_X1    g0398(.A1(G238), .A2(G1698), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n425), .A2(G1698), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n598), .B1(new_n601), .B2(new_n346), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n250), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n481), .B1(new_n207), .B2(G45), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n260), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT77), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n604), .A2(new_n260), .A3(KEYINPUT77), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n267), .A2(new_n489), .ZN(new_n610));
  AND4_X1   g0410(.A1(new_n596), .A2(new_n603), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n260), .A2(G274), .A3(new_n489), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n612), .B1(new_n602), .B2(new_n250), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n596), .B1(new_n613), .B2(new_n609), .ZN(new_n614));
  OAI21_X1  g0414(.A(G200), .B1(new_n611), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n208), .B1(new_n283), .B2(new_n406), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n347), .A2(new_n406), .A3(new_n454), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(KEYINPUT19), .A3(new_n617), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n208), .B(G68), .C1(new_n344), .C2(new_n345), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT19), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(new_n281), .B2(new_n406), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n618), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n329), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n278), .A2(new_n274), .A3(G87), .A4(new_n476), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n275), .A2(new_n430), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(G238), .A2(G1698), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(new_n425), .B2(G1698), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n597), .B1(new_n629), .B2(new_n245), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n610), .B1(new_n630), .B2(new_n260), .ZN(new_n631));
  INV_X1    g0431(.A(new_n608), .ZN(new_n632));
  AOI21_X1  g0432(.A(KEYINPUT77), .B1(new_n604), .B2(new_n260), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(KEYINPUT78), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n613), .A2(new_n596), .A3(new_n609), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(G190), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n615), .A2(new_n627), .A3(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n354), .B1(new_n611), .B2(new_n614), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n635), .A2(new_n303), .A3(new_n636), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n623), .B(new_n625), .C1(new_n430), .C2(new_n477), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT7), .B1(new_n346), .B2(new_n208), .ZN(new_n643));
  INV_X1    g0443(.A(new_n313), .ZN(new_n644));
  OAI21_X1  g0444(.A(G107), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n284), .A2(new_n392), .ZN(new_n646));
  AND2_X1   g0446(.A1(G97), .A2(G107), .ZN(new_n647));
  NOR2_X1   g0447(.A1(G97), .A2(G107), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n569), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n454), .A2(KEYINPUT6), .A3(G97), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n646), .B1(new_n651), .B2(G20), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n645), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n576), .B1(new_n653), .B2(new_n329), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n586), .A2(G190), .A3(new_n589), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n654), .B(new_n655), .C1(new_n300), .C2(new_n594), .ZN(new_n656));
  AND4_X1   g0456(.A1(new_n595), .A2(new_n638), .A3(new_n642), .A4(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n513), .A2(new_n557), .A3(new_n566), .A4(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n453), .A2(new_n658), .ZN(G372));
  NAND2_X1  g0459(.A1(new_n363), .A2(new_n364), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n340), .A2(new_n367), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n367), .B1(new_n340), .B2(new_n660), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n418), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n664), .B1(new_n420), .B2(new_n439), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n386), .A2(new_n388), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n663), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n295), .A2(new_n298), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n301), .A2(KEYINPUT10), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n306), .B1(new_n668), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n354), .B1(new_n631), .B2(new_n634), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n640), .A2(new_n641), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT26), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n300), .B1(new_n613), .B2(new_n609), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(new_n626), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n637), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n676), .B1(new_n680), .B2(new_n595), .ZN(new_n681));
  INV_X1    g0481(.A(new_n595), .ZN(new_n682));
  XOR2_X1   g0482(.A(KEYINPUT86), .B(KEYINPUT26), .Z(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n682), .A2(new_n642), .A3(new_n638), .A4(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n675), .B1(new_n681), .B2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT85), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n554), .A2(new_n556), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n552), .B1(new_n551), .B2(new_n523), .ZN(new_n690));
  AOI211_X1 g0490(.A(KEYINPUT21), .B(new_n522), .C1(new_n549), .C2(new_n550), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(new_n512), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n472), .A2(new_n479), .A3(new_n507), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n674), .A2(new_n679), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n595), .A2(new_n656), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n688), .B1(new_n693), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n465), .A2(new_n466), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT24), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n465), .A2(new_n464), .A3(new_n466), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(KEYINPUT82), .B1(new_n702), .B2(new_n329), .ZN(new_n703));
  INV_X1    g0503(.A(new_n471), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n479), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n510), .A2(new_n511), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n557), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n674), .A2(new_n595), .A3(new_n656), .A4(new_n679), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n478), .B1(new_n470), .B2(new_n471), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n709), .B1(new_n710), .B2(new_n507), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n708), .A2(new_n711), .A3(KEYINPUT85), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n687), .B1(new_n698), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n672), .B1(new_n453), .B2(new_n713), .ZN(G369));
  INV_X1    g0514(.A(new_n273), .ZN(new_n715));
  OR3_X1    g0515(.A1(new_n715), .A2(KEYINPUT27), .A3(G20), .ZN(new_n716));
  OAI21_X1  g0516(.A(KEYINPUT27), .B1(new_n715), .B2(G20), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n716), .A2(G213), .A3(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(G343), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n557), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n720), .ZN(new_n722));
  OR3_X1    g0522(.A1(new_n710), .A2(KEYINPUT87), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(KEYINPUT87), .B1(new_n710), .B2(new_n722), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n721), .A2(new_n513), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  XOR2_X1   g0525(.A(new_n720), .B(KEYINPUT88), .Z(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n512), .A2(new_n727), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n729), .A2(KEYINPUT89), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(KEYINPUT89), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n692), .B1(new_n562), .B2(new_n565), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n563), .A2(new_n720), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n735), .B1(new_n557), .B2(new_n734), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G330), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n513), .A2(new_n723), .A3(new_n724), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n739), .B1(new_n707), .B2(new_n722), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n732), .A2(new_n741), .ZN(G399));
  NAND2_X1  g0542(.A1(new_n211), .A2(new_n253), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n617), .A2(G116), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n743), .A2(G1), .A3(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n745), .B1(new_n215), .B2(new_n743), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT28), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT94), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n748), .B1(new_n658), .B2(new_n726), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n638), .A2(new_n642), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n707), .A2(new_n750), .A3(new_n694), .A4(new_n696), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n752), .A2(KEYINPUT94), .A3(new_n733), .A4(new_n727), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n611), .A2(new_n614), .ZN(new_n755));
  AND3_X1   g0555(.A1(new_n586), .A2(KEYINPUT30), .A3(new_n589), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n544), .A2(new_n303), .ZN(new_n757));
  AND3_X1   g0557(.A1(new_n757), .A2(new_n498), .A3(new_n504), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n755), .A2(new_n756), .A3(new_n758), .A4(new_n549), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT92), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n757), .A2(new_n498), .A3(new_n504), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n762), .A2(new_n611), .A3(new_n614), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n763), .A2(KEYINPUT92), .A3(new_n549), .A4(new_n756), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n755), .A2(new_n549), .A3(new_n758), .A4(new_n594), .ZN(new_n766));
  XOR2_X1   g0566(.A(KEYINPUT91), .B(KEYINPUT30), .Z(new_n767));
  AOI21_X1  g0567(.A(G179), .B1(new_n613), .B2(new_n609), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n505), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n594), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n766), .A2(new_n767), .B1(new_n770), .B2(new_n551), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n765), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(new_n720), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT93), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT31), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n722), .B1(new_n765), .B2(new_n771), .ZN(new_n777));
  OAI21_X1  g0577(.A(KEYINPUT93), .B1(new_n777), .B2(KEYINPUT31), .ZN(new_n778));
  XOR2_X1   g0578(.A(KEYINPUT90), .B(KEYINPUT31), .Z(new_n779));
  NOR2_X1   g0579(.A1(new_n727), .A2(new_n779), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n776), .A2(new_n778), .B1(new_n772), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n754), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G330), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n675), .B1(new_n708), .B2(new_n711), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n750), .A2(new_n682), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(new_n683), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n695), .A2(KEYINPUT26), .A3(new_n682), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n720), .B1(new_n784), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(KEYINPUT29), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n713), .A2(new_n726), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n790), .B1(new_n791), .B2(KEYINPUT29), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n783), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n747), .B1(new_n794), .B2(G1), .ZN(G364));
  NOR2_X1   g0595(.A1(new_n272), .A2(G20), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G45), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n743), .A2(G1), .A3(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n738), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(G330), .B2(new_n736), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n211), .A2(new_n245), .ZN(new_n802));
  INV_X1    g0602(.A(G355), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n802), .A2(new_n803), .B1(G116), .B2(new_n211), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n240), .A2(G45), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n211), .A2(new_n346), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(new_n254), .B2(new_n216), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n804), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(G13), .A2(G33), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(G20), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n217), .B1(G20), .B2(new_n354), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n799), .B1(new_n808), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n208), .A2(new_n383), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n816), .A2(new_n303), .A3(G200), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n303), .A2(G200), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n817), .A2(new_n347), .B1(new_n819), .B2(new_n202), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n208), .A2(G190), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n346), .B(new_n820), .C1(G77), .C2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(G179), .A2(G200), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n821), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(G159), .ZN(new_n828));
  OR2_X1    g0628(.A1(new_n828), .A2(KEYINPUT32), .ZN(new_n829));
  NAND3_X1  g0629(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(new_n383), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n828), .A2(KEYINPUT32), .B1(new_n831), .B2(G50), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n821), .A2(new_n303), .A3(G200), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT95), .Z(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(G107), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n824), .A2(new_n829), .A3(new_n832), .A4(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n208), .B1(new_n825), .B2(G190), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n837), .A2(new_n406), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n830), .A2(G190), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n838), .B1(new_n839), .B2(G68), .ZN(new_n840));
  XOR2_X1   g0640(.A(new_n840), .B(KEYINPUT96), .Z(new_n841));
  INV_X1    g0641(.A(new_n819), .ZN(new_n842));
  XNOR2_X1  g0642(.A(KEYINPUT33), .B(G317), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n842), .A2(G322), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT97), .Z(new_n845));
  NAND2_X1  g0645(.A1(new_n834), .A2(G283), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n245), .B1(new_n823), .B2(G311), .ZN(new_n847));
  INV_X1    g0647(.A(new_n817), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n848), .A2(G303), .B1(new_n827), .B2(G329), .ZN(new_n849));
  INV_X1    g0649(.A(new_n837), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n850), .A2(G294), .B1(G326), .B2(new_n831), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n846), .A2(new_n847), .A3(new_n849), .A4(new_n851), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n836), .A2(new_n841), .B1(new_n845), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n815), .B1(new_n853), .B2(new_n812), .ZN(new_n854));
  INV_X1    g0654(.A(new_n811), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n854), .B1(new_n736), .B2(new_n855), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n801), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(G396));
  INV_X1    g0658(.A(KEYINPUT98), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n438), .A2(new_n720), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n443), .A2(new_n444), .B1(new_n437), .B2(new_n722), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n860), .B1(new_n861), .B2(new_n438), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n791), .B(new_n862), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(new_n783), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n798), .ZN(new_n865));
  INV_X1    g0665(.A(new_n862), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n809), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n834), .A2(G87), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n245), .B(new_n838), .C1(G311), .C2(new_n827), .ZN(new_n869));
  AOI22_X1  g0669(.A1(G283), .A2(new_n839), .B1(new_n831), .B2(G303), .ZN(new_n870));
  INV_X1    g0670(.A(G294), .ZN(new_n871));
  OAI22_X1  g0671(.A1(new_n819), .A2(new_n871), .B1(new_n822), .B2(new_n457), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(G107), .B2(new_n848), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n868), .A2(new_n869), .A3(new_n870), .A4(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(G132), .ZN(new_n875));
  OAI221_X1 g0675(.A(new_n245), .B1(new_n826), .B2(new_n875), .C1(new_n817), .C2(new_n201), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(G58), .B2(new_n850), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n834), .A2(G68), .ZN(new_n878));
  AOI22_X1  g0678(.A1(G143), .A2(new_n842), .B1(new_n823), .B2(G159), .ZN(new_n879));
  INV_X1    g0679(.A(new_n839), .ZN(new_n880));
  INV_X1    g0680(.A(G137), .ZN(new_n881));
  INV_X1    g0681(.A(new_n831), .ZN(new_n882));
  OAI221_X1 g0682(.A(new_n879), .B1(new_n880), .B2(new_n282), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT34), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n877), .B(new_n878), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n883), .A2(new_n884), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n874), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n812), .A2(new_n809), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n887), .A2(new_n812), .B1(new_n392), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n798), .B1(new_n867), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n859), .B1(new_n865), .B2(new_n891), .ZN(new_n892));
  AOI211_X1 g0692(.A(KEYINPUT98), .B(new_n890), .C1(new_n864), .C2(new_n798), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(G384));
  OR2_X1    g0695(.A1(new_n651), .A2(KEYINPUT35), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n651), .A2(KEYINPUT35), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n896), .A2(new_n897), .A3(G116), .A4(new_n218), .ZN(new_n898));
  XOR2_X1   g0698(.A(new_n898), .B(KEYINPUT36), .Z(new_n899));
  NAND3_X1  g0699(.A1(new_n216), .A2(G77), .A3(new_n317), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n201), .A2(G68), .ZN(new_n901));
  AOI211_X1 g0701(.A(new_n207), .B(G13), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n402), .A2(new_n720), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n418), .A2(new_n420), .A3(new_n904), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n402), .B(new_n720), .C1(new_n416), .C2(new_n417), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT38), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n328), .A2(new_n329), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n377), .A2(KEYINPUT16), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n339), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n718), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n368), .A2(new_n372), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n914), .B1(new_n915), .B2(new_n666), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n385), .A2(new_n339), .A3(new_n334), .ZN(new_n917));
  INV_X1    g0717(.A(new_n660), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n315), .A2(new_n327), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n330), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n376), .B1(new_n378), .B2(new_n920), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n914), .B(new_n917), .C1(new_n918), .C2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n340), .B1(new_n371), .B2(new_n913), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT37), .B1(new_n379), .B2(new_n385), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n922), .A2(KEYINPUT37), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n909), .B1(new_n916), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n917), .B1(new_n921), .B2(new_n918), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n921), .A2(new_n718), .ZN(new_n928));
  OAI21_X1  g0728(.A(KEYINPUT37), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n923), .A2(new_n924), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n931), .B(KEYINPUT38), .C1(new_n389), .C2(new_n914), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n926), .A2(new_n932), .ZN(new_n933));
  NOR3_X1   g0733(.A1(new_n693), .A2(new_n688), .A3(new_n697), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT85), .B1(new_n708), .B2(new_n711), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n686), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n936), .A2(new_n727), .A3(new_n862), .ZN(new_n937));
  INV_X1    g0737(.A(new_n860), .ZN(new_n938));
  AOI211_X1 g0738(.A(new_n908), .B(new_n933), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n664), .A2(new_n722), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n340), .A2(new_n913), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n663), .B2(new_n666), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n942), .B(new_n917), .C1(new_n379), .C2(new_n918), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n944), .A2(KEYINPUT37), .B1(new_n923), .B2(new_n924), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n909), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT39), .ZN(new_n947));
  AND3_X1   g0747(.A1(new_n932), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n947), .B1(new_n926), .B2(new_n932), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n941), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n663), .A2(new_n913), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(KEYINPUT99), .B1(new_n939), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n937), .A2(new_n938), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n926), .A2(new_n932), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n955), .A2(new_n956), .A3(new_n907), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT99), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n957), .A2(new_n958), .A3(new_n950), .A4(new_n952), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n954), .A2(new_n959), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n452), .B(new_n790), .C1(KEYINPUT29), .C2(new_n791), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n672), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n960), .B(new_n962), .Z(new_n963));
  INV_X1    g0763(.A(G330), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n862), .A2(new_n907), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(KEYINPUT81), .B1(new_n564), .B2(new_n559), .ZN(new_n967));
  AND4_X1   g0767(.A1(KEYINPUT81), .A2(new_n558), .A3(new_n555), .A4(new_n559), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n557), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n969), .A2(new_n751), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT94), .B1(new_n970), .B2(new_n727), .ZN(new_n971));
  NOR4_X1   g0771(.A1(new_n969), .A2(new_n751), .A3(new_n748), .A4(new_n726), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT101), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n777), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n779), .B1(new_n777), .B2(new_n974), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n976), .A2(new_n977), .B1(new_n775), .B2(new_n773), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n956), .B(new_n966), .C1(new_n973), .C2(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(KEYINPUT100), .B(KEYINPUT40), .Z(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n773), .A2(new_n775), .ZN(new_n983));
  INV_X1    g0783(.A(new_n779), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(new_n773), .B2(KEYINPUT101), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n983), .B1(new_n985), .B2(new_n975), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n754), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n932), .A2(new_n946), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n988), .A2(KEYINPUT40), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n987), .A2(new_n989), .A3(new_n966), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n982), .A2(new_n990), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n452), .A2(new_n987), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n964), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n991), .B2(new_n992), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n963), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n207), .B2(new_n796), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n963), .A2(new_n994), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n903), .B1(new_n996), .B2(new_n997), .ZN(G367));
  NOR2_X1   g0798(.A1(new_n722), .A2(new_n627), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n675), .A2(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT102), .Z(new_n1001));
  NOR2_X1   g0801(.A1(new_n680), .A2(new_n999), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT103), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1005), .A2(KEYINPUT43), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n741), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n696), .B1(new_n727), .B2(new_n654), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT104), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(new_n682), .B2(new_n726), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1008), .A2(new_n1013), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1014), .A2(KEYINPUT106), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(KEYINPUT106), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1007), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1005), .A2(KEYINPUT43), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1012), .A2(new_n725), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT105), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1020), .B(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT42), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1020), .B(KEYINPUT105), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(KEYINPUT42), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n682), .B1(new_n1011), .B2(new_n512), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1024), .B(new_n1026), .C1(new_n726), .C2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1015), .A2(new_n1007), .A3(new_n1016), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1018), .A2(new_n1019), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1028), .A2(new_n1019), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1029), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1031), .B1(new_n1032), .B2(new_n1017), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n743), .B(KEYINPUT41), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n740), .A2(new_n721), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n725), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n738), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1037), .A2(new_n737), .A3(new_n725), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n794), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT108), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1042), .B(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(KEYINPUT44), .B1(new_n732), .B2(new_n1013), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT44), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n730), .A2(new_n1046), .A3(new_n731), .A4(new_n1012), .ZN(new_n1047));
  AOI21_X1  g0847(.A(KEYINPUT45), .B1(new_n732), .B2(new_n1013), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT45), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n1049), .B(new_n1012), .C1(new_n730), .C2(new_n731), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1045), .B(new_n1047), .C1(new_n1048), .C2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT107), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1051), .A2(new_n1052), .A3(new_n741), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n741), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1044), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1036), .B1(new_n1056), .B2(new_n794), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n797), .A2(G1), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1035), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1004), .A2(new_n811), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n236), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n813), .B1(new_n211), .B2(new_n430), .C1(new_n1061), .C2(new_n806), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n799), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n837), .A2(new_n203), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1065), .B(new_n245), .C1(new_n282), .C2(new_n819), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n817), .A2(new_n202), .B1(new_n822), .B2(new_n201), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n833), .A2(new_n392), .B1(new_n826), .B2(new_n881), .ZN(new_n1068));
  INV_X1    g0868(.A(G159), .ZN(new_n1069));
  INV_X1    g0869(.A(G143), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n880), .A2(new_n1069), .B1(new_n882), .B2(new_n1070), .ZN(new_n1071));
  NOR4_X1   g0871(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .A4(new_n1071), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT109), .Z(new_n1073));
  NOR2_X1   g0873(.A1(new_n817), .A2(new_n457), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1074), .A2(KEYINPUT46), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(G107), .B2(new_n850), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1074), .A2(KEYINPUT46), .B1(new_n831), .B2(G311), .ZN(new_n1077));
  INV_X1    g0877(.A(G283), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n833), .A2(new_n406), .B1(new_n822), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(G317), .B2(new_n827), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n346), .B1(new_n819), .B2(new_n531), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(G294), .B2(new_n839), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1076), .A2(new_n1077), .A3(new_n1080), .A4(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1073), .A2(new_n1083), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT47), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1063), .B1(new_n1085), .B2(new_n812), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1060), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1059), .A2(new_n1087), .ZN(G387));
  XNOR2_X1  g0888(.A(new_n1042), .B(KEYINPUT108), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n743), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n793), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  OR2_X1    g0892(.A1(new_n740), .A2(new_n855), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n802), .A2(new_n744), .B1(G107), .B2(new_n211), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n233), .A2(G45), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n744), .ZN(new_n1096));
  AOI211_X1 g0896(.A(G45), .B(new_n1096), .C1(G68), .C2(G77), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n280), .A2(G50), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT50), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n806), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1094), .B1(new_n1095), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n799), .B1(new_n1101), .B2(new_n814), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n834), .A2(G97), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n837), .A2(new_n430), .ZN(new_n1104));
  XOR2_X1   g0904(.A(KEYINPUT110), .B(G150), .Z(new_n1105));
  AOI211_X1 g0905(.A(new_n346), .B(new_n1104), .C1(new_n827), .C2(new_n1105), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n375), .A2(new_n839), .B1(G159), .B2(new_n831), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n817), .A2(new_n392), .B1(new_n822), .B2(new_n203), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(G50), .B2(new_n842), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1103), .A2(new_n1106), .A3(new_n1107), .A4(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n245), .B1(new_n827), .B2(G326), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n817), .A2(new_n871), .B1(new_n837), .B2(new_n1078), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT111), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(G317), .A2(new_n842), .B1(new_n823), .B2(G303), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n839), .A2(G311), .ZN(new_n1115));
  INV_X1    g0915(.A(G322), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1114), .B(new_n1115), .C1(new_n1116), .C2(new_n882), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT48), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1113), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n1118), .B2(new_n1117), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT49), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n1111), .B1(new_n457), .B2(new_n833), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1110), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1102), .B1(new_n1124), .B2(new_n812), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n1041), .A2(new_n1058), .B1(new_n1093), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1092), .A2(new_n1126), .ZN(G393));
  NAND2_X1  g0927(.A1(new_n732), .A2(new_n1013), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n1049), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n732), .A2(KEYINPUT45), .A3(new_n1013), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1131), .A2(new_n741), .A3(new_n1045), .A4(new_n1047), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1051), .A2(new_n1008), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT114), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n1134), .A2(new_n1135), .A3(new_n1089), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1135), .B1(new_n1134), .B2(new_n1089), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1090), .B(new_n1056), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1132), .A2(new_n1133), .A3(new_n1058), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n813), .B1(new_n406), .B2(new_n211), .C1(new_n243), .C2(new_n806), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n798), .B1(new_n1140), .B2(KEYINPUT112), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(KEYINPUT112), .B2(new_n1140), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n822), .A2(new_n280), .B1(new_n826), .B2(new_n1070), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n346), .B(new_n1143), .C1(G68), .C2(new_n848), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n882), .A2(new_n282), .B1(new_n819), .B2(new_n1069), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT51), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n837), .A2(new_n392), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(new_n839), .B2(G50), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1144), .A2(new_n1146), .A3(new_n868), .A4(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n245), .B1(new_n827), .B2(G322), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n835), .B(new_n1150), .C1(new_n1078), .C2(new_n817), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT113), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n842), .A2(G311), .B1(G317), .B2(new_n831), .ZN(new_n1153));
  XOR2_X1   g0953(.A(new_n1153), .B(KEYINPUT52), .Z(new_n1154));
  AOI22_X1  g0954(.A1(new_n823), .A2(G294), .B1(G303), .B2(new_n839), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1154), .B(new_n1155), .C1(new_n457), .C2(new_n837), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1149), .B1(new_n1152), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1142), .B1(new_n1157), .B2(new_n812), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n1013), .B2(new_n855), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1139), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1138), .A2(new_n1161), .ZN(G390));
  AOI21_X1  g0962(.A(new_n964), .B1(new_n754), .B2(new_n986), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n452), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n961), .A2(new_n672), .A3(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n782), .A2(G330), .A3(new_n966), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n861), .A2(new_n438), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n860), .B1(new_n789), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n907), .B1(new_n1163), .B2(new_n862), .ZN(new_n1170));
  OAI21_X1  g0970(.A(KEYINPUT115), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  OAI211_X1 g0971(.A(G330), .B(new_n862), .C1(new_n973), .C2(new_n978), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n908), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n789), .A2(new_n1167), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n938), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n964), .B1(new_n754), .B2(new_n781), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1175), .B1(new_n1176), .B2(new_n966), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT115), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1173), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1171), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1163), .A2(new_n966), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n907), .B1(new_n1176), .B2(new_n862), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n955), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1165), .B1(new_n1180), .B2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n948), .A2(new_n949), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n908), .B1(new_n937), .B2(new_n938), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1186), .B1(new_n1187), .B2(new_n941), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n940), .B(new_n988), .C1(new_n1168), .C2(new_n908), .ZN(new_n1189));
  AND3_X1   g0989(.A1(new_n1188), .A2(new_n1166), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1181), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(KEYINPUT116), .B1(new_n1185), .B2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n743), .B1(new_n1185), .B2(new_n1192), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n1173), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1178), .B1(new_n1173), .B2(new_n1177), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1184), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1165), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT116), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1188), .A2(new_n1166), .A3(new_n1189), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1201), .B1(new_n1202), .B2(new_n1181), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1199), .A2(new_n1200), .A3(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1193), .A2(new_n1194), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1186), .A2(new_n809), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n812), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n848), .A2(new_n1105), .ZN(new_n1208));
  XOR2_X1   g1008(.A(new_n1208), .B(KEYINPUT53), .Z(new_n1209));
  INV_X1    g1009(.A(G125), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n245), .B1(new_n826), .B2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(G159), .B2(new_n850), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G128), .A2(new_n831), .B1(new_n839), .B2(G137), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(KEYINPUT54), .B(G143), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n833), .A2(new_n201), .B1(new_n822), .B2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G132), .B2(new_n842), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1209), .A2(new_n1212), .A3(new_n1213), .A4(new_n1216), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n245), .B(new_n1147), .C1(G87), .C2(new_n848), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G107), .A2(new_n839), .B1(new_n831), .B2(G283), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n819), .A2(new_n457), .B1(new_n826), .B2(new_n871), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(G97), .B2(new_n823), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n878), .A2(new_n1218), .A3(new_n1219), .A4(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1207), .B1(new_n1217), .B2(new_n1222), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n798), .B(new_n1223), .C1(new_n280), .C2(new_n888), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1192), .A2(new_n1058), .B1(new_n1206), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1205), .A2(new_n1225), .ZN(G378));
  OAI22_X1  g1026(.A1(new_n882), .A2(new_n1210), .B1(new_n837), .B2(new_n282), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1214), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n848), .A2(new_n1228), .B1(new_n842), .B2(G128), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n881), .B2(new_n822), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n1227), .B(new_n1230), .C1(G132), .C2(new_n839), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  OR2_X1    g1032(.A1(new_n1232), .A2(KEYINPUT59), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(KEYINPUT59), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n283), .B(new_n253), .C1(new_n833), .C2(new_n1069), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G124), .B2(new_n827), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1233), .A2(new_n1234), .A3(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1065), .B1(new_n880), .B2(new_n406), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n819), .A2(new_n454), .B1(new_n826), .B2(new_n1078), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n833), .A2(new_n202), .B1(new_n822), .B2(new_n430), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n253), .B(new_n346), .C1(new_n817), .C2(new_n392), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n1239), .B(new_n1240), .C1(KEYINPUT117), .C2(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1242), .B1(KEYINPUT117), .B2(new_n1241), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n1238), .B(new_n1243), .C1(G116), .C2(new_n831), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1244), .A2(KEYINPUT58), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(KEYINPUT58), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n201), .B1(new_n344), .B2(G41), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1237), .A2(new_n1245), .A3(new_n1246), .A4(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n812), .ZN(new_n1249));
  XOR2_X1   g1049(.A(new_n1249), .B(KEYINPUT118), .Z(new_n1250));
  AOI211_X1 g1050(.A(new_n798), .B(new_n1250), .C1(new_n201), .C2(new_n888), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n671), .A2(new_n305), .A3(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1252), .B1(new_n302), .B2(new_n306), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n287), .A2(new_n913), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1256), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1251), .B1(new_n1260), .B2(new_n810), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n965), .B1(new_n754), .B2(new_n986), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n964), .B1(new_n1263), .B2(new_n989), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n982), .A2(new_n1264), .A3(new_n1259), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1259), .B1(new_n982), .B2(new_n1264), .ZN(new_n1266));
  OAI21_X1  g1066(.A(KEYINPUT119), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n990), .A2(G330), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n980), .B1(new_n1263), .B2(new_n956), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1260), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n982), .A2(new_n1264), .A3(new_n1259), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT119), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1270), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  AND3_X1   g1073(.A1(new_n954), .A2(KEYINPUT120), .A3(new_n959), .ZN(new_n1274));
  AOI21_X1  g1074(.A(KEYINPUT120), .B1(new_n954), .B2(new_n959), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1267), .B(new_n1273), .C1(new_n1274), .C2(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n960), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1262), .B1(new_n1278), .B2(new_n1058), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1165), .B1(new_n1192), .B2(new_n1197), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(new_n1277), .B2(new_n1276), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1090), .B1(new_n1281), .B2(KEYINPUT57), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT121), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1270), .A2(new_n954), .A3(new_n959), .A4(new_n1271), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(new_n1271), .A2(new_n1270), .B1(new_n954), .B2(new_n959), .ZN(new_n1286));
  OAI21_X1  g1086(.A(KEYINPUT57), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1283), .B1(new_n1287), .B2(new_n1280), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n908), .B1(new_n783), .B2(new_n866), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1181), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(new_n1171), .A2(new_n1179), .B1(new_n1290), .B2(new_n955), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1198), .B1(new_n1203), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1277), .A2(new_n1284), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1292), .A2(KEYINPUT121), .A3(KEYINPUT57), .A4(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1288), .A2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1279), .B1(new_n1282), .B2(new_n1295), .ZN(G375));
  INV_X1    g1096(.A(new_n1036), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1180), .A2(new_n1184), .A3(new_n1165), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1199), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n798), .B1(new_n203), .B2(new_n888), .ZN(new_n1300));
  OAI22_X1  g1100(.A1(new_n882), .A2(new_n875), .B1(new_n837), .B2(new_n201), .ZN(new_n1301));
  AOI22_X1  g1101(.A1(new_n848), .A2(G159), .B1(new_n827), .B2(G128), .ZN(new_n1302));
  OAI221_X1 g1102(.A(new_n1302), .B1(new_n881), .B2(new_n819), .C1(new_n282), .C2(new_n822), .ZN(new_n1303));
  AOI211_X1 g1103(.A(new_n1301), .B(new_n1303), .C1(new_n839), .C2(new_n1228), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n245), .B1(new_n833), .B2(new_n202), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(new_n1305), .B(KEYINPUT122), .ZN(new_n1306));
  AOI22_X1  g1106(.A1(new_n848), .A2(G97), .B1(new_n823), .B2(G107), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1307), .B1(new_n1078), .B2(new_n819), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1308), .B1(G77), .B2(new_n834), .ZN(new_n1309));
  OAI22_X1  g1109(.A1(new_n880), .A2(new_n457), .B1(new_n882), .B2(new_n871), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n346), .B1(new_n826), .B2(new_n531), .ZN(new_n1311));
  NOR3_X1   g1111(.A1(new_n1310), .A2(new_n1104), .A3(new_n1311), .ZN(new_n1312));
  AOI22_X1  g1112(.A1(new_n1304), .A2(new_n1306), .B1(new_n1309), .B2(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1300), .B1(new_n1313), .B2(new_n1207), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1314), .B1(new_n908), .B2(new_n809), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1315), .B1(new_n1197), .B2(new_n1058), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1299), .A2(new_n1316), .ZN(G381));
  NAND2_X1  g1117(.A1(new_n1134), .A2(new_n1089), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(KEYINPUT114), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1134), .A2(new_n1135), .A3(new_n1089), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n1008), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1089), .B1(new_n1323), .B2(new_n1053), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1324), .A2(new_n743), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1160), .B1(new_n1321), .B2(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1326), .A2(new_n1059), .A3(new_n1087), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(G375), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1092), .A2(new_n857), .A3(new_n1126), .ZN(new_n1330));
  NOR4_X1   g1130(.A1(G378), .A2(G384), .A3(G381), .A4(new_n1330), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1328), .A2(new_n1329), .A3(new_n1331), .ZN(G407));
  INV_X1    g1132(.A(G378), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n719), .A2(G213), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1334), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1329), .A2(new_n1333), .A3(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(G407), .A2(G213), .A3(new_n1336), .ZN(G409));
  INV_X1    g1137(.A(KEYINPUT60), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1298), .A2(new_n1338), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1291), .A2(KEYINPUT60), .A3(new_n1165), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1339), .A2(new_n1340), .A3(new_n1199), .A4(new_n1090), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1341), .A2(new_n1316), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(G384), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1341), .A2(new_n894), .A3(new_n1316), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1335), .A2(G2897), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1345), .A2(new_n1346), .ZN(new_n1347));
  NAND4_X1  g1147(.A1(new_n1343), .A2(G2897), .A3(new_n1335), .A4(new_n1344), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT124), .ZN(new_n1349));
  AND3_X1   g1149(.A1(new_n1347), .A2(new_n1348), .A3(new_n1349), .ZN(new_n1350));
  AOI21_X1  g1150(.A(new_n1349), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1351));
  NOR2_X1   g1151(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1352));
  OAI211_X1 g1152(.A(G378), .B(new_n1279), .C1(new_n1282), .C2(new_n1295), .ZN(new_n1353));
  OAI21_X1  g1153(.A(new_n1058), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1354), .A2(new_n1261), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1355), .B1(new_n1281), .B2(new_n1297), .ZN(new_n1356));
  OAI21_X1  g1156(.A(KEYINPUT123), .B1(new_n1356), .B2(G378), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1278), .A2(new_n1297), .A3(new_n1292), .ZN(new_n1358));
  INV_X1    g1158(.A(new_n1355), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1358), .A2(new_n1359), .ZN(new_n1360));
  INV_X1    g1160(.A(KEYINPUT123), .ZN(new_n1361));
  NAND4_X1  g1161(.A1(new_n1360), .A2(new_n1361), .A3(new_n1205), .A4(new_n1225), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1353), .A2(new_n1357), .A3(new_n1362), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1363), .A2(new_n1334), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1352), .A2(new_n1364), .ZN(new_n1365));
  OAI21_X1  g1165(.A(new_n1297), .B1(new_n1324), .B2(new_n793), .ZN(new_n1366));
  INV_X1    g1166(.A(new_n1058), .ZN(new_n1367));
  AOI21_X1  g1167(.A(new_n1034), .B1(new_n1366), .B2(new_n1367), .ZN(new_n1368));
  INV_X1    g1168(.A(new_n1087), .ZN(new_n1369));
  OAI21_X1  g1169(.A(G390), .B1(new_n1368), .B2(new_n1369), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1370), .A2(new_n1327), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(G393), .A2(G396), .ZN(new_n1372));
  AND3_X1   g1172(.A1(new_n1372), .A2(KEYINPUT125), .A3(new_n1330), .ZN(new_n1373));
  AOI21_X1  g1173(.A(KEYINPUT125), .B1(new_n1372), .B2(new_n1330), .ZN(new_n1374));
  OAI21_X1  g1174(.A(new_n1371), .B1(new_n1373), .B2(new_n1374), .ZN(new_n1375));
  INV_X1    g1175(.A(new_n1374), .ZN(new_n1376));
  NAND3_X1  g1176(.A1(new_n1370), .A2(new_n1327), .A3(new_n1376), .ZN(new_n1377));
  AOI21_X1  g1177(.A(KEYINPUT61), .B1(new_n1375), .B2(new_n1377), .ZN(new_n1378));
  NAND3_X1  g1178(.A1(new_n1363), .A2(new_n1334), .A3(new_n1345), .ZN(new_n1379));
  INV_X1    g1179(.A(KEYINPUT63), .ZN(new_n1380));
  OR2_X1    g1180(.A1(new_n1379), .A2(new_n1380), .ZN(new_n1381));
  NAND2_X1  g1181(.A1(new_n1379), .A2(new_n1380), .ZN(new_n1382));
  NAND4_X1  g1182(.A1(new_n1365), .A2(new_n1378), .A3(new_n1381), .A4(new_n1382), .ZN(new_n1383));
  AND2_X1   g1183(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1384));
  NAND2_X1  g1184(.A1(new_n1364), .A2(new_n1384), .ZN(new_n1385));
  INV_X1    g1185(.A(KEYINPUT61), .ZN(new_n1386));
  NAND2_X1  g1186(.A1(new_n1385), .A2(new_n1386), .ZN(new_n1387));
  NOR2_X1   g1187(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1388));
  OR2_X1    g1188(.A1(new_n1379), .A2(new_n1388), .ZN(new_n1389));
  AND2_X1   g1189(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1390));
  AOI21_X1  g1190(.A(new_n1390), .B1(new_n1379), .B2(new_n1388), .ZN(new_n1391));
  AOI21_X1  g1191(.A(new_n1387), .B1(new_n1389), .B2(new_n1391), .ZN(new_n1392));
  NAND2_X1  g1192(.A1(new_n1375), .A2(new_n1377), .ZN(new_n1393));
  OAI21_X1  g1193(.A(new_n1383), .B1(new_n1392), .B2(new_n1393), .ZN(G405));
  NAND2_X1  g1194(.A1(G375), .A2(new_n1333), .ZN(new_n1395));
  NAND2_X1  g1195(.A1(new_n1395), .A2(new_n1353), .ZN(new_n1396));
  NAND2_X1  g1196(.A1(new_n1396), .A2(new_n1345), .ZN(new_n1397));
  NAND4_X1  g1197(.A1(new_n1395), .A2(new_n1353), .A3(new_n1344), .A4(new_n1343), .ZN(new_n1398));
  NAND2_X1  g1198(.A1(new_n1397), .A2(new_n1398), .ZN(new_n1399));
  OAI21_X1  g1199(.A(KEYINPUT127), .B1(new_n1393), .B2(new_n1399), .ZN(new_n1400));
  INV_X1    g1200(.A(new_n1377), .ZN(new_n1401));
  NOR2_X1   g1201(.A1(new_n1373), .A2(new_n1374), .ZN(new_n1402));
  AOI21_X1  g1202(.A(new_n1402), .B1(new_n1370), .B2(new_n1327), .ZN(new_n1403));
  NOR2_X1   g1203(.A1(new_n1401), .A2(new_n1403), .ZN(new_n1404));
  INV_X1    g1204(.A(KEYINPUT127), .ZN(new_n1405));
  NAND4_X1  g1205(.A1(new_n1404), .A2(new_n1405), .A3(new_n1398), .A4(new_n1397), .ZN(new_n1406));
  NAND2_X1  g1206(.A1(new_n1393), .A2(new_n1399), .ZN(new_n1407));
  AND3_X1   g1207(.A1(new_n1400), .A2(new_n1406), .A3(new_n1407), .ZN(G402));
endmodule


