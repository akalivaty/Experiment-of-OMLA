

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747;

  AND2_X1 U367 ( .A1(n583), .A2(n578), .ZN(n590) );
  XNOR2_X1 U368 ( .A(n495), .B(n494), .ZN(n535) );
  NOR2_X1 U369 ( .A1(n688), .A2(n685), .ZN(n624) );
  XOR2_X1 U370 ( .A(KEYINPUT38), .B(n539), .Z(n620) );
  XNOR2_X1 U371 ( .A(n566), .B(KEYINPUT0), .ZN(n594) );
  XNOR2_X1 U372 ( .A(n478), .B(n477), .ZN(n527) );
  INV_X2 U373 ( .A(G953), .ZN(n713) );
  NAND2_X2 U374 ( .A1(n413), .A2(n411), .ZN(n548) );
  AND2_X2 U375 ( .A1(n414), .A2(n417), .ZN(n413) );
  XNOR2_X2 U376 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n362) );
  AND2_X1 U377 ( .A1(n736), .A2(n714), .ZN(n652) );
  AND2_X1 U378 ( .A1(n394), .A2(n348), .ZN(n392) );
  XNOR2_X1 U379 ( .A(n368), .B(KEYINPUT83), .ZN(n542) );
  NOR2_X2 U380 ( .A1(n535), .A2(n536), .ZN(n685) );
  XNOR2_X1 U381 ( .A(n457), .B(n456), .ZN(n519) );
  XNOR2_X1 U382 ( .A(n400), .B(G131), .ZN(n489) );
  XNOR2_X2 U383 ( .A(G143), .B(G128), .ZN(n463) );
  NOR2_X2 U384 ( .A1(n588), .A2(n506), .ZN(n437) );
  XNOR2_X1 U385 ( .A(n380), .B(KEYINPUT84), .ZN(n544) );
  NAND2_X1 U386 ( .A1(n542), .A2(KEYINPUT47), .ZN(n380) );
  XOR2_X1 U387 ( .A(KEYINPUT73), .B(KEYINPUT39), .Z(n479) );
  XNOR2_X1 U388 ( .A(n503), .B(n397), .ZN(n730) );
  XNOR2_X1 U389 ( .A(n489), .B(n398), .ZN(n397) );
  XNOR2_X1 U390 ( .A(n399), .B(G137), .ZN(n398) );
  INV_X1 U391 ( .A(KEYINPUT70), .ZN(n399) );
  XNOR2_X1 U392 ( .A(n722), .B(n451), .ZN(n466) );
  XNOR2_X1 U393 ( .A(n437), .B(KEYINPUT67), .ZN(n555) );
  XNOR2_X1 U394 ( .A(n365), .B(n358), .ZN(n583) );
  NOR2_X1 U395 ( .A1(n594), .A2(n575), .ZN(n365) );
  NOR2_X1 U396 ( .A1(n546), .A2(n545), .ZN(n547) );
  INV_X1 U397 ( .A(KEYINPUT44), .ZN(n586) );
  AND2_X1 U398 ( .A1(n643), .A2(n585), .ZN(n364) );
  XOR2_X1 U399 ( .A(KEYINPUT5), .B(KEYINPUT98), .Z(n452) );
  XNOR2_X1 U400 ( .A(n730), .B(n438), .ZN(n455) );
  NAND2_X1 U401 ( .A1(n349), .A2(n406), .ZN(n370) );
  XNOR2_X1 U402 ( .A(n529), .B(n528), .ZN(n559) );
  XNOR2_X1 U403 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U404 ( .A(KEYINPUT3), .B(KEYINPUT72), .ZN(n449) );
  XOR2_X1 U405 ( .A(KEYINPUT10), .B(KEYINPUT68), .Z(n424) );
  XNOR2_X1 U406 ( .A(n374), .B(n427), .ZN(n373) );
  XOR2_X1 U407 ( .A(G110), .B(G119), .Z(n427) );
  XNOR2_X1 U408 ( .A(n429), .B(n426), .ZN(n374) );
  XNOR2_X1 U409 ( .A(G128), .B(G137), .ZN(n426) );
  XNOR2_X1 U410 ( .A(n428), .B(n376), .ZN(n499) );
  XNOR2_X1 U411 ( .A(n509), .B(n508), .ZN(n512) );
  NAND2_X1 U412 ( .A1(n412), .A2(n415), .ZN(n411) );
  AND2_X1 U413 ( .A1(n620), .A2(n416), .ZN(n415) );
  NAND2_X1 U414 ( .A1(n523), .A2(n382), .ZN(n550) );
  XNOR2_X1 U415 ( .A(n384), .B(n383), .ZN(n382) );
  BUF_X1 U416 ( .A(n527), .Z(n539) );
  XNOR2_X1 U417 ( .A(n525), .B(n396), .ZN(n610) );
  INV_X1 U418 ( .A(KEYINPUT1), .ZN(n396) );
  AND2_X1 U419 ( .A1(n507), .A2(n605), .ZN(n520) );
  XNOR2_X1 U420 ( .A(G902), .B(KEYINPUT15), .ZN(n647) );
  INV_X1 U421 ( .A(KEYINPUT48), .ZN(n377) );
  INV_X1 U422 ( .A(n362), .ZN(n429) );
  INV_X1 U423 ( .A(KEYINPUT69), .ZN(n400) );
  XNOR2_X1 U424 ( .A(G104), .B(G122), .ZN(n485) );
  XNOR2_X1 U425 ( .A(n381), .B(G101), .ZN(n450) );
  INV_X1 U426 ( .A(KEYINPUT4), .ZN(n381) );
  XNOR2_X1 U427 ( .A(n363), .B(n461), .ZN(n465) );
  XOR2_X1 U428 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n461) );
  XNOR2_X1 U429 ( .A(n460), .B(KEYINPUT91), .ZN(n363) );
  AND2_X1 U430 ( .A1(n603), .A2(n423), .ZN(n393) );
  INV_X1 U431 ( .A(n620), .ZN(n418) );
  INV_X1 U432 ( .A(KEYINPUT104), .ZN(n383) );
  XNOR2_X1 U433 ( .A(n455), .B(n385), .ZN(n669) );
  XNOR2_X1 U434 ( .A(n466), .B(n386), .ZN(n385) );
  XNOR2_X1 U435 ( .A(n453), .B(n454), .ZN(n386) );
  XNOR2_X1 U436 ( .A(G110), .B(G104), .ZN(n443) );
  XNOR2_X1 U437 ( .A(KEYINPUT77), .B(KEYINPUT90), .ZN(n442) );
  XNOR2_X1 U438 ( .A(G122), .B(G116), .ZN(n471) );
  XNOR2_X1 U439 ( .A(n463), .B(G134), .ZN(n503) );
  XNOR2_X1 U440 ( .A(n455), .B(n389), .ZN(n699) );
  XNOR2_X1 U441 ( .A(n391), .B(n390), .ZN(n389) );
  XNOR2_X1 U442 ( .A(n450), .B(n356), .ZN(n390) );
  XNOR2_X1 U443 ( .A(n441), .B(n468), .ZN(n391) );
  AND2_X2 U444 ( .A1(n420), .A2(n419), .ZN(n698) );
  NAND2_X1 U445 ( .A1(n652), .A2(KEYINPUT2), .ZN(n419) );
  XNOR2_X1 U446 ( .A(n421), .B(KEYINPUT64), .ZN(n420) );
  NAND2_X1 U447 ( .A1(n422), .A2(n361), .ZN(n421) );
  NOR2_X1 U448 ( .A1(n530), .A2(n559), .ZN(n368) );
  NAND2_X1 U449 ( .A1(n555), .A2(n410), .ZN(n409) );
  NAND2_X1 U450 ( .A1(n371), .A2(n407), .ZN(n406) );
  XNOR2_X1 U451 ( .A(n669), .B(KEYINPUT62), .ZN(n670) );
  INV_X1 U452 ( .A(G101), .ZN(n723) );
  XNOR2_X1 U453 ( .A(n372), .B(n401), .ZN(n403) );
  XNOR2_X1 U454 ( .A(n373), .B(n375), .ZN(n372) );
  NAND2_X1 U455 ( .A1(n499), .A2(G221), .ZN(n375) );
  XNOR2_X1 U456 ( .A(n663), .B(n662), .ZN(n664) );
  BUF_X1 U457 ( .A(n698), .Z(n708) );
  NOR2_X1 U458 ( .A1(n550), .A2(n395), .ZN(n551) );
  XNOR2_X1 U459 ( .A(KEYINPUT107), .B(KEYINPUT40), .ZN(n504) );
  AND2_X1 U460 ( .A1(n526), .A2(n395), .ZN(n691) );
  XNOR2_X1 U461 ( .A(n580), .B(KEYINPUT32), .ZN(n643) );
  NOR2_X1 U462 ( .A1(n610), .A2(n604), .ZN(n579) );
  NOR2_X1 U463 ( .A1(n581), .A2(n395), .ZN(n582) );
  AND2_X1 U464 ( .A1(n610), .A2(n604), .ZN(n589) );
  XOR2_X1 U465 ( .A(G113), .B(G119), .Z(n347) );
  AND2_X1 U466 ( .A1(n554), .A2(n360), .ZN(n348) );
  INV_X1 U467 ( .A(n610), .ZN(n395) );
  AND2_X1 U468 ( .A1(n409), .A2(n405), .ZN(n349) );
  OR2_X1 U469 ( .A1(n705), .A2(G902), .ZN(n350) );
  BUF_X1 U470 ( .A(n588), .Z(n369) );
  OR2_X1 U471 ( .A1(n564), .A2(n563), .ZN(n351) );
  XOR2_X1 U472 ( .A(KEYINPUT71), .B(n547), .Z(n352) );
  XOR2_X1 U473 ( .A(KEYINPUT30), .B(n459), .Z(n353) );
  XOR2_X1 U474 ( .A(KEYINPUT118), .B(n640), .Z(n354) );
  OR2_X1 U475 ( .A1(n563), .A2(n448), .ZN(n355) );
  AND2_X1 U476 ( .A1(G227), .A2(n713), .ZN(n356) );
  AND2_X1 U477 ( .A1(n409), .A2(n408), .ZN(n357) );
  XOR2_X1 U478 ( .A(n576), .B(KEYINPUT22), .Z(n358) );
  XOR2_X1 U479 ( .A(KEYINPUT86), .B(KEYINPUT45), .Z(n359) );
  NAND2_X1 U480 ( .A1(n648), .A2(n647), .ZN(n360) );
  NAND2_X1 U481 ( .A1(n360), .A2(n651), .ZN(n361) );
  INV_X1 U482 ( .A(G146), .ZN(n438) );
  NAND2_X1 U483 ( .A1(n548), .A2(n685), .ZN(n505) );
  NAND2_X1 U484 ( .A1(n364), .A2(n742), .ZN(n587) );
  NAND2_X1 U485 ( .A1(n366), .A2(n352), .ZN(n378) );
  XNOR2_X1 U486 ( .A(n379), .B(KEYINPUT46), .ZN(n366) );
  NOR2_X2 U487 ( .A1(n659), .A2(n712), .ZN(n661) );
  NOR2_X2 U488 ( .A1(n666), .A2(n712), .ZN(n668) );
  NAND2_X1 U489 ( .A1(n520), .A2(n519), .ZN(n509) );
  XNOR2_X1 U490 ( .A(n367), .B(n673), .ZN(G57) );
  NOR2_X2 U491 ( .A1(n672), .A2(n712), .ZN(n367) );
  XNOR2_X1 U492 ( .A(n370), .B(KEYINPUT79), .ZN(n388) );
  INV_X1 U493 ( .A(n555), .ZN(n371) );
  INV_X1 U494 ( .A(KEYINPUT8), .ZN(n376) );
  XNOR2_X2 U495 ( .A(n378), .B(n377), .ZN(n394) );
  NOR2_X2 U496 ( .A1(n743), .A2(n746), .ZN(n379) );
  INV_X1 U497 ( .A(n542), .ZN(n683) );
  NAND2_X1 U498 ( .A1(n577), .A2(n520), .ZN(n384) );
  XNOR2_X1 U499 ( .A(n519), .B(n518), .ZN(n577) );
  XNOR2_X2 U500 ( .A(n387), .B(KEYINPUT78), .ZN(n534) );
  NAND2_X1 U501 ( .A1(n388), .A2(n353), .ZN(n387) );
  XNOR2_X1 U502 ( .A(n524), .B(KEYINPUT36), .ZN(n526) );
  NOR2_X2 U503 ( .A1(n699), .A2(G902), .ZN(n511) );
  AND2_X1 U504 ( .A1(n394), .A2(n554), .ZN(n736) );
  NAND2_X1 U505 ( .A1(n392), .A2(n714), .ZN(n422) );
  XNOR2_X2 U506 ( .A(n393), .B(n359), .ZN(n714) );
  NAND2_X1 U507 ( .A1(n403), .A2(n402), .ZN(n404) );
  INV_X1 U508 ( .A(n480), .ZN(n401) );
  INV_X1 U509 ( .A(n403), .ZN(n710) );
  INV_X1 U510 ( .A(G902), .ZN(n402) );
  XNOR2_X2 U511 ( .A(n404), .B(n433), .ZN(n588) );
  AND2_X1 U512 ( .A1(n408), .A2(n355), .ZN(n405) );
  NAND2_X1 U513 ( .A1(n444), .A2(n410), .ZN(n408) );
  NAND2_X1 U514 ( .A1(n357), .A2(n406), .ZN(n596) );
  NOR2_X1 U515 ( .A1(n444), .A2(n410), .ZN(n407) );
  INV_X1 U516 ( .A(KEYINPUT97), .ZN(n410) );
  INV_X1 U517 ( .A(n534), .ZN(n412) );
  NAND2_X1 U518 ( .A1(n534), .A2(n479), .ZN(n414) );
  INV_X1 U519 ( .A(n479), .ZN(n416) );
  NAND2_X1 U520 ( .A1(n418), .A2(n479), .ZN(n417) );
  XNOR2_X1 U521 ( .A(n425), .B(n424), .ZN(n480) );
  XNOR2_X1 U522 ( .A(n462), .B(G140), .ZN(n425) );
  AND2_X1 U523 ( .A1(n355), .A2(n588), .ZN(n507) );
  AND2_X1 U524 ( .A1(n602), .A2(n601), .ZN(n423) );
  INV_X1 U525 ( .A(n619), .ZN(n521) );
  XNOR2_X1 U526 ( .A(n452), .B(G116), .ZN(n453) );
  XNOR2_X1 U527 ( .A(n587), .B(n586), .ZN(n603) );
  AND2_X1 U528 ( .A1(n658), .A2(G953), .ZN(n712) );
  BUF_X1 U529 ( .A(n743), .Z(n744) );
  XNOR2_X1 U530 ( .A(n642), .B(n641), .ZN(G75) );
  XOR2_X2 U531 ( .A(G146), .B(G125), .Z(n462) );
  NAND2_X1 U532 ( .A1(G234), .A2(n713), .ZN(n428) );
  NAND2_X1 U533 ( .A1(G234), .A2(n647), .ZN(n430) );
  XNOR2_X1 U534 ( .A(KEYINPUT20), .B(n430), .ZN(n434) );
  AND2_X1 U535 ( .A1(n434), .A2(G217), .ZN(n432) );
  XNOR2_X1 U536 ( .A(KEYINPUT95), .B(KEYINPUT25), .ZN(n431) );
  NAND2_X1 U537 ( .A1(G221), .A2(n434), .ZN(n436) );
  XNOR2_X1 U538 ( .A(KEYINPUT96), .B(KEYINPUT21), .ZN(n435) );
  XNOR2_X1 U539 ( .A(n436), .B(n435), .ZN(n506) );
  XOR2_X1 U540 ( .A(KEYINPUT80), .B(KEYINPUT81), .Z(n440) );
  XNOR2_X1 U541 ( .A(G107), .B(G140), .ZN(n439) );
  XNOR2_X1 U542 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U543 ( .A(n443), .B(n442), .ZN(n468) );
  INV_X1 U544 ( .A(G469), .ZN(n510) );
  XNOR2_X1 U545 ( .A(n511), .B(G469), .ZN(n444) );
  NAND2_X1 U546 ( .A1(G234), .A2(G237), .ZN(n445) );
  XNOR2_X1 U547 ( .A(n445), .B(KEYINPUT14), .ZN(n446) );
  NAND2_X1 U548 ( .A1(G952), .A2(n446), .ZN(n633) );
  NOR2_X1 U549 ( .A1(n633), .A2(G953), .ZN(n563) );
  NAND2_X1 U550 ( .A1(G902), .A2(n446), .ZN(n561) );
  OR2_X1 U551 ( .A1(n713), .A2(n561), .ZN(n447) );
  NOR2_X1 U552 ( .A1(G900), .A2(n447), .ZN(n448) );
  NOR2_X1 U553 ( .A1(G953), .A2(G237), .ZN(n482) );
  NAND2_X1 U554 ( .A1(G210), .A2(n482), .ZN(n454) );
  XNOR2_X1 U555 ( .A(n347), .B(n449), .ZN(n722) );
  INV_X1 U556 ( .A(n450), .ZN(n451) );
  NOR2_X1 U557 ( .A1(G902), .A2(n669), .ZN(n457) );
  INV_X1 U558 ( .A(G472), .ZN(n456) );
  BUF_X2 U559 ( .A(n519), .Z(n608) );
  INV_X1 U560 ( .A(G237), .ZN(n458) );
  NAND2_X1 U561 ( .A1(n402), .A2(n458), .ZN(n474) );
  NAND2_X1 U562 ( .A1(n474), .A2(G214), .ZN(n619) );
  NAND2_X1 U563 ( .A1(n608), .A2(n619), .ZN(n459) );
  NAND2_X1 U564 ( .A1(G224), .A2(n713), .ZN(n460) );
  XNOR2_X1 U565 ( .A(n462), .B(n463), .ZN(n464) );
  XNOR2_X1 U566 ( .A(n465), .B(n464), .ZN(n467) );
  XNOR2_X1 U567 ( .A(n467), .B(n466), .ZN(n473) );
  INV_X1 U568 ( .A(n468), .ZN(n470) );
  XNOR2_X1 U569 ( .A(KEYINPUT75), .B(KEYINPUT16), .ZN(n469) );
  XNOR2_X1 U570 ( .A(n470), .B(n469), .ZN(n472) );
  XNOR2_X1 U571 ( .A(n471), .B(G107), .ZN(n498) );
  XNOR2_X1 U572 ( .A(n472), .B(n498), .ZN(n725) );
  XNOR2_X1 U573 ( .A(n473), .B(n725), .ZN(n655) );
  NAND2_X1 U574 ( .A1(n655), .A2(n647), .ZN(n478) );
  NAND2_X1 U575 ( .A1(n474), .A2(G210), .ZN(n476) );
  INV_X1 U576 ( .A(KEYINPUT92), .ZN(n475) );
  XNOR2_X1 U577 ( .A(n476), .B(n475), .ZN(n477) );
  BUF_X1 U578 ( .A(n480), .Z(n481) );
  XOR2_X1 U579 ( .A(n481), .B(G113), .Z(n493) );
  XOR2_X1 U580 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n484) );
  NAND2_X1 U581 ( .A1(G214), .A2(n482), .ZN(n483) );
  XNOR2_X1 U582 ( .A(n484), .B(n483), .ZN(n488) );
  XOR2_X1 U583 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n486) );
  XNOR2_X1 U584 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U585 ( .A(n488), .B(n487), .ZN(n491) );
  XNOR2_X1 U586 ( .A(G143), .B(n489), .ZN(n490) );
  XNOR2_X1 U587 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U588 ( .A(n493), .B(n492), .ZN(n663) );
  NAND2_X1 U589 ( .A1(n663), .A2(n402), .ZN(n495) );
  XNOR2_X1 U590 ( .A(KEYINPUT13), .B(G475), .ZN(n494) );
  XNOR2_X1 U591 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n496) );
  XNOR2_X1 U592 ( .A(n496), .B(KEYINPUT101), .ZN(n497) );
  XOR2_X1 U593 ( .A(n498), .B(n497), .Z(n501) );
  NAND2_X1 U594 ( .A1(G217), .A2(n499), .ZN(n500) );
  XNOR2_X1 U595 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U596 ( .A(n503), .B(n502), .ZN(n705) );
  XNOR2_X1 U597 ( .A(G478), .B(n350), .ZN(n536) );
  XNOR2_X2 U598 ( .A(n505), .B(n504), .ZN(n743) );
  INV_X1 U599 ( .A(n506), .ZN(n605) );
  XNOR2_X1 U600 ( .A(KEYINPUT105), .B(KEYINPUT28), .ZN(n508) );
  XNOR2_X1 U601 ( .A(n511), .B(n510), .ZN(n525) );
  NAND2_X1 U602 ( .A1(n512), .A2(n525), .ZN(n513) );
  XNOR2_X1 U603 ( .A(n513), .B(KEYINPUT106), .ZN(n530) );
  INV_X1 U604 ( .A(n536), .ZN(n514) );
  AND2_X1 U605 ( .A1(n535), .A2(n514), .ZN(n574) );
  INV_X1 U606 ( .A(n574), .ZN(n622) );
  NAND2_X1 U607 ( .A1(n620), .A2(n619), .ZN(n623) );
  NOR2_X1 U608 ( .A1(n622), .A2(n623), .ZN(n516) );
  XNOR2_X1 U609 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n515) );
  XNOR2_X1 U610 ( .A(n516), .B(n515), .ZN(n635) );
  NOR2_X1 U611 ( .A1(n530), .A2(n635), .ZN(n517) );
  XNOR2_X1 U612 ( .A(n517), .B(KEYINPUT42), .ZN(n746) );
  INV_X1 U613 ( .A(KEYINPUT6), .ZN(n518) );
  INV_X1 U614 ( .A(n685), .ZN(n522) );
  NOR2_X1 U615 ( .A1(n522), .A2(n521), .ZN(n523) );
  INV_X1 U616 ( .A(n539), .ZN(n552) );
  NOR2_X1 U617 ( .A1(n550), .A2(n552), .ZN(n524) );
  NAND2_X1 U618 ( .A1(n527), .A2(n619), .ZN(n529) );
  XNOR2_X1 U619 ( .A(KEYINPUT65), .B(KEYINPUT19), .ZN(n528) );
  AND2_X1 U620 ( .A1(n535), .A2(n536), .ZN(n688) );
  NOR2_X1 U621 ( .A1(KEYINPUT47), .A2(n624), .ZN(n531) );
  XOR2_X1 U622 ( .A(KEYINPUT76), .B(n531), .Z(n532) );
  NOR2_X1 U623 ( .A1(n542), .A2(n532), .ZN(n533) );
  NOR2_X1 U624 ( .A1(n691), .A2(n533), .ZN(n541) );
  BUF_X1 U625 ( .A(n534), .Z(n538) );
  INV_X1 U626 ( .A(n535), .ZN(n537) );
  NAND2_X1 U627 ( .A1(n537), .A2(n536), .ZN(n568) );
  NOR2_X1 U628 ( .A1(n538), .A2(n568), .ZN(n540) );
  NAND2_X1 U629 ( .A1(n540), .A2(n539), .ZN(n644) );
  NAND2_X1 U630 ( .A1(n541), .A2(n644), .ZN(n546) );
  NAND2_X1 U631 ( .A1(n624), .A2(KEYINPUT47), .ZN(n543) );
  NAND2_X1 U632 ( .A1(n544), .A2(n543), .ZN(n545) );
  BUF_X1 U633 ( .A(n548), .Z(n549) );
  NAND2_X1 U634 ( .A1(n549), .A2(n688), .ZN(n695) );
  XOR2_X1 U635 ( .A(n551), .B(KEYINPUT43), .Z(n553) );
  NAND2_X1 U636 ( .A1(n553), .A2(n552), .ZN(n696) );
  AND2_X1 U637 ( .A1(n695), .A2(n696), .ZN(n554) );
  XOR2_X1 U638 ( .A(KEYINPUT88), .B(KEYINPUT33), .Z(n558) );
  BUF_X1 U639 ( .A(n555), .Z(n556) );
  NOR2_X1 U640 ( .A1(n610), .A2(n556), .ZN(n593) );
  NAND2_X1 U641 ( .A1(n593), .A2(n577), .ZN(n557) );
  XNOR2_X1 U642 ( .A(n558), .B(n557), .ZN(n634) );
  INV_X1 U643 ( .A(n559), .ZN(n565) );
  NOR2_X1 U644 ( .A1(G898), .A2(n713), .ZN(n560) );
  XNOR2_X1 U645 ( .A(KEYINPUT93), .B(n560), .ZN(n726) );
  NOR2_X1 U646 ( .A1(n561), .A2(n726), .ZN(n562) );
  XNOR2_X1 U647 ( .A(n562), .B(KEYINPUT94), .ZN(n564) );
  NAND2_X1 U648 ( .A1(n565), .A2(n351), .ZN(n566) );
  NOR2_X1 U649 ( .A1(n634), .A2(n594), .ZN(n567) );
  XNOR2_X1 U650 ( .A(n567), .B(KEYINPUT34), .ZN(n570) );
  INV_X1 U651 ( .A(n568), .ZN(n569) );
  NAND2_X1 U652 ( .A1(n570), .A2(n569), .ZN(n573) );
  INV_X1 U653 ( .A(KEYINPUT82), .ZN(n571) );
  XNOR2_X1 U654 ( .A(n571), .B(KEYINPUT35), .ZN(n572) );
  XNOR2_X1 U655 ( .A(n573), .B(n572), .ZN(n742) );
  NAND2_X1 U656 ( .A1(n574), .A2(n605), .ZN(n575) );
  INV_X1 U657 ( .A(KEYINPUT74), .ZN(n576) );
  INV_X1 U658 ( .A(n577), .ZN(n578) );
  NAND2_X1 U659 ( .A1(n590), .A2(n579), .ZN(n580) );
  INV_X1 U660 ( .A(n369), .ZN(n604) );
  OR2_X1 U661 ( .A1(n608), .A2(n604), .ZN(n581) );
  NAND2_X1 U662 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U663 ( .A(n584), .B(KEYINPUT103), .ZN(n741) );
  INV_X1 U664 ( .A(n741), .ZN(n585) );
  NAND2_X1 U665 ( .A1(n590), .A2(n589), .ZN(n592) );
  INV_X1 U666 ( .A(KEYINPUT102), .ZN(n591) );
  XNOR2_X1 U667 ( .A(n592), .B(n591), .ZN(n747) );
  INV_X1 U668 ( .A(n747), .ZN(n602) );
  AND2_X1 U669 ( .A1(n593), .A2(n608), .ZN(n615) );
  INV_X1 U670 ( .A(n594), .ZN(n597) );
  NAND2_X1 U671 ( .A1(n615), .A2(n597), .ZN(n595) );
  XNOR2_X1 U672 ( .A(n595), .B(KEYINPUT31), .ZN(n689) );
  NOR2_X1 U673 ( .A1(n596), .A2(n608), .ZN(n598) );
  AND2_X1 U674 ( .A1(n598), .A2(n597), .ZN(n676) );
  OR2_X1 U675 ( .A1(n689), .A2(n676), .ZN(n600) );
  INV_X1 U676 ( .A(n624), .ZN(n599) );
  NAND2_X1 U677 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U678 ( .A(n652), .B(KEYINPUT2), .ZN(n639) );
  XNOR2_X1 U679 ( .A(KEYINPUT51), .B(KEYINPUT116), .ZN(n617) );
  NOR2_X1 U680 ( .A1(n605), .A2(n604), .ZN(n606) );
  XOR2_X1 U681 ( .A(KEYINPUT49), .B(n606), .Z(n607) );
  NOR2_X1 U682 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U683 ( .A(KEYINPUT115), .B(n609), .ZN(n613) );
  NAND2_X1 U684 ( .A1(n610), .A2(n556), .ZN(n611) );
  XOR2_X1 U685 ( .A(KEYINPUT50), .B(n611), .Z(n612) );
  NOR2_X1 U686 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U687 ( .A1(n615), .A2(n614), .ZN(n616) );
  XOR2_X1 U688 ( .A(n617), .B(n616), .Z(n618) );
  NOR2_X1 U689 ( .A1(n635), .A2(n618), .ZN(n629) );
  NOR2_X1 U690 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U691 ( .A1(n622), .A2(n621), .ZN(n626) );
  NOR2_X1 U692 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U693 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U694 ( .A1(n634), .A2(n627), .ZN(n628) );
  NOR2_X1 U695 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U696 ( .A(n630), .B(KEYINPUT117), .Z(n631) );
  XNOR2_X1 U697 ( .A(KEYINPUT52), .B(n631), .ZN(n632) );
  NOR2_X1 U698 ( .A1(n633), .A2(n632), .ZN(n637) );
  NOR2_X1 U699 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U700 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U701 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U702 ( .A1(n713), .A2(n354), .ZN(n642) );
  XNOR2_X1 U703 ( .A(KEYINPUT119), .B(KEYINPUT53), .ZN(n641) );
  XNOR2_X1 U704 ( .A(n643), .B(G119), .ZN(G21) );
  XNOR2_X1 U705 ( .A(n644), .B(G143), .ZN(G45) );
  INV_X1 U706 ( .A(n647), .ZN(n646) );
  NAND2_X1 U707 ( .A1(KEYINPUT2), .A2(KEYINPUT85), .ZN(n645) );
  NOR2_X1 U708 ( .A1(n646), .A2(n645), .ZN(n649) );
  INV_X1 U709 ( .A(n649), .ZN(n648) );
  INV_X1 U710 ( .A(KEYINPUT2), .ZN(n653) );
  NOR2_X1 U711 ( .A1(n653), .A2(KEYINPUT85), .ZN(n650) );
  OR2_X1 U712 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U713 ( .A1(n698), .A2(G210), .ZN(n657) );
  XNOR2_X1 U714 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n654) );
  XNOR2_X1 U715 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U716 ( .A(n657), .B(n656), .ZN(n659) );
  INV_X1 U717 ( .A(G952), .ZN(n658) );
  XNOR2_X1 U718 ( .A(KEYINPUT120), .B(KEYINPUT56), .ZN(n660) );
  XNOR2_X1 U719 ( .A(n661), .B(n660), .ZN(G51) );
  NAND2_X1 U720 ( .A1(n698), .A2(G475), .ZN(n665) );
  XOR2_X1 U721 ( .A(KEYINPUT89), .B(KEYINPUT59), .Z(n662) );
  XNOR2_X1 U722 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U723 ( .A(KEYINPUT66), .B(KEYINPUT60), .ZN(n667) );
  XNOR2_X1 U724 ( .A(n668), .B(n667), .ZN(G60) );
  NAND2_X1 U725 ( .A1(n698), .A2(G472), .ZN(n671) );
  XNOR2_X1 U726 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U727 ( .A(KEYINPUT63), .B(KEYINPUT87), .ZN(n673) );
  XOR2_X1 U728 ( .A(G104), .B(KEYINPUT109), .Z(n675) );
  NAND2_X1 U729 ( .A1(n676), .A2(n685), .ZN(n674) );
  XNOR2_X1 U730 ( .A(n675), .B(n674), .ZN(G6) );
  XNOR2_X1 U731 ( .A(G107), .B(KEYINPUT110), .ZN(n680) );
  XOR2_X1 U732 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n678) );
  NAND2_X1 U733 ( .A1(n676), .A2(n688), .ZN(n677) );
  XNOR2_X1 U734 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U735 ( .A(n680), .B(n679), .ZN(G9) );
  XOR2_X1 U736 ( .A(G128), .B(KEYINPUT29), .Z(n682) );
  NAND2_X1 U737 ( .A1(n683), .A2(n688), .ZN(n681) );
  XNOR2_X1 U738 ( .A(n682), .B(n681), .ZN(G30) );
  NAND2_X1 U739 ( .A1(n683), .A2(n685), .ZN(n684) );
  XNOR2_X1 U740 ( .A(n684), .B(G146), .ZN(G48) );
  XOR2_X1 U741 ( .A(G113), .B(KEYINPUT111), .Z(n687) );
  NAND2_X1 U742 ( .A1(n689), .A2(n685), .ZN(n686) );
  XNOR2_X1 U743 ( .A(n687), .B(n686), .ZN(G15) );
  NAND2_X1 U744 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U745 ( .A(n690), .B(G116), .ZN(G18) );
  XNOR2_X1 U746 ( .A(n691), .B(KEYINPUT37), .ZN(n692) );
  XNOR2_X1 U747 ( .A(n692), .B(KEYINPUT112), .ZN(n693) );
  XNOR2_X1 U748 ( .A(G125), .B(n693), .ZN(G27) );
  XOR2_X1 U749 ( .A(G134), .B(KEYINPUT113), .Z(n694) );
  XNOR2_X1 U750 ( .A(n695), .B(n694), .ZN(G36) );
  XNOR2_X1 U751 ( .A(n696), .B(G140), .ZN(n697) );
  XNOR2_X1 U752 ( .A(KEYINPUT114), .B(n697), .ZN(G42) );
  NAND2_X1 U753 ( .A1(n708), .A2(G469), .ZN(n703) );
  XNOR2_X1 U754 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n701) );
  XNOR2_X1 U755 ( .A(n699), .B(KEYINPUT57), .ZN(n700) );
  XNOR2_X1 U756 ( .A(n701), .B(n700), .ZN(n702) );
  XNOR2_X1 U757 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U758 ( .A1(n712), .A2(n704), .ZN(G54) );
  NAND2_X1 U759 ( .A1(n708), .A2(G478), .ZN(n706) );
  XNOR2_X1 U760 ( .A(n706), .B(n705), .ZN(n707) );
  NOR2_X1 U761 ( .A1(n712), .A2(n707), .ZN(G63) );
  NAND2_X1 U762 ( .A1(n708), .A2(G217), .ZN(n709) );
  XNOR2_X1 U763 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X1 U764 ( .A1(n712), .A2(n711), .ZN(G66) );
  NAND2_X1 U765 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U766 ( .A(n715), .B(KEYINPUT123), .ZN(n720) );
  NAND2_X1 U767 ( .A1(G953), .A2(G224), .ZN(n716) );
  XNOR2_X1 U768 ( .A(KEYINPUT61), .B(n716), .ZN(n717) );
  NAND2_X1 U769 ( .A1(n717), .A2(G898), .ZN(n718) );
  XOR2_X1 U770 ( .A(n718), .B(KEYINPUT122), .Z(n719) );
  NOR2_X1 U771 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U772 ( .A(KEYINPUT124), .B(n721), .Z(n729) );
  XNOR2_X1 U773 ( .A(n722), .B(n723), .ZN(n724) );
  XNOR2_X1 U774 ( .A(n725), .B(n724), .ZN(n727) );
  NAND2_X1 U775 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U776 ( .A(n729), .B(n728), .Z(G69) );
  XNOR2_X1 U777 ( .A(n730), .B(KEYINPUT4), .ZN(n731) );
  XNOR2_X1 U778 ( .A(n481), .B(n731), .ZN(n735) );
  XNOR2_X1 U779 ( .A(G227), .B(n735), .ZN(n732) );
  NAND2_X1 U780 ( .A1(n732), .A2(G900), .ZN(n733) );
  NAND2_X1 U781 ( .A1(n733), .A2(G953), .ZN(n734) );
  XNOR2_X1 U782 ( .A(n734), .B(KEYINPUT125), .ZN(n739) );
  XNOR2_X1 U783 ( .A(n736), .B(n735), .ZN(n737) );
  NOR2_X1 U784 ( .A1(n737), .A2(G953), .ZN(n738) );
  NOR2_X1 U785 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U786 ( .A(KEYINPUT126), .B(n740), .Z(G72) );
  XOR2_X1 U787 ( .A(G110), .B(n741), .Z(G12) );
  XNOR2_X1 U788 ( .A(G122), .B(n742), .ZN(G24) );
  XNOR2_X1 U789 ( .A(G131), .B(KEYINPUT127), .ZN(n745) );
  XNOR2_X1 U790 ( .A(n745), .B(n744), .ZN(G33) );
  XOR2_X1 U791 ( .A(G137), .B(n746), .Z(G39) );
  XOR2_X1 U792 ( .A(G101), .B(n747), .Z(G3) );
endmodule

