

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U548 ( .A(KEYINPUT30), .B(KEYINPUT98), .ZN(n647) );
  XNOR2_X1 U549 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U550 ( .A(KEYINPUT101), .B(KEYINPUT31), .ZN(n656) );
  XNOR2_X1 U551 ( .A(n657), .B(n656), .ZN(n658) );
  AND2_X1 U552 ( .A1(n666), .A2(n661), .ZN(n664) );
  XNOR2_X1 U553 ( .A(n580), .B(KEYINPUT23), .ZN(n581) );
  NOR2_X1 U554 ( .A1(n530), .A2(G2105), .ZN(n579) );
  NOR2_X1 U555 ( .A1(n588), .A2(n587), .ZN(n590) );
  XNOR2_X1 U556 ( .A(n592), .B(n591), .ZN(n758) );
  XOR2_X1 U557 ( .A(G543), .B(KEYINPUT0), .Z(n565) );
  NOR2_X1 U558 ( .A1(G651), .A2(n565), .ZN(n787) );
  NAND2_X1 U559 ( .A1(G52), .A2(n787), .ZN(n521) );
  INV_X1 U560 ( .A(G651), .ZN(n523) );
  NOR2_X1 U561 ( .A1(G543), .A2(n523), .ZN(n518) );
  XOR2_X1 U562 ( .A(KEYINPUT68), .B(n518), .Z(n519) );
  XNOR2_X1 U563 ( .A(KEYINPUT1), .B(n519), .ZN(n788) );
  NAND2_X1 U564 ( .A1(G64), .A2(n788), .ZN(n520) );
  NAND2_X1 U565 ( .A1(n521), .A2(n520), .ZN(n528) );
  NOR2_X1 U566 ( .A1(G651), .A2(G543), .ZN(n783) );
  NAND2_X1 U567 ( .A1(n783), .A2(G90), .ZN(n522) );
  XNOR2_X1 U568 ( .A(n522), .B(KEYINPUT70), .ZN(n525) );
  NOR2_X1 U569 ( .A1(n565), .A2(n523), .ZN(n784) );
  NAND2_X1 U570 ( .A1(G77), .A2(n784), .ZN(n524) );
  NAND2_X1 U571 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U572 ( .A(KEYINPUT9), .B(n526), .Z(n527) );
  NOR2_X1 U573 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U574 ( .A(KEYINPUT71), .B(n529), .Z(G171) );
  INV_X1 U575 ( .A(G171), .ZN(G301) );
  INV_X1 U576 ( .A(G2104), .ZN(n530) );
  BUF_X1 U577 ( .A(n579), .Z(n994) );
  NAND2_X1 U578 ( .A1(G102), .A2(n994), .ZN(n533) );
  NOR2_X1 U579 ( .A1(G2104), .A2(G2105), .ZN(n531) );
  XOR2_X1 U580 ( .A(KEYINPUT17), .B(n531), .Z(n585) );
  BUF_X1 U581 ( .A(n585), .Z(n995) );
  NAND2_X1 U582 ( .A1(G138), .A2(n995), .ZN(n532) );
  NAND2_X1 U583 ( .A1(n533), .A2(n532), .ZN(n538) );
  AND2_X1 U584 ( .A1(G2104), .A2(G2105), .ZN(n990) );
  NAND2_X1 U585 ( .A1(G114), .A2(n990), .ZN(n535) );
  AND2_X1 U586 ( .A1(n530), .A2(G2105), .ZN(n991) );
  NAND2_X1 U587 ( .A1(G126), .A2(n991), .ZN(n534) );
  NAND2_X1 U588 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U589 ( .A(KEYINPUT87), .B(n536), .Z(n537) );
  NOR2_X1 U590 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U591 ( .A(KEYINPUT88), .B(n539), .ZN(G164) );
  NAND2_X1 U592 ( .A1(n783), .A2(G89), .ZN(n540) );
  XNOR2_X1 U593 ( .A(n540), .B(KEYINPUT4), .ZN(n542) );
  NAND2_X1 U594 ( .A1(G76), .A2(n784), .ZN(n541) );
  NAND2_X1 U595 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U596 ( .A(n543), .B(KEYINPUT5), .ZN(n548) );
  NAND2_X1 U597 ( .A1(G51), .A2(n787), .ZN(n545) );
  NAND2_X1 U598 ( .A1(G63), .A2(n788), .ZN(n544) );
  NAND2_X1 U599 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U600 ( .A(KEYINPUT6), .B(n546), .Z(n547) );
  NAND2_X1 U601 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U602 ( .A(n549), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U603 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U604 ( .A1(G88), .A2(n783), .ZN(n551) );
  NAND2_X1 U605 ( .A1(G75), .A2(n784), .ZN(n550) );
  NAND2_X1 U606 ( .A1(n551), .A2(n550), .ZN(n556) );
  NAND2_X1 U607 ( .A1(n787), .A2(G50), .ZN(n552) );
  XNOR2_X1 U608 ( .A(n552), .B(KEYINPUT84), .ZN(n554) );
  NAND2_X1 U609 ( .A1(G62), .A2(n788), .ZN(n553) );
  NAND2_X1 U610 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U611 ( .A1(n556), .A2(n555), .ZN(G166) );
  XNOR2_X1 U612 ( .A(G166), .B(KEYINPUT89), .ZN(G303) );
  NAND2_X1 U613 ( .A1(G86), .A2(n783), .ZN(n558) );
  NAND2_X1 U614 ( .A1(G48), .A2(n787), .ZN(n557) );
  NAND2_X1 U615 ( .A1(n558), .A2(n557), .ZN(n561) );
  NAND2_X1 U616 ( .A1(n784), .A2(G73), .ZN(n559) );
  XOR2_X1 U617 ( .A(KEYINPUT2), .B(n559), .Z(n560) );
  NOR2_X1 U618 ( .A1(n561), .A2(n560), .ZN(n563) );
  NAND2_X1 U619 ( .A1(G61), .A2(n788), .ZN(n562) );
  NAND2_X1 U620 ( .A1(n563), .A2(n562), .ZN(G305) );
  NAND2_X1 U621 ( .A1(G49), .A2(n787), .ZN(n564) );
  XNOR2_X1 U622 ( .A(n564), .B(KEYINPUT82), .ZN(n570) );
  NAND2_X1 U623 ( .A1(G87), .A2(n565), .ZN(n567) );
  NAND2_X1 U624 ( .A1(G74), .A2(G651), .ZN(n566) );
  NAND2_X1 U625 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U626 ( .A1(n788), .A2(n568), .ZN(n569) );
  NAND2_X1 U627 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U628 ( .A(KEYINPUT83), .B(n571), .Z(G288) );
  NAND2_X1 U629 ( .A1(G85), .A2(n783), .ZN(n573) );
  NAND2_X1 U630 ( .A1(G72), .A2(n784), .ZN(n572) );
  NAND2_X1 U631 ( .A1(n573), .A2(n572), .ZN(n577) );
  NAND2_X1 U632 ( .A1(G47), .A2(n787), .ZN(n575) );
  NAND2_X1 U633 ( .A1(G60), .A2(n788), .ZN(n574) );
  NAND2_X1 U634 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U635 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U636 ( .A(KEYINPUT69), .B(n578), .ZN(G290) );
  INV_X1 U637 ( .A(KEYINPUT64), .ZN(n592) );
  NAND2_X1 U638 ( .A1(G101), .A2(n579), .ZN(n580) );
  XNOR2_X1 U639 ( .A(n581), .B(KEYINPUT65), .ZN(n583) );
  NAND2_X1 U640 ( .A1(G125), .A2(n991), .ZN(n582) );
  NAND2_X1 U641 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U642 ( .A(n584), .B(KEYINPUT66), .ZN(n588) );
  NAND2_X1 U643 ( .A1(G137), .A2(n585), .ZN(n586) );
  XNOR2_X1 U644 ( .A(KEYINPUT67), .B(n586), .ZN(n587) );
  NAND2_X1 U645 ( .A1(n990), .A2(G113), .ZN(n589) );
  NAND2_X1 U646 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U647 ( .A1(G40), .A2(n758), .ZN(n686) );
  XNOR2_X1 U648 ( .A(KEYINPUT95), .B(n686), .ZN(n593) );
  NOR2_X1 U649 ( .A1(G1384), .A2(G164), .ZN(n687) );
  NAND2_X1 U650 ( .A1(n593), .A2(n687), .ZN(n669) );
  NAND2_X1 U651 ( .A1(G1961), .A2(n669), .ZN(n595) );
  INV_X1 U652 ( .A(n669), .ZN(n667) );
  XOR2_X1 U653 ( .A(G2078), .B(KEYINPUT25), .Z(n865) );
  NAND2_X1 U654 ( .A1(n667), .A2(n865), .ZN(n594) );
  NAND2_X1 U655 ( .A1(n595), .A2(n594), .ZN(n652) );
  OR2_X1 U656 ( .A1(G301), .A2(n652), .ZN(n643) );
  NAND2_X1 U657 ( .A1(G53), .A2(n787), .ZN(n597) );
  NAND2_X1 U658 ( .A1(G65), .A2(n788), .ZN(n596) );
  NAND2_X1 U659 ( .A1(n597), .A2(n596), .ZN(n601) );
  NAND2_X1 U660 ( .A1(G91), .A2(n783), .ZN(n599) );
  NAND2_X1 U661 ( .A1(G78), .A2(n784), .ZN(n598) );
  NAND2_X1 U662 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U663 ( .A1(n601), .A2(n600), .ZN(n884) );
  NAND2_X1 U664 ( .A1(n667), .A2(G2072), .ZN(n602) );
  XNOR2_X1 U665 ( .A(n602), .B(KEYINPUT27), .ZN(n604) );
  INV_X1 U666 ( .A(G1956), .ZN(n847) );
  NOR2_X1 U667 ( .A1(n847), .A2(n667), .ZN(n603) );
  NOR2_X1 U668 ( .A1(n604), .A2(n603), .ZN(n606) );
  NOR2_X1 U669 ( .A1(n884), .A2(n606), .ZN(n605) );
  XOR2_X1 U670 ( .A(n605), .B(KEYINPUT28), .Z(n640) );
  NAND2_X1 U671 ( .A1(n884), .A2(n606), .ZN(n638) );
  NAND2_X1 U672 ( .A1(n783), .A2(G81), .ZN(n607) );
  XNOR2_X1 U673 ( .A(n607), .B(KEYINPUT12), .ZN(n609) );
  NAND2_X1 U674 ( .A1(G68), .A2(n784), .ZN(n608) );
  NAND2_X1 U675 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U676 ( .A(n610), .B(KEYINPUT13), .ZN(n612) );
  NAND2_X1 U677 ( .A1(G43), .A2(n787), .ZN(n611) );
  NAND2_X1 U678 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U679 ( .A1(n788), .A2(G56), .ZN(n613) );
  XNOR2_X1 U680 ( .A(n613), .B(KEYINPUT75), .ZN(n614) );
  XNOR2_X1 U681 ( .A(n614), .B(KEYINPUT14), .ZN(n615) );
  NOR2_X1 U682 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U683 ( .A(KEYINPUT76), .B(n617), .Z(n1012) );
  NAND2_X1 U684 ( .A1(G1996), .A2(n667), .ZN(n618) );
  XOR2_X1 U685 ( .A(KEYINPUT26), .B(n618), .Z(n619) );
  NOR2_X1 U686 ( .A1(n1012), .A2(n619), .ZN(n621) );
  NAND2_X1 U687 ( .A1(G1341), .A2(n669), .ZN(n620) );
  NAND2_X1 U688 ( .A1(n621), .A2(n620), .ZN(n634) );
  NAND2_X1 U689 ( .A1(G54), .A2(n787), .ZN(n623) );
  NAND2_X1 U690 ( .A1(G66), .A2(n788), .ZN(n622) );
  NAND2_X1 U691 ( .A1(n623), .A2(n622), .ZN(n627) );
  NAND2_X1 U692 ( .A1(G92), .A2(n783), .ZN(n625) );
  NAND2_X1 U693 ( .A1(G79), .A2(n784), .ZN(n624) );
  NAND2_X1 U694 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U695 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U696 ( .A(n628), .B(KEYINPUT15), .ZN(n1011) );
  NOR2_X1 U697 ( .A1(n634), .A2(n1011), .ZN(n629) );
  XNOR2_X1 U698 ( .A(n629), .B(KEYINPUT97), .ZN(n633) );
  NOR2_X1 U699 ( .A1(n667), .A2(G1348), .ZN(n631) );
  NOR2_X1 U700 ( .A1(G2067), .A2(n669), .ZN(n630) );
  NOR2_X1 U701 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U702 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U703 ( .A1(n634), .A2(n1011), .ZN(n635) );
  NAND2_X1 U704 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U705 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U706 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U707 ( .A(KEYINPUT29), .B(n641), .Z(n642) );
  NAND2_X1 U708 ( .A1(n643), .A2(n642), .ZN(n659) );
  INV_X1 U709 ( .A(G8), .ZN(n668) );
  OR2_X1 U710 ( .A1(n668), .A2(G1966), .ZN(n644) );
  NOR2_X1 U711 ( .A1(n667), .A2(n644), .ZN(n660) );
  NOR2_X1 U712 ( .A1(n669), .A2(G2084), .ZN(n645) );
  XNOR2_X1 U713 ( .A(n645), .B(KEYINPUT96), .ZN(n662) );
  NOR2_X1 U714 ( .A1(n660), .A2(n662), .ZN(n646) );
  NAND2_X1 U715 ( .A1(n646), .A2(G8), .ZN(n648) );
  NOR2_X1 U716 ( .A1(n649), .A2(G168), .ZN(n651) );
  INV_X1 U717 ( .A(KEYINPUT99), .ZN(n650) );
  XNOR2_X1 U718 ( .A(n651), .B(n650), .ZN(n655) );
  NAND2_X1 U719 ( .A1(G301), .A2(n652), .ZN(n653) );
  XOR2_X1 U720 ( .A(KEYINPUT100), .B(n653), .Z(n654) );
  NOR2_X1 U721 ( .A1(n655), .A2(n654), .ZN(n657) );
  NAND2_X1 U722 ( .A1(n659), .A2(n658), .ZN(n666) );
  INV_X1 U723 ( .A(n660), .ZN(n661) );
  NAND2_X1 U724 ( .A1(G8), .A2(n662), .ZN(n663) );
  NAND2_X1 U725 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U726 ( .A(KEYINPUT102), .B(n665), .ZN(n679) );
  NAND2_X1 U727 ( .A1(n666), .A2(G286), .ZN(n674) );
  OR2_X1 U728 ( .A1(n668), .A2(n667), .ZN(n729) );
  NOR2_X1 U729 ( .A1(G1971), .A2(n729), .ZN(n671) );
  NOR2_X1 U730 ( .A1(G2090), .A2(n669), .ZN(n670) );
  NOR2_X1 U731 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U732 ( .A1(G303), .A2(n672), .ZN(n673) );
  NAND2_X1 U733 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U734 ( .A1(n675), .A2(G8), .ZN(n677) );
  XOR2_X1 U735 ( .A(KEYINPUT103), .B(KEYINPUT32), .Z(n676) );
  XNOR2_X1 U736 ( .A(n677), .B(n676), .ZN(n678) );
  NAND2_X1 U737 ( .A1(n679), .A2(n678), .ZN(n726) );
  NOR2_X1 U738 ( .A1(G2090), .A2(G303), .ZN(n680) );
  NAND2_X1 U739 ( .A1(G8), .A2(n680), .ZN(n684) );
  NOR2_X1 U740 ( .A1(G1981), .A2(G305), .ZN(n681) );
  XOR2_X1 U741 ( .A(n681), .B(KEYINPUT24), .Z(n682) );
  NOR2_X1 U742 ( .A1(n729), .A2(n682), .ZN(n718) );
  INV_X1 U743 ( .A(n718), .ZN(n683) );
  AND2_X1 U744 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U745 ( .A1(n726), .A2(n685), .ZN(n721) );
  NOR2_X1 U746 ( .A1(n687), .A2(n686), .ZN(n753) );
  NAND2_X1 U747 ( .A1(G105), .A2(n994), .ZN(n688) );
  XNOR2_X1 U748 ( .A(n688), .B(KEYINPUT38), .ZN(n695) );
  NAND2_X1 U749 ( .A1(G117), .A2(n990), .ZN(n690) );
  NAND2_X1 U750 ( .A1(G141), .A2(n995), .ZN(n689) );
  NAND2_X1 U751 ( .A1(n690), .A2(n689), .ZN(n693) );
  NAND2_X1 U752 ( .A1(n991), .A2(G129), .ZN(n691) );
  XOR2_X1 U753 ( .A(KEYINPUT92), .B(n691), .Z(n692) );
  NOR2_X1 U754 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U755 ( .A1(n695), .A2(n694), .ZN(n983) );
  NAND2_X1 U756 ( .A1(G1996), .A2(n983), .ZN(n696) );
  XOR2_X1 U757 ( .A(KEYINPUT93), .B(n696), .Z(n705) );
  NAND2_X1 U758 ( .A1(G95), .A2(n994), .ZN(n698) );
  NAND2_X1 U759 ( .A1(G131), .A2(n995), .ZN(n697) );
  NAND2_X1 U760 ( .A1(n698), .A2(n697), .ZN(n701) );
  NAND2_X1 U761 ( .A1(G107), .A2(n990), .ZN(n699) );
  XNOR2_X1 U762 ( .A(KEYINPUT91), .B(n699), .ZN(n700) );
  NOR2_X1 U763 ( .A1(n701), .A2(n700), .ZN(n703) );
  NAND2_X1 U764 ( .A1(n991), .A2(G119), .ZN(n702) );
  NAND2_X1 U765 ( .A1(n703), .A2(n702), .ZN(n982) );
  NAND2_X1 U766 ( .A1(G1991), .A2(n982), .ZN(n704) );
  NAND2_X1 U767 ( .A1(n705), .A2(n704), .ZN(n914) );
  NAND2_X1 U768 ( .A1(n753), .A2(n914), .ZN(n706) );
  XOR2_X1 U769 ( .A(KEYINPUT94), .B(n706), .Z(n747) );
  INV_X1 U770 ( .A(n747), .ZN(n717) );
  NAND2_X1 U771 ( .A1(G104), .A2(n994), .ZN(n708) );
  NAND2_X1 U772 ( .A1(G140), .A2(n995), .ZN(n707) );
  NAND2_X1 U773 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U774 ( .A(KEYINPUT34), .B(n709), .ZN(n714) );
  NAND2_X1 U775 ( .A1(G116), .A2(n990), .ZN(n711) );
  NAND2_X1 U776 ( .A1(G128), .A2(n991), .ZN(n710) );
  NAND2_X1 U777 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U778 ( .A(n712), .B(KEYINPUT35), .Z(n713) );
  NOR2_X1 U779 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U780 ( .A(KEYINPUT36), .B(n715), .Z(n716) );
  XOR2_X1 U781 ( .A(KEYINPUT90), .B(n716), .Z(n1003) );
  XNOR2_X1 U782 ( .A(G2067), .B(KEYINPUT37), .ZN(n744) );
  NOR2_X1 U783 ( .A1(n1003), .A2(n744), .ZN(n913) );
  NAND2_X1 U784 ( .A1(n753), .A2(n913), .ZN(n750) );
  NAND2_X1 U785 ( .A1(n717), .A2(n750), .ZN(n733) );
  NOR2_X1 U786 ( .A1(n718), .A2(n729), .ZN(n719) );
  NOR2_X1 U787 ( .A1(n733), .A2(n719), .ZN(n720) );
  NAND2_X1 U788 ( .A1(n721), .A2(n720), .ZN(n741) );
  NOR2_X1 U789 ( .A1(G1976), .A2(G288), .ZN(n894) );
  NOR2_X1 U790 ( .A1(G1971), .A2(G303), .ZN(n722) );
  NOR2_X1 U791 ( .A1(n894), .A2(n722), .ZN(n724) );
  INV_X1 U792 ( .A(KEYINPUT33), .ZN(n723) );
  AND2_X1 U793 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U794 ( .A1(n726), .A2(n725), .ZN(n739) );
  INV_X1 U795 ( .A(n729), .ZN(n727) );
  NAND2_X1 U796 ( .A1(G1976), .A2(G288), .ZN(n892) );
  AND2_X1 U797 ( .A1(n727), .A2(n892), .ZN(n728) );
  OR2_X1 U798 ( .A1(KEYINPUT33), .A2(n728), .ZN(n737) );
  NAND2_X1 U799 ( .A1(n894), .A2(KEYINPUT33), .ZN(n730) );
  NOR2_X1 U800 ( .A1(n730), .A2(n729), .ZN(n732) );
  XOR2_X1 U801 ( .A(G1981), .B(G305), .Z(n902) );
  INV_X1 U802 ( .A(n902), .ZN(n731) );
  NOR2_X1 U803 ( .A1(n732), .A2(n731), .ZN(n735) );
  INV_X1 U804 ( .A(n733), .ZN(n734) );
  AND2_X1 U805 ( .A1(n735), .A2(n734), .ZN(n736) );
  AND2_X1 U806 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U807 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U808 ( .A1(n741), .A2(n740), .ZN(n743) );
  XNOR2_X1 U809 ( .A(G1986), .B(G290), .ZN(n886) );
  NAND2_X1 U810 ( .A1(n886), .A2(n753), .ZN(n742) );
  NAND2_X1 U811 ( .A1(n743), .A2(n742), .ZN(n756) );
  NAND2_X1 U812 ( .A1(n1003), .A2(n744), .ZN(n934) );
  NOR2_X1 U813 ( .A1(G1996), .A2(n983), .ZN(n930) );
  NOR2_X1 U814 ( .A1(G1986), .A2(G290), .ZN(n745) );
  NOR2_X1 U815 ( .A1(G1991), .A2(n982), .ZN(n910) );
  NOR2_X1 U816 ( .A1(n745), .A2(n910), .ZN(n746) );
  NOR2_X1 U817 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U818 ( .A1(n930), .A2(n748), .ZN(n749) );
  XNOR2_X1 U819 ( .A(KEYINPUT39), .B(n749), .ZN(n751) );
  NAND2_X1 U820 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U821 ( .A1(n934), .A2(n752), .ZN(n754) );
  NAND2_X1 U822 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U823 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U824 ( .A(n757), .B(KEYINPUT40), .ZN(G329) );
  BUF_X1 U825 ( .A(n758), .Z(G160) );
  AND2_X1 U826 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U827 ( .A1(G123), .A2(n991), .ZN(n759) );
  XNOR2_X1 U828 ( .A(n759), .B(KEYINPUT18), .ZN(n766) );
  NAND2_X1 U829 ( .A1(G99), .A2(n994), .ZN(n761) );
  NAND2_X1 U830 ( .A1(G135), .A2(n995), .ZN(n760) );
  NAND2_X1 U831 ( .A1(n761), .A2(n760), .ZN(n764) );
  NAND2_X1 U832 ( .A1(n990), .A2(G111), .ZN(n762) );
  XOR2_X1 U833 ( .A(KEYINPUT80), .B(n762), .Z(n763) );
  NOR2_X1 U834 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U835 ( .A1(n766), .A2(n765), .ZN(n985) );
  XNOR2_X1 U836 ( .A(G2096), .B(n985), .ZN(n767) );
  OR2_X1 U837 ( .A1(G2100), .A2(n767), .ZN(G156) );
  INV_X1 U838 ( .A(G860), .ZN(n795) );
  OR2_X1 U839 ( .A1(n795), .A2(n1012), .ZN(G153) );
  INV_X1 U840 ( .A(G69), .ZN(G235) );
  INV_X1 U841 ( .A(G108), .ZN(G238) );
  INV_X1 U842 ( .A(G120), .ZN(G236) );
  INV_X1 U843 ( .A(G132), .ZN(G219) );
  INV_X1 U844 ( .A(G82), .ZN(G220) );
  NAND2_X1 U845 ( .A1(G7), .A2(G661), .ZN(n768) );
  XNOR2_X1 U846 ( .A(n768), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U847 ( .A(KEYINPUT11), .B(KEYINPUT74), .Z(n770) );
  INV_X1 U848 ( .A(G223), .ZN(n823) );
  NAND2_X1 U849 ( .A1(G567), .A2(n823), .ZN(n769) );
  XNOR2_X1 U850 ( .A(n770), .B(n769), .ZN(G234) );
  INV_X1 U851 ( .A(n1011), .ZN(n793) );
  NOR2_X1 U852 ( .A1(n793), .A2(G868), .ZN(n771) );
  XNOR2_X1 U853 ( .A(n771), .B(KEYINPUT77), .ZN(n773) );
  NAND2_X1 U854 ( .A1(G868), .A2(G301), .ZN(n772) );
  NAND2_X1 U855 ( .A1(n773), .A2(n772), .ZN(G284) );
  XOR2_X1 U856 ( .A(n884), .B(KEYINPUT72), .Z(G299) );
  NOR2_X1 U857 ( .A1(G299), .A2(G868), .ZN(n774) );
  XNOR2_X1 U858 ( .A(n774), .B(KEYINPUT78), .ZN(n776) );
  INV_X1 U859 ( .A(G868), .ZN(n805) );
  NOR2_X1 U860 ( .A1(n805), .A2(G286), .ZN(n775) );
  NOR2_X1 U861 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U862 ( .A(KEYINPUT79), .B(n777), .Z(G297) );
  NAND2_X1 U863 ( .A1(n795), .A2(G559), .ZN(n778) );
  NAND2_X1 U864 ( .A1(n778), .A2(n793), .ZN(n779) );
  XNOR2_X1 U865 ( .A(n779), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U866 ( .A1(n1012), .A2(G868), .ZN(n782) );
  NAND2_X1 U867 ( .A1(G868), .A2(n793), .ZN(n780) );
  NOR2_X1 U868 ( .A1(G559), .A2(n780), .ZN(n781) );
  NOR2_X1 U869 ( .A1(n782), .A2(n781), .ZN(G282) );
  NAND2_X1 U870 ( .A1(G93), .A2(n783), .ZN(n786) );
  NAND2_X1 U871 ( .A1(G80), .A2(n784), .ZN(n785) );
  NAND2_X1 U872 ( .A1(n786), .A2(n785), .ZN(n792) );
  NAND2_X1 U873 ( .A1(G55), .A2(n787), .ZN(n790) );
  NAND2_X1 U874 ( .A1(G67), .A2(n788), .ZN(n789) );
  NAND2_X1 U875 ( .A1(n790), .A2(n789), .ZN(n791) );
  OR2_X1 U876 ( .A1(n792), .A2(n791), .ZN(n806) );
  NAND2_X1 U877 ( .A1(G559), .A2(n793), .ZN(n794) );
  XOR2_X1 U878 ( .A(n1012), .B(n794), .Z(n803) );
  NAND2_X1 U879 ( .A1(n795), .A2(n803), .ZN(n796) );
  XNOR2_X1 U880 ( .A(n796), .B(KEYINPUT81), .ZN(n797) );
  XOR2_X1 U881 ( .A(n806), .B(n797), .Z(G145) );
  XOR2_X1 U882 ( .A(KEYINPUT19), .B(n806), .Z(n802) );
  XNOR2_X1 U883 ( .A(G299), .B(G290), .ZN(n798) );
  XNOR2_X1 U884 ( .A(n798), .B(G288), .ZN(n799) );
  XNOR2_X1 U885 ( .A(G166), .B(n799), .ZN(n800) );
  XNOR2_X1 U886 ( .A(n800), .B(G305), .ZN(n801) );
  XNOR2_X1 U887 ( .A(n802), .B(n801), .ZN(n1013) );
  XNOR2_X1 U888 ( .A(n803), .B(n1013), .ZN(n804) );
  NAND2_X1 U889 ( .A1(n804), .A2(G868), .ZN(n808) );
  NAND2_X1 U890 ( .A1(n806), .A2(n805), .ZN(n807) );
  NAND2_X1 U891 ( .A1(n808), .A2(n807), .ZN(G295) );
  NAND2_X1 U892 ( .A1(G2078), .A2(G2084), .ZN(n809) );
  XOR2_X1 U893 ( .A(KEYINPUT20), .B(n809), .Z(n810) );
  NAND2_X1 U894 ( .A1(G2090), .A2(n810), .ZN(n811) );
  XNOR2_X1 U895 ( .A(KEYINPUT21), .B(n811), .ZN(n812) );
  NAND2_X1 U896 ( .A1(n812), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U897 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U898 ( .A(KEYINPUT73), .B(G57), .ZN(G237) );
  NOR2_X1 U899 ( .A1(G220), .A2(G219), .ZN(n813) );
  XOR2_X1 U900 ( .A(KEYINPUT22), .B(n813), .Z(n814) );
  NOR2_X1 U901 ( .A1(G218), .A2(n814), .ZN(n815) );
  XOR2_X1 U902 ( .A(KEYINPUT85), .B(n815), .Z(n816) );
  NAND2_X1 U903 ( .A1(G96), .A2(n816), .ZN(n949) );
  NAND2_X1 U904 ( .A1(n949), .A2(G2106), .ZN(n821) );
  NOR2_X1 U905 ( .A1(G237), .A2(G236), .ZN(n818) );
  NOR2_X1 U906 ( .A1(G238), .A2(G235), .ZN(n817) );
  NAND2_X1 U907 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U908 ( .A(KEYINPUT86), .B(n819), .ZN(n950) );
  NAND2_X1 U909 ( .A1(n950), .A2(G567), .ZN(n820) );
  NAND2_X1 U910 ( .A1(n821), .A2(n820), .ZN(n981) );
  NAND2_X1 U911 ( .A1(G483), .A2(G661), .ZN(n822) );
  NOR2_X1 U912 ( .A1(n981), .A2(n822), .ZN(n826) );
  NAND2_X1 U913 ( .A1(n826), .A2(G36), .ZN(G176) );
  NAND2_X1 U914 ( .A1(G2106), .A2(n823), .ZN(G217) );
  AND2_X1 U915 ( .A1(G15), .A2(G2), .ZN(n824) );
  NAND2_X1 U916 ( .A1(G661), .A2(n824), .ZN(G259) );
  NAND2_X1 U917 ( .A1(G3), .A2(G1), .ZN(n825) );
  XNOR2_X1 U918 ( .A(KEYINPUT106), .B(n825), .ZN(n827) );
  NAND2_X1 U919 ( .A1(n827), .A2(n826), .ZN(G188) );
  NAND2_X1 U921 ( .A1(G124), .A2(n991), .ZN(n828) );
  XNOR2_X1 U922 ( .A(n828), .B(KEYINPUT44), .ZN(n829) );
  XNOR2_X1 U923 ( .A(KEYINPUT110), .B(n829), .ZN(n832) );
  NAND2_X1 U924 ( .A1(G112), .A2(n990), .ZN(n830) );
  XOR2_X1 U925 ( .A(KEYINPUT111), .B(n830), .Z(n831) );
  NAND2_X1 U926 ( .A1(n832), .A2(n831), .ZN(n836) );
  NAND2_X1 U927 ( .A1(G100), .A2(n994), .ZN(n834) );
  NAND2_X1 U928 ( .A1(G136), .A2(n995), .ZN(n833) );
  NAND2_X1 U929 ( .A1(n834), .A2(n833), .ZN(n835) );
  NOR2_X1 U930 ( .A1(n836), .A2(n835), .ZN(G162) );
  XOR2_X1 U931 ( .A(G1966), .B(G21), .Z(n846) );
  XNOR2_X1 U932 ( .A(G1986), .B(KEYINPUT126), .ZN(n837) );
  XNOR2_X1 U933 ( .A(n837), .B(G24), .ZN(n843) );
  XNOR2_X1 U934 ( .A(G1971), .B(G22), .ZN(n838) );
  XNOR2_X1 U935 ( .A(n838), .B(KEYINPUT124), .ZN(n840) );
  XNOR2_X1 U936 ( .A(G23), .B(G1976), .ZN(n839) );
  NOR2_X1 U937 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U938 ( .A(n841), .B(KEYINPUT125), .ZN(n842) );
  NOR2_X1 U939 ( .A1(n843), .A2(n842), .ZN(n844) );
  XNOR2_X1 U940 ( .A(KEYINPUT58), .B(n844), .ZN(n845) );
  NAND2_X1 U941 ( .A1(n846), .A2(n845), .ZN(n859) );
  XOR2_X1 U942 ( .A(G1961), .B(G5), .Z(n857) );
  XNOR2_X1 U943 ( .A(G20), .B(n847), .ZN(n851) );
  XNOR2_X1 U944 ( .A(G1341), .B(G19), .ZN(n849) );
  XNOR2_X1 U945 ( .A(G1981), .B(G6), .ZN(n848) );
  NOR2_X1 U946 ( .A1(n849), .A2(n848), .ZN(n850) );
  NAND2_X1 U947 ( .A1(n851), .A2(n850), .ZN(n854) );
  XOR2_X1 U948 ( .A(KEYINPUT59), .B(G1348), .Z(n852) );
  XNOR2_X1 U949 ( .A(G4), .B(n852), .ZN(n853) );
  NOR2_X1 U950 ( .A1(n854), .A2(n853), .ZN(n855) );
  XNOR2_X1 U951 ( .A(n855), .B(KEYINPUT60), .ZN(n856) );
  NAND2_X1 U952 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U953 ( .A1(n859), .A2(n858), .ZN(n860) );
  XNOR2_X1 U954 ( .A(n860), .B(KEYINPUT61), .ZN(n862) );
  XNOR2_X1 U955 ( .A(G16), .B(KEYINPUT123), .ZN(n861) );
  NAND2_X1 U956 ( .A1(n862), .A2(n861), .ZN(n947) );
  INV_X1 U957 ( .A(KEYINPUT55), .ZN(n939) );
  XNOR2_X1 U958 ( .A(G2090), .B(G35), .ZN(n876) );
  XNOR2_X1 U959 ( .A(G2067), .B(G26), .ZN(n864) );
  XNOR2_X1 U960 ( .A(G2072), .B(G33), .ZN(n863) );
  NOR2_X1 U961 ( .A1(n864), .A2(n863), .ZN(n869) );
  XNOR2_X1 U962 ( .A(G1996), .B(G32), .ZN(n867) );
  XNOR2_X1 U963 ( .A(G27), .B(n865), .ZN(n866) );
  NOR2_X1 U964 ( .A1(n867), .A2(n866), .ZN(n868) );
  NAND2_X1 U965 ( .A1(n869), .A2(n868), .ZN(n873) );
  XOR2_X1 U966 ( .A(G1991), .B(G25), .Z(n870) );
  NAND2_X1 U967 ( .A1(n870), .A2(G28), .ZN(n871) );
  XOR2_X1 U968 ( .A(KEYINPUT119), .B(n871), .Z(n872) );
  NOR2_X1 U969 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U970 ( .A(KEYINPUT53), .B(n874), .ZN(n875) );
  NOR2_X1 U971 ( .A1(n876), .A2(n875), .ZN(n879) );
  XOR2_X1 U972 ( .A(G2084), .B(KEYINPUT54), .Z(n877) );
  XNOR2_X1 U973 ( .A(G34), .B(n877), .ZN(n878) );
  NAND2_X1 U974 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U975 ( .A(n939), .B(n880), .ZN(n882) );
  INV_X1 U976 ( .A(G29), .ZN(n881) );
  NAND2_X1 U977 ( .A1(n882), .A2(n881), .ZN(n883) );
  NAND2_X1 U978 ( .A1(G11), .A2(n883), .ZN(n945) );
  XNOR2_X1 U979 ( .A(G16), .B(KEYINPUT56), .ZN(n908) );
  XNOR2_X1 U980 ( .A(n884), .B(G1956), .ZN(n888) );
  XNOR2_X1 U981 ( .A(G1348), .B(n1011), .ZN(n885) );
  NOR2_X1 U982 ( .A1(n886), .A2(n885), .ZN(n887) );
  NAND2_X1 U983 ( .A1(n888), .A2(n887), .ZN(n890) );
  XNOR2_X1 U984 ( .A(G1341), .B(n1012), .ZN(n889) );
  NOR2_X1 U985 ( .A1(n890), .A2(n889), .ZN(n898) );
  XOR2_X1 U986 ( .A(G1971), .B(G303), .Z(n891) );
  XNOR2_X1 U987 ( .A(n891), .B(KEYINPUT120), .ZN(n893) );
  NAND2_X1 U988 ( .A1(n893), .A2(n892), .ZN(n895) );
  NOR2_X1 U989 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U990 ( .A(KEYINPUT121), .B(n896), .Z(n897) );
  NAND2_X1 U991 ( .A1(n898), .A2(n897), .ZN(n900) );
  XNOR2_X1 U992 ( .A(G1961), .B(G301), .ZN(n899) );
  NOR2_X1 U993 ( .A1(n900), .A2(n899), .ZN(n901) );
  XNOR2_X1 U994 ( .A(KEYINPUT122), .B(n901), .ZN(n906) );
  XNOR2_X1 U995 ( .A(G168), .B(G1966), .ZN(n903) );
  NAND2_X1 U996 ( .A1(n903), .A2(n902), .ZN(n904) );
  XNOR2_X1 U997 ( .A(KEYINPUT57), .B(n904), .ZN(n905) );
  NAND2_X1 U998 ( .A1(n906), .A2(n905), .ZN(n907) );
  NAND2_X1 U999 ( .A1(n908), .A2(n907), .ZN(n943) );
  XOR2_X1 U1000 ( .A(G2084), .B(G160), .Z(n909) );
  NOR2_X1 U1001 ( .A1(n910), .A2(n909), .ZN(n911) );
  NAND2_X1 U1002 ( .A1(n911), .A2(n985), .ZN(n912) );
  XNOR2_X1 U1003 ( .A(KEYINPUT117), .B(n912), .ZN(n916) );
  NOR2_X1 U1004 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1005 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1006 ( .A(KEYINPUT118), .B(n917), .ZN(n937) );
  NAND2_X1 U1007 ( .A1(G103), .A2(n994), .ZN(n919) );
  NAND2_X1 U1008 ( .A1(G139), .A2(n995), .ZN(n918) );
  NAND2_X1 U1009 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1010 ( .A(KEYINPUT113), .B(n920), .Z(n925) );
  NAND2_X1 U1011 ( .A1(G115), .A2(n990), .ZN(n922) );
  NAND2_X1 U1012 ( .A1(G127), .A2(n991), .ZN(n921) );
  NAND2_X1 U1013 ( .A1(n922), .A2(n921), .ZN(n923) );
  XOR2_X1 U1014 ( .A(KEYINPUT47), .B(n923), .Z(n924) );
  NOR2_X1 U1015 ( .A1(n925), .A2(n924), .ZN(n1007) );
  XOR2_X1 U1016 ( .A(G2072), .B(n1007), .Z(n927) );
  XOR2_X1 U1017 ( .A(G164), .B(G2078), .Z(n926) );
  NOR2_X1 U1018 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1019 ( .A(KEYINPUT50), .B(n928), .Z(n933) );
  XOR2_X1 U1020 ( .A(G2090), .B(G162), .Z(n929) );
  NOR2_X1 U1021 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1022 ( .A(KEYINPUT51), .B(n931), .ZN(n932) );
  NOR2_X1 U1023 ( .A1(n933), .A2(n932), .ZN(n935) );
  NAND2_X1 U1024 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1025 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1026 ( .A(KEYINPUT52), .B(n938), .ZN(n940) );
  NAND2_X1 U1027 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1028 ( .A1(n941), .A2(G29), .ZN(n942) );
  NAND2_X1 U1029 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1030 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1031 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1032 ( .A(KEYINPUT62), .B(n948), .Z(G311) );
  XNOR2_X1 U1033 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1034 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1035 ( .A1(n950), .A2(n949), .ZN(G325) );
  INV_X1 U1036 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U1037 ( .A(G1348), .B(G2454), .ZN(n951) );
  XNOR2_X1 U1038 ( .A(n951), .B(G2430), .ZN(n952) );
  XNOR2_X1 U1039 ( .A(n952), .B(G1341), .ZN(n958) );
  XOR2_X1 U1040 ( .A(G2443), .B(G2427), .Z(n954) );
  XNOR2_X1 U1041 ( .A(G2438), .B(G2446), .ZN(n953) );
  XNOR2_X1 U1042 ( .A(n954), .B(n953), .ZN(n956) );
  XOR2_X1 U1043 ( .A(G2451), .B(G2435), .Z(n955) );
  XNOR2_X1 U1044 ( .A(n956), .B(n955), .ZN(n957) );
  XNOR2_X1 U1045 ( .A(n958), .B(n957), .ZN(n959) );
  NAND2_X1 U1046 ( .A1(n959), .A2(G14), .ZN(n960) );
  XNOR2_X1 U1047 ( .A(KEYINPUT104), .B(n960), .ZN(n1021) );
  XNOR2_X1 U1048 ( .A(n1021), .B(KEYINPUT105), .ZN(G401) );
  XOR2_X1 U1049 ( .A(KEYINPUT109), .B(G2474), .Z(n962) );
  XNOR2_X1 U1050 ( .A(G1986), .B(G1976), .ZN(n961) );
  XNOR2_X1 U1051 ( .A(n962), .B(n961), .ZN(n963) );
  XOR2_X1 U1052 ( .A(n963), .B(G1956), .Z(n965) );
  XNOR2_X1 U1053 ( .A(G1996), .B(G1991), .ZN(n964) );
  XNOR2_X1 U1054 ( .A(n965), .B(n964), .ZN(n969) );
  XOR2_X1 U1055 ( .A(KEYINPUT108), .B(KEYINPUT41), .Z(n967) );
  XNOR2_X1 U1056 ( .A(G1971), .B(G1961), .ZN(n966) );
  XNOR2_X1 U1057 ( .A(n967), .B(n966), .ZN(n968) );
  XOR2_X1 U1058 ( .A(n969), .B(n968), .Z(n971) );
  XNOR2_X1 U1059 ( .A(G1966), .B(G1981), .ZN(n970) );
  XNOR2_X1 U1060 ( .A(n971), .B(n970), .ZN(G229) );
  XOR2_X1 U1061 ( .A(KEYINPUT42), .B(G2084), .Z(n973) );
  XNOR2_X1 U1062 ( .A(G2067), .B(G2078), .ZN(n972) );
  XNOR2_X1 U1063 ( .A(n973), .B(n972), .ZN(n974) );
  XOR2_X1 U1064 ( .A(n974), .B(G2678), .Z(n976) );
  XNOR2_X1 U1065 ( .A(G2072), .B(KEYINPUT107), .ZN(n975) );
  XNOR2_X1 U1066 ( .A(n976), .B(n975), .ZN(n980) );
  XOR2_X1 U1067 ( .A(G2100), .B(G2096), .Z(n978) );
  XNOR2_X1 U1068 ( .A(G2090), .B(KEYINPUT43), .ZN(n977) );
  XNOR2_X1 U1069 ( .A(n978), .B(n977), .ZN(n979) );
  XOR2_X1 U1070 ( .A(n980), .B(n979), .Z(G227) );
  INV_X1 U1071 ( .A(n981), .ZN(G319) );
  XOR2_X1 U1072 ( .A(n983), .B(n982), .Z(n984) );
  XNOR2_X1 U1073 ( .A(n985), .B(n984), .ZN(n989) );
  XOR2_X1 U1074 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n987) );
  XNOR2_X1 U1075 ( .A(G162), .B(KEYINPUT114), .ZN(n986) );
  XNOR2_X1 U1076 ( .A(n987), .B(n986), .ZN(n988) );
  XOR2_X1 U1077 ( .A(n989), .B(n988), .Z(n1005) );
  NAND2_X1 U1078 ( .A1(G118), .A2(n990), .ZN(n993) );
  NAND2_X1 U1079 ( .A1(G130), .A2(n991), .ZN(n992) );
  NAND2_X1 U1080 ( .A1(n993), .A2(n992), .ZN(n1001) );
  NAND2_X1 U1081 ( .A1(G106), .A2(n994), .ZN(n997) );
  NAND2_X1 U1082 ( .A1(G142), .A2(n995), .ZN(n996) );
  NAND2_X1 U1083 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1084 ( .A(KEYINPUT45), .B(n998), .Z(n999) );
  XNOR2_X1 U1085 ( .A(KEYINPUT112), .B(n999), .ZN(n1000) );
  NOR2_X1 U1086 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1087 ( .A(n1003), .B(n1002), .ZN(n1004) );
  XNOR2_X1 U1088 ( .A(n1005), .B(n1004), .ZN(n1006) );
  XOR2_X1 U1089 ( .A(n1007), .B(n1006), .Z(n1008) );
  XNOR2_X1 U1090 ( .A(G164), .B(n1008), .ZN(n1009) );
  XOR2_X1 U1091 ( .A(n1009), .B(G160), .Z(n1010) );
  NOR2_X1 U1092 ( .A1(G37), .A2(n1010), .ZN(G395) );
  XNOR2_X1 U1093 ( .A(KEYINPUT115), .B(n1011), .ZN(n1016) );
  XNOR2_X1 U1094 ( .A(G171), .B(n1012), .ZN(n1014) );
  XNOR2_X1 U1095 ( .A(n1014), .B(n1013), .ZN(n1015) );
  XNOR2_X1 U1096 ( .A(n1016), .B(n1015), .ZN(n1017) );
  XNOR2_X1 U1097 ( .A(n1017), .B(G286), .ZN(n1018) );
  NOR2_X1 U1098 ( .A1(G37), .A2(n1018), .ZN(G397) );
  XNOR2_X1 U1099 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n1020) );
  NOR2_X1 U1100 ( .A1(G229), .A2(G227), .ZN(n1019) );
  XNOR2_X1 U1101 ( .A(n1020), .B(n1019), .ZN(n1023) );
  NAND2_X1 U1102 ( .A1(G319), .A2(n1021), .ZN(n1022) );
  NOR2_X1 U1103 ( .A1(n1023), .A2(n1022), .ZN(n1025) );
  NOR2_X1 U1104 ( .A1(G395), .A2(G397), .ZN(n1024) );
  NAND2_X1 U1105 ( .A1(n1025), .A2(n1024), .ZN(G225) );
  INV_X1 U1106 ( .A(G225), .ZN(G308) );
endmodule

