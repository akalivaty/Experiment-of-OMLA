

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742;

  XNOR2_X2 U382 ( .A(n526), .B(n525), .ZN(n710) );
  INV_X2 U383 ( .A(G953), .ZN(n734) );
  NAND2_X1 U384 ( .A1(n656), .A2(n655), .ZN(n510) );
  XOR2_X1 U385 ( .A(G146), .B(G125), .Z(n408) );
  INV_X1 U386 ( .A(KEYINPUT3), .ZN(n384) );
  XNOR2_X1 U387 ( .A(G113), .B(G119), .ZN(n382) );
  OR2_X1 U388 ( .A1(n588), .A2(n372), .ZN(n732) );
  NAND2_X1 U389 ( .A1(n739), .A2(n635), .ZN(n501) );
  NAND2_X1 U390 ( .A1(n517), .A2(n478), .ZN(n381) );
  XNOR2_X1 U391 ( .A(n466), .B(n465), .ZN(n545) );
  XNOR2_X1 U392 ( .A(n383), .B(n382), .ZN(n439) );
  XNOR2_X1 U393 ( .A(n384), .B(KEYINPUT91), .ZN(n383) );
  XNOR2_X1 U394 ( .A(G143), .B(G128), .ZN(n424) );
  XNOR2_X1 U395 ( .A(G131), .B(G134), .ZN(n725) );
  XNOR2_X2 U396 ( .A(n399), .B(n398), .ZN(n552) );
  XNOR2_X1 U397 ( .A(n726), .B(G101), .ZN(n445) );
  NOR2_X1 U398 ( .A1(n545), .A2(n544), .ZN(n567) );
  XNOR2_X1 U399 ( .A(n547), .B(KEYINPUT28), .ZN(n558) );
  NAND2_X1 U400 ( .A1(n567), .A2(n546), .ZN(n547) );
  XOR2_X1 U401 ( .A(KEYINPUT10), .B(n408), .Z(n450) );
  NOR2_X1 U402 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U403 ( .A(n368), .B(n367), .ZN(n601) );
  INV_X1 U404 ( .A(n445), .ZN(n367) );
  XNOR2_X1 U405 ( .A(n450), .B(n409), .ZN(n410) );
  XNOR2_X1 U406 ( .A(G140), .B(KEYINPUT97), .ZN(n409) );
  XNOR2_X1 U407 ( .A(G143), .B(G113), .ZN(n407) );
  INV_X1 U408 ( .A(KEYINPUT18), .ZN(n388) );
  NAND2_X1 U409 ( .A1(n362), .A2(n376), .ZN(n375) );
  NAND2_X1 U410 ( .A1(n552), .A2(n670), .ZN(n570) );
  AND2_X1 U411 ( .A1(n539), .A2(n538), .ZN(n553) );
  NOR2_X1 U412 ( .A1(n536), .A2(n544), .ZN(n539) );
  XNOR2_X1 U413 ( .A(n570), .B(KEYINPUT19), .ZN(n557) );
  XNOR2_X1 U414 ( .A(n660), .B(n479), .ZN(n546) );
  XNOR2_X1 U415 ( .A(n444), .B(n441), .ZN(n370) );
  XNOR2_X1 U416 ( .A(KEYINPUT30), .B(KEYINPUT108), .ZN(n527) );
  NAND2_X1 U417 ( .A1(n373), .A2(n650), .ZN(n372) );
  XNOR2_X1 U418 ( .A(G128), .B(G119), .ZN(n452) );
  NOR2_X1 U419 ( .A1(n710), .A2(n598), .ZN(n693) );
  OR2_X1 U420 ( .A1(n588), .A2(n371), .ZN(n598) );
  NAND2_X1 U421 ( .A1(n373), .A2(n597), .ZN(n371) );
  NAND2_X1 U422 ( .A1(n374), .A2(n670), .ZN(n582) );
  INV_X1 U423 ( .A(n556), .ZN(n548) );
  NAND2_X1 U424 ( .A1(n557), .A2(n363), .ZN(n385) );
  XNOR2_X1 U425 ( .A(n463), .B(n462), .ZN(n466) );
  XNOR2_X1 U426 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U427 ( .A(n446), .B(G472), .ZN(n447) );
  XNOR2_X1 U428 ( .A(n361), .B(n415), .ZN(n416) );
  BUF_X1 U429 ( .A(n621), .Z(n705) );
  XNOR2_X1 U430 ( .A(n391), .B(n390), .ZN(n392) );
  AND2_X1 U431 ( .A1(n698), .A2(n734), .ZN(n380) );
  XNOR2_X1 U432 ( .A(n375), .B(KEYINPUT110), .ZN(n569) );
  XOR2_X1 U433 ( .A(n560), .B(KEYINPUT78), .Z(n640) );
  OR2_X1 U434 ( .A1(n514), .A2(n513), .ZN(n645) );
  XNOR2_X1 U435 ( .A(n378), .B(n377), .ZN(G75) );
  INV_X1 U436 ( .A(KEYINPUT53), .ZN(n377) );
  OR2_X1 U437 ( .A1(n694), .A2(n379), .ZN(n378) );
  NAND2_X1 U438 ( .A1(n360), .A2(n380), .ZN(n379) );
  INV_X1 U439 ( .A(n642), .ZN(n376) );
  OR2_X1 U440 ( .A1(n687), .A2(n686), .ZN(n360) );
  XOR2_X1 U441 ( .A(n413), .B(n412), .Z(n361) );
  XNOR2_X1 U442 ( .A(KEYINPUT105), .B(n568), .ZN(n362) );
  OR2_X1 U443 ( .A1(n533), .A2(n403), .ZN(n363) );
  XOR2_X1 U444 ( .A(n405), .B(n404), .Z(n364) );
  XOR2_X1 U445 ( .A(n601), .B(KEYINPUT62), .Z(n365) );
  XOR2_X1 U446 ( .A(KEYINPUT48), .B(KEYINPUT86), .Z(n366) );
  NOR2_X1 U447 ( .A1(n601), .A2(G902), .ZN(n448) );
  XNOR2_X1 U448 ( .A(n370), .B(n369), .ZN(n368) );
  XNOR2_X1 U449 ( .A(n439), .B(n472), .ZN(n369) );
  INV_X1 U450 ( .A(n738), .ZN(n373) );
  INV_X1 U451 ( .A(n375), .ZN(n374) );
  XNOR2_X2 U452 ( .A(n381), .B(KEYINPUT32), .ZN(n739) );
  NOR2_X2 U453 ( .A1(n482), .A2(n566), .ZN(n517) );
  NAND2_X1 U454 ( .A1(n511), .A2(n437), .ZN(n438) );
  XNOR2_X2 U455 ( .A(n385), .B(n364), .ZN(n511) );
  AND2_X2 U456 ( .A1(n600), .A2(n599), .ZN(n621) );
  NAND2_X1 U457 ( .A1(n524), .A2(n523), .ZN(n526) );
  INV_X1 U458 ( .A(KEYINPUT76), .ZN(n390) );
  INV_X1 U459 ( .A(KEYINPUT25), .ZN(n460) );
  XNOR2_X1 U460 ( .A(n393), .B(n392), .ZN(n394) );
  NOR2_X1 U461 ( .A1(n677), .A2(n674), .ZN(n543) );
  INV_X1 U462 ( .A(KEYINPUT66), .ZN(n404) );
  INV_X1 U463 ( .A(n693), .ZN(n599) );
  INV_X1 U464 ( .A(KEYINPUT102), .ZN(n479) );
  XNOR2_X1 U465 ( .A(n417), .B(n416), .ZN(n624) );
  NOR2_X1 U466 ( .A1(n558), .A2(n548), .ZN(n549) );
  INV_X1 U467 ( .A(n709), .ZN(n604) );
  XNOR2_X1 U468 ( .A(n439), .B(KEYINPUT16), .ZN(n387) );
  XOR2_X1 U469 ( .A(G116), .B(G107), .Z(n420) );
  XOR2_X1 U470 ( .A(G122), .B(G104), .Z(n406) );
  XOR2_X1 U471 ( .A(n420), .B(n406), .Z(n386) );
  XNOR2_X1 U472 ( .A(n387), .B(n386), .ZN(n716) );
  XNOR2_X1 U473 ( .A(n408), .B(KEYINPUT17), .ZN(n389) );
  XNOR2_X1 U474 ( .A(n389), .B(n388), .ZN(n393) );
  NAND2_X1 U475 ( .A1(G224), .A2(n734), .ZN(n391) );
  XNOR2_X1 U476 ( .A(n716), .B(n394), .ZN(n397) );
  XNOR2_X1 U477 ( .A(n424), .B(KEYINPUT4), .ZN(n726) );
  XNOR2_X1 U478 ( .A(KEYINPUT73), .B(KEYINPUT90), .ZN(n395) );
  XNOR2_X1 U479 ( .A(n395), .B(G110), .ZN(n717) );
  XNOR2_X1 U480 ( .A(n717), .B(KEYINPUT68), .ZN(n396) );
  XNOR2_X1 U481 ( .A(n445), .B(n396), .ZN(n474) );
  XNOR2_X1 U482 ( .A(n397), .B(n474), .ZN(n611) );
  XNOR2_X1 U483 ( .A(G902), .B(KEYINPUT15), .ZN(n592) );
  NAND2_X1 U484 ( .A1(n611), .A2(n592), .ZN(n399) );
  OR2_X1 U485 ( .A1(G237), .A2(G902), .ZN(n400) );
  AND2_X1 U486 ( .A1(G210), .A2(n400), .ZN(n398) );
  NAND2_X1 U487 ( .A1(G214), .A2(n400), .ZN(n670) );
  NAND2_X1 U488 ( .A1(G234), .A2(G237), .ZN(n401) );
  XNOR2_X1 U489 ( .A(n401), .B(KEYINPUT14), .ZN(n402) );
  NAND2_X1 U490 ( .A1(G952), .A2(n402), .ZN(n687) );
  NOR2_X1 U491 ( .A1(G953), .A2(n687), .ZN(n533) );
  NAND2_X1 U492 ( .A1(G902), .A2(n402), .ZN(n529) );
  OR2_X1 U493 ( .A1(n734), .A2(G898), .ZN(n722) );
  NOR2_X1 U494 ( .A1(n529), .A2(n722), .ZN(n403) );
  INV_X1 U495 ( .A(KEYINPUT0), .ZN(n405) );
  XNOR2_X1 U496 ( .A(KEYINPUT13), .B(G475), .ZN(n419) );
  XNOR2_X1 U497 ( .A(n407), .B(n406), .ZN(n411) );
  XOR2_X1 U498 ( .A(n411), .B(n410), .Z(n417) );
  XOR2_X1 U499 ( .A(KEYINPUT98), .B(KEYINPUT12), .Z(n413) );
  XNOR2_X1 U500 ( .A(G131), .B(KEYINPUT11), .ZN(n412) );
  NOR2_X1 U501 ( .A1(G237), .A2(G953), .ZN(n414) );
  XNOR2_X1 U502 ( .A(n414), .B(KEYINPUT74), .ZN(n440) );
  NAND2_X1 U503 ( .A1(G214), .A2(n440), .ZN(n415) );
  NOR2_X1 U504 ( .A1(G902), .A2(n624), .ZN(n418) );
  XNOR2_X1 U505 ( .A(n419), .B(n418), .ZN(n514) );
  INV_X1 U506 ( .A(n514), .ZN(n432) );
  XNOR2_X1 U507 ( .A(n420), .B(KEYINPUT7), .ZN(n430) );
  NAND2_X1 U508 ( .A1(n734), .A2(G234), .ZN(n422) );
  XNOR2_X1 U509 ( .A(KEYINPUT67), .B(KEYINPUT8), .ZN(n421) );
  XNOR2_X1 U510 ( .A(n422), .B(n421), .ZN(n451) );
  NAND2_X1 U511 ( .A1(n451), .A2(G217), .ZN(n428) );
  XNOR2_X1 U512 ( .A(KEYINPUT9), .B(KEYINPUT99), .ZN(n423) );
  XNOR2_X1 U513 ( .A(n424), .B(n423), .ZN(n426) );
  XNOR2_X1 U514 ( .A(G134), .B(G122), .ZN(n425) );
  XNOR2_X1 U515 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U516 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U517 ( .A(n430), .B(n429), .ZN(n706) );
  NOR2_X1 U518 ( .A1(G902), .A2(n706), .ZN(n431) );
  XNOR2_X1 U519 ( .A(G478), .B(n431), .ZN(n513) );
  NAND2_X1 U520 ( .A1(n432), .A2(n513), .ZN(n674) );
  NAND2_X1 U521 ( .A1(G234), .A2(n592), .ZN(n433) );
  XNOR2_X1 U522 ( .A(KEYINPUT20), .B(n433), .ZN(n464) );
  NAND2_X1 U523 ( .A1(n464), .A2(G221), .ZN(n435) );
  INV_X1 U524 ( .A(KEYINPUT21), .ZN(n434) );
  XNOR2_X1 U525 ( .A(n435), .B(n434), .ZN(n651) );
  INV_X1 U526 ( .A(n651), .ZN(n436) );
  NOR2_X1 U527 ( .A1(n674), .A2(n436), .ZN(n437) );
  XNOR2_X1 U528 ( .A(n438), .B(KEYINPUT22), .ZN(n482) );
  XNOR2_X1 U529 ( .A(n725), .B(G146), .ZN(n472) );
  NAND2_X1 U530 ( .A1(G210), .A2(n440), .ZN(n441) );
  XOR2_X1 U531 ( .A(KEYINPUT72), .B(KEYINPUT5), .Z(n443) );
  XNOR2_X1 U532 ( .A(G137), .B(G116), .ZN(n442) );
  XNOR2_X1 U533 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U534 ( .A(KEYINPUT70), .B(KEYINPUT96), .ZN(n446) );
  XNOR2_X2 U535 ( .A(n448), .B(n447), .ZN(n660) );
  XNOR2_X1 U536 ( .A(KEYINPUT100), .B(KEYINPUT6), .ZN(n449) );
  XNOR2_X1 U537 ( .A(n660), .B(n449), .ZN(n566) );
  XNOR2_X1 U538 ( .A(G140), .B(G137), .ZN(n469) );
  XNOR2_X1 U539 ( .A(n450), .B(n469), .ZN(n728) );
  NAND2_X1 U540 ( .A1(n451), .A2(G221), .ZN(n453) );
  XNOR2_X1 U541 ( .A(n453), .B(n452), .ZN(n458) );
  XOR2_X1 U542 ( .A(KEYINPUT93), .B(KEYINPUT83), .Z(n455) );
  XNOR2_X1 U543 ( .A(G110), .B(KEYINPUT24), .ZN(n454) );
  XNOR2_X1 U544 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U545 ( .A(n456), .B(KEYINPUT23), .Z(n457) );
  XNOR2_X1 U546 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U547 ( .A(n728), .B(n459), .ZN(n617) );
  NOR2_X1 U548 ( .A1(G902), .A2(n617), .ZN(n463) );
  XNOR2_X1 U549 ( .A(KEYINPUT94), .B(KEYINPUT75), .ZN(n461) );
  NAND2_X1 U550 ( .A1(n464), .A2(G217), .ZN(n465) );
  XOR2_X1 U551 ( .A(KEYINPUT101), .B(n545), .Z(n652) );
  XNOR2_X1 U552 ( .A(G107), .B(G104), .ZN(n468) );
  NAND2_X1 U553 ( .A1(n734), .A2(G227), .ZN(n467) );
  XNOR2_X1 U554 ( .A(n468), .B(n467), .ZN(n470) );
  XNOR2_X1 U555 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U556 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U557 ( .A(n474), .B(n473), .ZN(n701) );
  OR2_X1 U558 ( .A1(n701), .A2(G902), .ZN(n476) );
  INV_X1 U559 ( .A(G469), .ZN(n475) );
  XNOR2_X1 U560 ( .A(n476), .B(n475), .ZN(n505) );
  XNOR2_X1 U561 ( .A(n505), .B(KEYINPUT1), .ZN(n518) );
  XNOR2_X1 U562 ( .A(n518), .B(KEYINPUT89), .ZN(n572) );
  INV_X1 U563 ( .A(n572), .ZN(n477) );
  NOR2_X1 U564 ( .A1(n652), .A2(n477), .ZN(n478) );
  NOR2_X1 U565 ( .A1(n546), .A2(n545), .ZN(n480) );
  NAND2_X1 U566 ( .A1(n480), .A2(n518), .ZN(n481) );
  OR2_X1 U567 ( .A1(n482), .A2(n481), .ZN(n635) );
  XNOR2_X1 U568 ( .A(n501), .B(KEYINPUT87), .ZN(n493) );
  AND2_X1 U569 ( .A1(n545), .A2(n651), .ZN(n656) );
  INV_X1 U570 ( .A(n518), .ZN(n655) );
  XNOR2_X1 U571 ( .A(n510), .B(KEYINPUT103), .ZN(n483) );
  NAND2_X1 U572 ( .A1(n483), .A2(n566), .ZN(n487) );
  XNOR2_X1 U573 ( .A(KEYINPUT88), .B(KEYINPUT33), .ZN(n485) );
  INV_X1 U574 ( .A(KEYINPUT69), .ZN(n484) );
  XNOR2_X1 U575 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U576 ( .A(n487), .B(n486), .ZN(n681) );
  XNOR2_X1 U577 ( .A(n511), .B(KEYINPUT92), .ZN(n504) );
  NAND2_X1 U578 ( .A1(n681), .A2(n504), .ZN(n488) );
  XNOR2_X1 U579 ( .A(n488), .B(KEYINPUT34), .ZN(n490) );
  INV_X1 U580 ( .A(n513), .ZN(n489) );
  NAND2_X1 U581 ( .A1(n514), .A2(n489), .ZN(n555) );
  OR2_X1 U582 ( .A1(n490), .A2(n555), .ZN(n492) );
  XNOR2_X1 U583 ( .A(KEYINPUT77), .B(KEYINPUT35), .ZN(n491) );
  XNOR2_X2 U584 ( .A(n492), .B(n491), .ZN(n608) );
  NAND2_X1 U585 ( .A1(n493), .A2(n608), .ZN(n496) );
  INV_X1 U586 ( .A(KEYINPUT44), .ZN(n494) );
  AND2_X1 U587 ( .A1(n494), .A2(KEYINPUT64), .ZN(n495) );
  NAND2_X1 U588 ( .A1(n496), .A2(n495), .ZN(n500) );
  NAND2_X1 U589 ( .A1(n501), .A2(KEYINPUT64), .ZN(n497) );
  AND2_X1 U590 ( .A1(n497), .A2(KEYINPUT44), .ZN(n498) );
  NAND2_X1 U591 ( .A1(n498), .A2(n608), .ZN(n499) );
  NAND2_X1 U592 ( .A1(n500), .A2(n499), .ZN(n524) );
  INV_X1 U593 ( .A(n501), .ZN(n503) );
  INV_X1 U594 ( .A(KEYINPUT64), .ZN(n502) );
  NAND2_X1 U595 ( .A1(n503), .A2(n502), .ZN(n522) );
  INV_X1 U596 ( .A(n504), .ZN(n507) );
  INV_X1 U597 ( .A(n505), .ZN(n556) );
  NAND2_X1 U598 ( .A1(n656), .A2(n556), .ZN(n506) );
  NOR2_X1 U599 ( .A1(n507), .A2(n506), .ZN(n508) );
  XOR2_X1 U600 ( .A(KEYINPUT95), .B(n508), .Z(n509) );
  NAND2_X1 U601 ( .A1(n509), .A2(n660), .ZN(n630) );
  NOR2_X1 U602 ( .A1(n510), .A2(n660), .ZN(n663) );
  AND2_X1 U603 ( .A1(n511), .A2(n663), .ZN(n512) );
  XNOR2_X1 U604 ( .A(n512), .B(KEYINPUT31), .ZN(n644) );
  NAND2_X1 U605 ( .A1(n630), .A2(n644), .ZN(n516) );
  NAND2_X1 U606 ( .A1(n513), .A2(n514), .ZN(n642) );
  NAND2_X1 U607 ( .A1(n642), .A2(n645), .ZN(n676) );
  XOR2_X1 U608 ( .A(n676), .B(KEYINPUT82), .Z(n561) );
  INV_X1 U609 ( .A(n561), .ZN(n515) );
  NAND2_X1 U610 ( .A1(n516), .A2(n515), .ZN(n520) );
  AND2_X1 U611 ( .A1(n652), .A2(n517), .ZN(n519) );
  NAND2_X1 U612 ( .A1(n519), .A2(n518), .ZN(n607) );
  AND2_X1 U613 ( .A1(n520), .A2(n607), .ZN(n521) );
  AND2_X1 U614 ( .A1(n522), .A2(n521), .ZN(n523) );
  INV_X1 U615 ( .A(KEYINPUT45), .ZN(n525) );
  INV_X1 U616 ( .A(n710), .ZN(n591) );
  NAND2_X1 U617 ( .A1(n546), .A2(n670), .ZN(n528) );
  XNOR2_X1 U618 ( .A(n528), .B(n527), .ZN(n536) );
  NOR2_X1 U619 ( .A1(G900), .A2(n529), .ZN(n530) );
  NAND2_X1 U620 ( .A1(G953), .A2(n530), .ZN(n531) );
  XOR2_X1 U621 ( .A(KEYINPUT104), .B(n531), .Z(n532) );
  NOR2_X1 U622 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U623 ( .A(n534), .B(KEYINPUT79), .ZN(n535) );
  NAND2_X1 U624 ( .A1(n535), .A2(n651), .ZN(n544) );
  INV_X1 U625 ( .A(n545), .ZN(n537) );
  NOR2_X1 U626 ( .A1(n537), .A2(n548), .ZN(n538) );
  XOR2_X1 U627 ( .A(KEYINPUT38), .B(n552), .Z(n671) );
  NAND2_X1 U628 ( .A1(n553), .A2(n671), .ZN(n540) );
  XNOR2_X1 U629 ( .A(n540), .B(KEYINPUT39), .ZN(n589) );
  AND2_X1 U630 ( .A1(n376), .A2(n589), .ZN(n542) );
  XNOR2_X1 U631 ( .A(KEYINPUT109), .B(KEYINPUT40), .ZN(n541) );
  XNOR2_X1 U632 ( .A(n542), .B(n541), .ZN(n740) );
  NAND2_X1 U633 ( .A1(n671), .A2(n670), .ZN(n677) );
  XNOR2_X1 U634 ( .A(n543), .B(KEYINPUT41), .ZN(n696) );
  INV_X1 U635 ( .A(n696), .ZN(n668) );
  NAND2_X1 U636 ( .A1(n668), .A2(n549), .ZN(n550) );
  XNOR2_X1 U637 ( .A(n550), .B(KEYINPUT42), .ZN(n741) );
  NAND2_X1 U638 ( .A1(n740), .A2(n741), .ZN(n551) );
  XNOR2_X1 U639 ( .A(n551), .B(KEYINPUT46), .ZN(n579) );
  BUF_X1 U640 ( .A(n552), .Z(n581) );
  NAND2_X1 U641 ( .A1(n553), .A2(n581), .ZN(n554) );
  NOR2_X1 U642 ( .A1(n555), .A2(n554), .ZN(n639) );
  NAND2_X1 U643 ( .A1(n557), .A2(n556), .ZN(n559) );
  OR2_X1 U644 ( .A1(n559), .A2(n558), .ZN(n560) );
  INV_X1 U645 ( .A(n640), .ZN(n564) );
  NOR2_X1 U646 ( .A1(KEYINPUT47), .A2(n561), .ZN(n562) );
  XNOR2_X1 U647 ( .A(n562), .B(KEYINPUT71), .ZN(n563) );
  NOR2_X1 U648 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U649 ( .A1(n639), .A2(n565), .ZN(n574) );
  NAND2_X1 U650 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U651 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U652 ( .A(n571), .B(KEYINPUT36), .ZN(n573) );
  NAND2_X1 U653 ( .A1(n573), .A2(n572), .ZN(n649) );
  AND2_X1 U654 ( .A1(n574), .A2(n649), .ZN(n577) );
  NAND2_X1 U655 ( .A1(n676), .A2(n640), .ZN(n575) );
  NAND2_X1 U656 ( .A1(n575), .A2(KEYINPUT47), .ZN(n576) );
  NAND2_X1 U657 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U658 ( .A(n580), .B(n366), .ZN(n588) );
  INV_X1 U659 ( .A(n581), .ZN(n586) );
  NOR2_X1 U660 ( .A1(n582), .A2(n655), .ZN(n584) );
  XOR2_X1 U661 ( .A(KEYINPUT43), .B(KEYINPUT106), .Z(n583) );
  XNOR2_X1 U662 ( .A(n584), .B(n583), .ZN(n585) );
  NAND2_X1 U663 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U664 ( .A(KEYINPUT107), .B(n587), .ZN(n738) );
  INV_X1 U665 ( .A(n645), .ZN(n636) );
  NAND2_X1 U666 ( .A1(n589), .A2(n636), .ZN(n650) );
  NOR2_X1 U667 ( .A1(n732), .A2(n592), .ZN(n590) );
  NAND2_X1 U668 ( .A1(n591), .A2(n590), .ZN(n595) );
  XNOR2_X1 U669 ( .A(n592), .B(KEYINPUT85), .ZN(n593) );
  NAND2_X1 U670 ( .A1(n593), .A2(KEYINPUT2), .ZN(n594) );
  NAND2_X1 U671 ( .A1(n595), .A2(n594), .ZN(n600) );
  NAND2_X1 U672 ( .A1(KEYINPUT2), .A2(n650), .ZN(n596) );
  XOR2_X1 U673 ( .A(KEYINPUT80), .B(n596), .Z(n597) );
  NAND2_X1 U674 ( .A1(n621), .A2(G472), .ZN(n602) );
  XNOR2_X1 U675 ( .A(n602), .B(n365), .ZN(n605) );
  INV_X1 U676 ( .A(G952), .ZN(n603) );
  AND2_X1 U677 ( .A1(n603), .A2(G953), .ZN(n709) );
  NAND2_X1 U678 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U679 ( .A(n606), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U680 ( .A(n607), .B(G101), .ZN(G3) );
  XNOR2_X1 U681 ( .A(n608), .B(G122), .ZN(G24) );
  NAND2_X1 U682 ( .A1(n621), .A2(G210), .ZN(n613) );
  XOR2_X1 U683 ( .A(KEYINPUT81), .B(KEYINPUT54), .Z(n609) );
  XNOR2_X1 U684 ( .A(n609), .B(KEYINPUT55), .ZN(n610) );
  XNOR2_X1 U685 ( .A(n611), .B(n610), .ZN(n612) );
  XNOR2_X1 U686 ( .A(n613), .B(n612), .ZN(n614) );
  NOR2_X2 U687 ( .A1(n614), .A2(n709), .ZN(n615) );
  XNOR2_X1 U688 ( .A(n615), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U689 ( .A1(n705), .A2(G217), .ZN(n619) );
  XOR2_X1 U690 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n616) );
  XNOR2_X1 U691 ( .A(n617), .B(n616), .ZN(n618) );
  XNOR2_X1 U692 ( .A(n619), .B(n618), .ZN(n620) );
  NOR2_X1 U693 ( .A1(n620), .A2(n709), .ZN(G66) );
  NAND2_X1 U694 ( .A1(n621), .A2(G475), .ZN(n626) );
  XNOR2_X1 U695 ( .A(KEYINPUT65), .B(KEYINPUT120), .ZN(n622) );
  XNOR2_X1 U696 ( .A(n622), .B(KEYINPUT59), .ZN(n623) );
  XNOR2_X1 U697 ( .A(n624), .B(n623), .ZN(n625) );
  XNOR2_X1 U698 ( .A(n626), .B(n625), .ZN(n627) );
  NOR2_X2 U699 ( .A1(n627), .A2(n709), .ZN(n628) );
  XNOR2_X1 U700 ( .A(n628), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X1 U701 ( .A1(n642), .A2(n630), .ZN(n629) );
  XOR2_X1 U702 ( .A(G104), .B(n629), .Z(G6) );
  NOR2_X1 U703 ( .A1(n630), .A2(n645), .ZN(n634) );
  XOR2_X1 U704 ( .A(KEYINPUT111), .B(KEYINPUT26), .Z(n632) );
  XNOR2_X1 U705 ( .A(G107), .B(KEYINPUT27), .ZN(n631) );
  XNOR2_X1 U706 ( .A(n632), .B(n631), .ZN(n633) );
  XNOR2_X1 U707 ( .A(n634), .B(n633), .ZN(G9) );
  XNOR2_X1 U708 ( .A(G110), .B(n635), .ZN(G12) );
  XOR2_X1 U709 ( .A(G128), .B(KEYINPUT29), .Z(n638) );
  NAND2_X1 U710 ( .A1(n636), .A2(n640), .ZN(n637) );
  XNOR2_X1 U711 ( .A(n638), .B(n637), .ZN(G30) );
  XOR2_X1 U712 ( .A(G143), .B(n639), .Z(G45) );
  NAND2_X1 U713 ( .A1(n640), .A2(n376), .ZN(n641) );
  XNOR2_X1 U714 ( .A(n641), .B(G146), .ZN(G48) );
  NOR2_X1 U715 ( .A1(n642), .A2(n644), .ZN(n643) );
  XOR2_X1 U716 ( .A(G113), .B(n643), .Z(G15) );
  NOR2_X1 U717 ( .A1(n645), .A2(n644), .ZN(n646) );
  XOR2_X1 U718 ( .A(KEYINPUT112), .B(n646), .Z(n647) );
  XNOR2_X1 U719 ( .A(G116), .B(n647), .ZN(G18) );
  XOR2_X1 U720 ( .A(G125), .B(KEYINPUT37), .Z(n648) );
  XNOR2_X1 U721 ( .A(n649), .B(n648), .ZN(G27) );
  XNOR2_X1 U722 ( .A(G134), .B(n650), .ZN(G36) );
  NOR2_X1 U723 ( .A1(n652), .A2(n651), .ZN(n654) );
  XNOR2_X1 U724 ( .A(KEYINPUT49), .B(KEYINPUT113), .ZN(n653) );
  XNOR2_X1 U725 ( .A(n654), .B(n653), .ZN(n659) );
  NOR2_X1 U726 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U727 ( .A(n657), .B(KEYINPUT50), .ZN(n658) );
  NOR2_X1 U728 ( .A1(n659), .A2(n658), .ZN(n661) );
  NAND2_X1 U729 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U730 ( .A(n662), .B(KEYINPUT114), .ZN(n665) );
  INV_X1 U731 ( .A(n663), .ZN(n664) );
  NAND2_X1 U732 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U733 ( .A(KEYINPUT51), .B(n666), .Z(n667) );
  NAND2_X1 U734 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U735 ( .A(n669), .B(KEYINPUT115), .ZN(n684) );
  NOR2_X1 U736 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U737 ( .A(n672), .B(KEYINPUT116), .ZN(n673) );
  NOR2_X1 U738 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U739 ( .A(KEYINPUT117), .B(n675), .Z(n680) );
  INV_X1 U740 ( .A(n676), .ZN(n678) );
  NOR2_X1 U741 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U742 ( .A1(n680), .A2(n679), .ZN(n682) );
  INV_X1 U743 ( .A(n681), .ZN(n695) );
  NOR2_X1 U744 ( .A1(n682), .A2(n695), .ZN(n683) );
  NOR2_X1 U745 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U746 ( .A(n685), .B(KEYINPUT52), .ZN(n686) );
  INV_X1 U747 ( .A(KEYINPUT2), .ZN(n688) );
  NAND2_X1 U748 ( .A1(n710), .A2(n688), .ZN(n691) );
  NAND2_X1 U749 ( .A1(n732), .A2(n688), .ZN(n689) );
  XNOR2_X1 U750 ( .A(n689), .B(KEYINPUT84), .ZN(n690) );
  NAND2_X1 U751 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U752 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U753 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U754 ( .A(KEYINPUT118), .B(n697), .Z(n698) );
  NAND2_X1 U755 ( .A1(n705), .A2(G469), .ZN(n703) );
  XOR2_X1 U756 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n699) );
  XOR2_X1 U757 ( .A(n699), .B(KEYINPUT119), .Z(n700) );
  XNOR2_X1 U758 ( .A(n701), .B(n700), .ZN(n702) );
  XNOR2_X1 U759 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U760 ( .A1(n709), .A2(n704), .ZN(G54) );
  NAND2_X1 U761 ( .A1(n705), .A2(G478), .ZN(n707) );
  XNOR2_X1 U762 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U763 ( .A1(n709), .A2(n708), .ZN(G63) );
  NAND2_X1 U764 ( .A1(n591), .A2(n734), .ZN(n715) );
  XOR2_X1 U765 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n712) );
  NAND2_X1 U766 ( .A1(G224), .A2(G953), .ZN(n711) );
  XNOR2_X1 U767 ( .A(n712), .B(n711), .ZN(n713) );
  NAND2_X1 U768 ( .A1(n713), .A2(G898), .ZN(n714) );
  NAND2_X1 U769 ( .A1(n715), .A2(n714), .ZN(n724) );
  XNOR2_X1 U770 ( .A(G101), .B(KEYINPUT124), .ZN(n720) );
  XNOR2_X1 U771 ( .A(n716), .B(n717), .ZN(n718) );
  XNOR2_X1 U772 ( .A(n718), .B(KEYINPUT125), .ZN(n719) );
  XNOR2_X1 U773 ( .A(n720), .B(n719), .ZN(n721) );
  NAND2_X1 U774 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U775 ( .A(n724), .B(n723), .Z(G69) );
  XOR2_X1 U776 ( .A(n726), .B(n725), .Z(n727) );
  XNOR2_X1 U777 ( .A(n728), .B(n727), .ZN(n733) );
  XNOR2_X1 U778 ( .A(G227), .B(n733), .ZN(n729) );
  NAND2_X1 U779 ( .A1(n729), .A2(G900), .ZN(n730) );
  NAND2_X1 U780 ( .A1(n730), .A2(G953), .ZN(n731) );
  XNOR2_X1 U781 ( .A(n731), .B(KEYINPUT126), .ZN(n737) );
  XNOR2_X1 U782 ( .A(n733), .B(n732), .ZN(n735) );
  NAND2_X1 U783 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U784 ( .A1(n737), .A2(n736), .ZN(G72) );
  XOR2_X1 U785 ( .A(G140), .B(n738), .Z(G42) );
  XNOR2_X1 U786 ( .A(G119), .B(n739), .ZN(G21) );
  XNOR2_X1 U787 ( .A(n740), .B(G131), .ZN(G33) );
  XOR2_X1 U788 ( .A(G137), .B(n741), .Z(n742) );
  XNOR2_X1 U789 ( .A(KEYINPUT127), .B(n742), .ZN(G39) );
endmodule

