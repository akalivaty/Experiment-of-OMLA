//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 0 0 1 0 0 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n556, new_n557, new_n558,
    new_n559, new_n562, new_n563, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n614, new_n617, new_n618,
    new_n619, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1142;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT64), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT65), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  AND2_X1   g032(.A1(new_n456), .A2(new_n457), .ZN(G319));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n461), .A2(G125), .ZN(new_n462));
  AND2_X1   g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  XNOR2_X1  g041(.A(new_n466), .B(KEYINPUT66), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n459), .A2(new_n460), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G137), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n464), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n470), .A2(G136), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n469), .A2(new_n465), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  OR2_X1    g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n477), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n474), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G162));
  INV_X1    g055(.A(KEYINPUT4), .ZN(new_n481));
  OAI211_X1 g056(.A(G138), .B(new_n465), .C1(new_n459), .C2(new_n460), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT67), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n484), .B1(new_n483), .B2(new_n482), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n482), .A2(new_n483), .A3(new_n481), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(new_n488), .B2(G2105), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n489), .B1(new_n475), .B2(G126), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n485), .A2(new_n486), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AND2_X1   g068(.A1(new_n490), .A2(new_n486), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n494), .A2(KEYINPUT68), .A3(new_n485), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  INV_X1    g072(.A(KEYINPUT6), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G651), .ZN(new_n499));
  XNOR2_X1  g074(.A(new_n499), .B(KEYINPUT69), .ZN(new_n500));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT6), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n504), .B1(new_n506), .B2(KEYINPUT70), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT5), .A3(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n503), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(G50), .A2(new_n505), .B1(new_n512), .B2(G88), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n510), .A2(G62), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n514), .A2(new_n515), .B1(G75), .B2(G543), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n516), .B1(new_n515), .B2(new_n514), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n513), .A2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND2_X1  g095(.A1(new_n512), .A2(G89), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n505), .A2(G51), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  AND3_X1   g099(.A1(new_n507), .A2(KEYINPUT72), .A3(new_n509), .ZN(new_n525));
  AOI21_X1  g100(.A(KEYINPUT72), .B1(new_n507), .B2(new_n509), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n527), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n521), .A2(new_n522), .A3(new_n524), .A4(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  NAND4_X1  g105(.A1(new_n500), .A2(G52), .A3(G543), .A4(new_n502), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n500), .A2(G90), .A3(new_n510), .A4(new_n502), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT72), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n508), .A2(KEYINPUT5), .A3(G543), .ZN(new_n535));
  AOI21_X1  g110(.A(G543), .B1(new_n508), .B2(KEYINPUT5), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n507), .A2(KEYINPUT72), .A3(new_n509), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n537), .A2(G64), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n501), .B1(new_n541), .B2(KEYINPUT73), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT73), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n539), .A2(new_n543), .A3(new_n540), .ZN(new_n544));
  AOI211_X1 g119(.A(KEYINPUT74), .B(new_n533), .C1(new_n542), .C2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT74), .ZN(new_n546));
  INV_X1    g121(.A(G64), .ZN(new_n547));
  NOR3_X1   g122(.A1(new_n525), .A2(new_n526), .A3(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n540), .ZN(new_n549));
  OAI21_X1  g124(.A(KEYINPUT73), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n550), .A2(G651), .A3(new_n544), .ZN(new_n551));
  INV_X1    g126(.A(new_n533), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n546), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n545), .A2(new_n553), .ZN(G301));
  INV_X1    g129(.A(G301), .ZN(G171));
  AOI22_X1  g130(.A1(G43), .A2(new_n505), .B1(new_n512), .B2(G81), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n527), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n501), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(G860), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n558), .A2(new_n559), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  AND2_X1   g139(.A1(new_n500), .A2(new_n502), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G543), .ZN(new_n566));
  INV_X1    g141(.A(G53), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT9), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n505), .A2(new_n569), .A3(G53), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n572));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n511), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n512), .A2(G91), .B1(G651), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n571), .A2(new_n572), .A3(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n572), .B1(new_n571), .B2(new_n576), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(G299));
  NAND4_X1  g155(.A1(new_n500), .A2(G87), .A3(new_n510), .A4(new_n502), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT76), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n500), .A2(G49), .A3(G543), .A4(new_n502), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT77), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n583), .B(new_n584), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n527), .B2(G74), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n582), .A2(new_n585), .A3(new_n586), .ZN(G288));
  NAND2_X1  g162(.A1(new_n505), .A2(G48), .ZN(new_n588));
  AND2_X1   g163(.A1(new_n510), .A2(G61), .ZN(new_n589));
  AND2_X1   g164(.A1(G73), .A2(G543), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AND2_X1   g166(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n512), .A2(G86), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(G305));
  AOI22_X1  g169(.A1(G47), .A2(new_n505), .B1(new_n512), .B2(G85), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n527), .A2(G60), .ZN(new_n597));
  NAND2_X1  g172(.A1(G72), .A2(G543), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n501), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G290));
  NAND2_X1  g176(.A1(new_n512), .A2(G92), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n512), .A2(KEYINPUT10), .A3(G92), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n505), .A2(G54), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n510), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n606), .B(new_n607), .C1(new_n501), .C2(new_n608), .ZN(new_n609));
  MUX2_X1   g184(.A(new_n609), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g185(.A(new_n609), .B(G301), .S(G868), .Z(G321));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NOR2_X1   g187(.A1(G286), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g188(.A(G299), .B(KEYINPUT78), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(new_n612), .ZN(G297));
  AOI21_X1  g190(.A(new_n613), .B1(new_n614), .B2(new_n612), .ZN(G280));
  OAI21_X1  g191(.A(new_n607), .B1(new_n501), .B2(new_n608), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n617), .B1(new_n604), .B2(new_n605), .ZN(new_n618));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(G860), .ZN(G148));
  NAND2_X1  g195(.A1(new_n558), .A2(new_n612), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n609), .A2(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(new_n612), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n467), .A2(new_n461), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT12), .Z(new_n626));
  XOR2_X1   g201(.A(KEYINPUT79), .B(KEYINPUT13), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(G2100), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n470), .A2(G135), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n475), .A2(G123), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  INV_X1    g209(.A(G111), .ZN(new_n635));
  AOI22_X1  g210(.A1(new_n634), .A2(KEYINPUT80), .B1(new_n635), .B2(G2105), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(KEYINPUT80), .B2(new_n634), .ZN(new_n637));
  AND3_X1   g212(.A1(new_n632), .A2(new_n633), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2096), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n630), .A2(new_n631), .A3(new_n639), .ZN(G156));
  XOR2_X1   g215(.A(KEYINPUT15), .B(G2435), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2438), .ZN(new_n642));
  XOR2_X1   g217(.A(G2427), .B(G2430), .Z(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT82), .B(KEYINPUT14), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n642), .A2(new_n643), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2443), .B(G2446), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2451), .B(G2454), .Z(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n649), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT83), .Z(new_n656));
  OAI211_X1 g231(.A(new_n656), .B(G14), .C1(new_n654), .C2(new_n653), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(G401));
  XOR2_X1   g233(.A(G2072), .B(G2078), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT17), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n662), .B2(new_n659), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n663), .B1(KEYINPUT84), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n666), .B1(KEYINPUT84), .B2(new_n665), .ZN(new_n667));
  INV_X1    g242(.A(new_n659), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n668), .A2(new_n664), .A3(new_n661), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT18), .Z(new_n670));
  NAND3_X1  g245(.A1(new_n660), .A2(new_n664), .A3(new_n662), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2096), .B(G2100), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G227));
  XOR2_X1   g249(.A(G1971), .B(G1976), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n677), .A2(new_n678), .ZN(new_n681));
  NOR3_X1   g256(.A1(new_n676), .A2(new_n681), .A3(new_n679), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n676), .A2(new_n681), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n684));
  AOI211_X1 g259(.A(new_n680), .B(new_n682), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(new_n683), .B2(new_n684), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G1981), .B(G1986), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(G229));
  MUX2_X1   g267(.A(G6), .B(G305), .S(G16), .Z(new_n693));
  XOR2_X1   g268(.A(KEYINPUT32), .B(G1981), .Z(new_n694));
  XOR2_X1   g269(.A(new_n693), .B(new_n694), .Z(new_n695));
  INV_X1    g270(.A(G16), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n696), .A2(G23), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(G288), .B2(G16), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT33), .B(G1976), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n696), .A2(G22), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT86), .Z(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G166), .B2(new_n696), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n703), .A2(G1971), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(G1971), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(new_n698), .B2(new_n699), .ZN(new_n706));
  NOR4_X1   g281(.A1(new_n695), .A2(new_n700), .A3(new_n704), .A4(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT34), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n600), .A2(new_n696), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(new_n696), .B2(G24), .ZN(new_n712));
  INV_X1    g287(.A(G1986), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(G29), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G25), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n470), .A2(G131), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n475), .A2(G119), .ZN(new_n718));
  OR2_X1    g293(.A1(G95), .A2(G2105), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n719), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n716), .B1(new_n722), .B2(new_n715), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT35), .B(G1991), .Z(new_n724));
  XOR2_X1   g299(.A(new_n723), .B(new_n724), .Z(new_n725));
  INV_X1    g300(.A(new_n712), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(G1986), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n709), .A2(new_n710), .A3(new_n714), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT36), .ZN(new_n729));
  AOI22_X1  g304(.A1(G105), .A2(new_n467), .B1(new_n470), .B2(G141), .ZN(new_n730));
  NAND3_X1  g305(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT26), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G129), .B2(new_n475), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n735), .A2(new_n715), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n715), .B2(G32), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT27), .B(G1996), .Z(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT87), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n737), .A2(new_n739), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT25), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n461), .A2(G127), .ZN(new_n744));
  NAND2_X1  g319(.A1(G115), .A2(G2104), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n465), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  AOI211_X1 g321(.A(new_n743), .B(new_n746), .C1(G139), .C2(new_n470), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G29), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G29), .B2(G33), .ZN(new_n749));
  INV_X1    g324(.A(G2072), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n741), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G1966), .ZN(new_n752));
  NOR2_X1   g327(.A1(G168), .A2(new_n696), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n696), .B2(G21), .ZN(new_n754));
  AOI211_X1 g329(.A(new_n740), .B(new_n751), .C1(new_n752), .C2(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G34), .ZN(new_n756));
  AOI21_X1  g331(.A(G29), .B1(new_n756), .B2(KEYINPUT24), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(KEYINPUT24), .B2(new_n756), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n472), .B2(new_n715), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G2084), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n749), .A2(new_n750), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n715), .A2(G26), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT28), .Z(new_n763));
  NAND2_X1  g338(.A1(new_n470), .A2(G140), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n475), .A2(G128), .ZN(new_n765));
  OR2_X1    g340(.A1(G104), .A2(G2105), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n766), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n764), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n763), .B1(new_n768), .B2(G29), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G2067), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT89), .B(KEYINPUT31), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G11), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT30), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G28), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n715), .B1(new_n773), .B2(G28), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(KEYINPUT90), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(KEYINPUT90), .B2(new_n775), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n772), .B(new_n777), .C1(new_n638), .C2(G29), .ZN(new_n778));
  AND4_X1   g353(.A1(new_n760), .A2(new_n761), .A3(new_n770), .A4(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(G4), .A2(G16), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n618), .B2(G16), .ZN(new_n781));
  INV_X1    g356(.A(G1348), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n755), .A2(new_n779), .A3(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n754), .A2(new_n752), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT88), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n715), .A2(G35), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT91), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G162), .B2(new_n715), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT29), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(G2090), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n715), .A2(G27), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G164), .B2(new_n715), .ZN(new_n793));
  INV_X1    g368(.A(G2078), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  MUX2_X1   g370(.A(G19), .B(new_n558), .S(G16), .Z(new_n796));
  OR2_X1    g371(.A1(new_n796), .A2(G1341), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(G1341), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n791), .A2(new_n795), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  NOR3_X1   g374(.A1(new_n784), .A2(new_n786), .A3(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(G5), .A2(G16), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G171), .B2(G16), .ZN(new_n802));
  INV_X1    g377(.A(G1961), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n696), .A2(G20), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT92), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT23), .ZN(new_n807));
  INV_X1    g382(.A(G299), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(new_n696), .ZN(new_n809));
  INV_X1    g384(.A(G1956), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n800), .A2(new_n804), .A3(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT93), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n729), .A2(new_n813), .ZN(G150));
  INV_X1    g389(.A(G150), .ZN(G311));
  NAND3_X1  g390(.A1(new_n565), .A2(G93), .A3(new_n510), .ZN(new_n816));
  INV_X1    g391(.A(G55), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n566), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n527), .A2(G67), .ZN(new_n819));
  NAND2_X1  g394(.A1(G80), .A2(G543), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n501), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n822), .A2(new_n559), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT95), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT37), .Z(new_n825));
  NAND2_X1  g400(.A1(new_n618), .A2(G559), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT38), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n558), .B(new_n822), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n827), .B(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(KEYINPUT39), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT94), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n559), .B1(new_n831), .B2(KEYINPUT39), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n825), .B1(new_n833), .B2(new_n834), .ZN(G145));
  NAND2_X1  g410(.A1(new_n470), .A2(G142), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT96), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n475), .A2(G130), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n465), .A2(G118), .ZN(new_n839));
  OAI21_X1  g414(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n837), .B(new_n838), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT98), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(new_n722), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n747), .B(new_n735), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n626), .B(KEYINPUT97), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n491), .B(new_n768), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n845), .B(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n472), .B(G162), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n638), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(G37), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n849), .A2(new_n851), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XOR2_X1   g431(.A(KEYINPUT99), .B(KEYINPUT40), .Z(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(G395));
  OAI21_X1  g433(.A(new_n609), .B1(new_n578), .B2(new_n579), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(KEYINPUT100), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n571), .A2(new_n576), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT75), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n862), .A2(new_n577), .A3(new_n618), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT100), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n864), .B(new_n609), .C1(new_n578), .C2(new_n579), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n860), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT41), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n859), .A2(new_n863), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n870), .A2(KEYINPUT101), .A3(KEYINPUT41), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT101), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n872), .B1(new_n869), .B2(new_n867), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n868), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n828), .B(new_n622), .Z(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(new_n870), .B2(new_n875), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n600), .B(G303), .ZN(new_n878));
  XNOR2_X1  g453(.A(G305), .B(G288), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT42), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n877), .A2(new_n881), .ZN(new_n883));
  OAI21_X1  g458(.A(G868), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n884), .B1(G868), .B2(new_n822), .ZN(G295));
  OAI21_X1  g460(.A(new_n884), .B1(G868), .B2(new_n822), .ZN(G331));
  OAI21_X1  g461(.A(KEYINPUT102), .B1(new_n545), .B2(new_n553), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n539), .A2(new_n543), .A3(new_n540), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n543), .B1(new_n539), .B2(new_n540), .ZN(new_n889));
  NOR3_X1   g464(.A1(new_n888), .A2(new_n889), .A3(new_n501), .ZN(new_n890));
  OAI21_X1  g465(.A(KEYINPUT74), .B1(new_n890), .B2(new_n533), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT102), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n551), .A2(new_n546), .A3(new_n552), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n887), .A2(new_n894), .A3(G286), .ZN(new_n895));
  OAI211_X1 g470(.A(KEYINPUT102), .B(G168), .C1(new_n545), .C2(new_n553), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(new_n829), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n895), .A2(new_n828), .A3(new_n896), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n874), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n902));
  AOI21_X1  g477(.A(KEYINPUT103), .B1(new_n897), .B2(new_n829), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n904));
  AOI211_X1 g479(.A(new_n904), .B(new_n828), .C1(new_n895), .C2(new_n896), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n899), .A2(new_n869), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n902), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n898), .A2(new_n904), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n897), .A2(KEYINPUT103), .A3(new_n829), .ZN(new_n910));
  AND4_X1   g485(.A1(new_n902), .A2(new_n909), .A3(new_n907), .A4(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n901), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(G37), .B1(new_n912), .B2(new_n880), .ZN(new_n913));
  INV_X1    g488(.A(new_n880), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n914), .B(new_n901), .C1(new_n908), .C2(new_n911), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT43), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n907), .A2(new_n898), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n909), .A2(new_n899), .A3(new_n910), .ZN(new_n918));
  NOR3_X1   g493(.A1(new_n578), .A2(new_n609), .A3(new_n579), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n618), .B1(new_n862), .B2(new_n577), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n867), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT105), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n860), .A2(KEYINPUT41), .A3(new_n863), .A4(new_n865), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n869), .A2(new_n924), .A3(new_n867), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n922), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n917), .B1(new_n918), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(G37), .B1(new_n927), .B2(new_n880), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n928), .A2(KEYINPUT43), .A3(new_n915), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT44), .B1(new_n916), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n932), .B1(new_n913), .B2(new_n915), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n928), .A2(new_n932), .A3(new_n915), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n930), .A2(new_n935), .ZN(G397));
  XNOR2_X1  g511(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n937));
  NAND2_X1  g512(.A1(G160), .A2(G40), .ZN(new_n938));
  AOI21_X1  g513(.A(G1384), .B1(new_n494), .B2(new_n485), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(G1384), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n491), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT107), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n938), .B1(new_n945), .B2(KEYINPUT50), .ZN(new_n946));
  AOI21_X1  g521(.A(G1384), .B1(new_n493), .B2(new_n495), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT50), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n947), .A2(KEYINPUT115), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT115), .B1(new_n947), .B2(new_n948), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n946), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G40), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n472), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n953), .B1(new_n943), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n496), .A2(new_n942), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n955), .B1(new_n956), .B2(new_n954), .ZN(new_n957));
  XNOR2_X1  g532(.A(KEYINPUT56), .B(G2072), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n951), .A2(new_n810), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT116), .ZN(new_n960));
  OR2_X1    g535(.A1(new_n960), .A2(KEYINPUT57), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(KEYINPUT57), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n571), .A2(new_n576), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n861), .A2(new_n960), .A3(KEYINPUT57), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n959), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n963), .ZN(new_n966));
  INV_X1    g541(.A(new_n955), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n967), .B(new_n958), .C1(KEYINPUT45), .C2(new_n947), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  AOI211_X1 g544(.A(new_n966), .B(new_n969), .C1(new_n951), .C2(new_n810), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n937), .B1(new_n965), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n972), .B1(new_n945), .B2(KEYINPUT50), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n938), .B1(new_n956), .B2(KEYINPUT50), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n941), .A2(new_n944), .A3(KEYINPUT108), .A4(new_n948), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G2067), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n941), .A2(new_n944), .A3(new_n953), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n976), .A2(new_n782), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n980), .A2(KEYINPUT60), .A3(new_n609), .ZN(new_n981));
  XNOR2_X1  g556(.A(KEYINPUT119), .B(G1996), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n957), .A2(new_n982), .ZN(new_n983));
  XOR2_X1   g558(.A(KEYINPUT58), .B(G1341), .Z(new_n984));
  NAND2_X1  g559(.A1(new_n978), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n558), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  OR2_X1    g561(.A1(new_n986), .A2(KEYINPUT59), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(KEYINPUT59), .ZN(new_n988));
  AND3_X1   g563(.A1(new_n981), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n970), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT61), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n609), .B1(new_n980), .B2(KEYINPUT60), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(KEYINPUT60), .B2(new_n980), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n971), .A2(new_n989), .A3(new_n991), .A4(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n980), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n995), .A2(KEYINPUT117), .A3(new_n618), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT117), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(new_n980), .B2(new_n609), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT118), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n959), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n966), .B1(new_n959), .B2(new_n999), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n996), .B(new_n998), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n990), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n994), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1981), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n592), .A2(new_n1005), .A3(new_n593), .ZN(new_n1006));
  INV_X1    g581(.A(new_n512), .ZN(new_n1007));
  XOR2_X1   g582(.A(KEYINPUT112), .B(G86), .Z(new_n1008));
  OAI211_X1 g583(.A(new_n588), .B(new_n591), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(G1981), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1006), .B(new_n1010), .C1(KEYINPUT113), .C2(KEYINPUT49), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT49), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1011), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G8), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n979), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1006), .A2(new_n1010), .A3(KEYINPUT113), .A4(KEYINPUT49), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  XOR2_X1   g593(.A(KEYINPUT110), .B(G1976), .Z(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT52), .B1(G288), .B2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n582), .A2(new_n585), .A3(G1976), .A4(new_n586), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1020), .A2(new_n978), .A3(G8), .A4(new_n1021), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1022), .A2(KEYINPUT111), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1022), .A2(KEYINPUT111), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1018), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n978), .A2(G8), .A3(new_n1021), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT52), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT109), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n1027), .B(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1025), .A2(new_n1029), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n957), .A2(G1971), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1031), .B1(new_n976), .B2(G2090), .ZN(new_n1032));
  NAND2_X1  g607(.A1(G303), .A2(G8), .ZN(new_n1033));
  XOR2_X1   g608(.A(new_n1033), .B(KEYINPUT55), .Z(new_n1034));
  NAND3_X1  g609(.A1(new_n1032), .A2(G8), .A3(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1031), .B1(new_n951), .B2(G2090), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1036), .A2(G8), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1030), .B(new_n1035), .C1(new_n1034), .C2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n945), .A2(new_n954), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n947), .A2(KEYINPUT45), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1039), .A2(new_n1040), .A3(new_n953), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n752), .ZN(new_n1042));
  INV_X1    g617(.A(G2084), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n973), .A2(new_n974), .A3(new_n1043), .A4(new_n975), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(G286), .A2(G8), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n1046), .B(KEYINPUT121), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1015), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1048), .B(KEYINPUT51), .C1(new_n1049), .C2(new_n1047), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1049), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1047), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1050), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n957), .A2(new_n794), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n976), .A2(new_n803), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n794), .A2(KEYINPUT53), .ZN(new_n1059));
  OR2_X1    g634(.A1(new_n1041), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(G171), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n939), .A2(KEYINPUT45), .ZN(new_n1063));
  NOR3_X1   g638(.A1(new_n955), .A2(new_n1063), .A3(new_n1059), .ZN(new_n1064));
  XNOR2_X1  g639(.A(new_n1064), .B(KEYINPUT122), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1058), .A2(G301), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT54), .B1(new_n1062), .B2(new_n1066), .ZN(new_n1067));
  NOR3_X1   g642(.A1(new_n1038), .A2(new_n1055), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1058), .A2(new_n1065), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(G171), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1058), .A2(G301), .A3(new_n1060), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(KEYINPUT54), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT123), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT123), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1070), .A2(new_n1074), .A3(KEYINPUT54), .A4(new_n1071), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1004), .A2(new_n1068), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT62), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT124), .B1(new_n1055), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT124), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1050), .A2(new_n1054), .A3(new_n1080), .A4(KEYINPUT62), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT62), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n1083), .A2(new_n1038), .A3(new_n1062), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1032), .A2(G8), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1030), .A2(new_n1034), .A3(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(G288), .A2(G1976), .ZN(new_n1088));
  XOR2_X1   g663(.A(new_n1088), .B(KEYINPUT114), .Z(new_n1089));
  AND2_X1   g664(.A1(new_n1018), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1006), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1016), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1087), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT63), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1049), .A2(G168), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1094), .B1(new_n1038), .B2(new_n1095), .ZN(new_n1096));
  OR2_X1    g671(.A1(new_n1086), .A2(new_n1034), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1095), .A2(new_n1094), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1097), .A2(new_n1030), .A3(new_n1035), .A4(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1093), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1077), .A2(new_n1085), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1063), .A2(new_n953), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1102), .B(KEYINPUT106), .ZN(new_n1103));
  XOR2_X1   g678(.A(new_n721), .B(new_n724), .Z(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n768), .B(new_n977), .ZN(new_n1106));
  INV_X1    g681(.A(G1996), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1106), .B1(new_n1107), .B2(new_n735), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1103), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1102), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1110), .A2(new_n1107), .A3(new_n735), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1105), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n600), .B(new_n713), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1112), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1101), .A2(new_n1114), .ZN(new_n1115));
  NOR3_X1   g690(.A1(G290), .A2(new_n1102), .A3(G1986), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1116), .B(KEYINPUT127), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n1117), .B(KEYINPUT48), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT126), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1112), .A2(new_n1119), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1112), .A2(new_n1119), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n1118), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1110), .A2(new_n1107), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT46), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1125), .B(KEYINPUT125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1106), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1103), .B1(new_n734), .B2(new_n1127), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1126), .B(new_n1128), .C1(new_n1124), .C2(new_n1123), .ZN(new_n1129));
  XOR2_X1   g704(.A(new_n1129), .B(KEYINPUT47), .Z(new_n1130));
  NAND2_X1  g705(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n722), .A2(new_n724), .ZN(new_n1132));
  OAI22_X1  g707(.A1(new_n1131), .A2(new_n1132), .B1(G2067), .B2(new_n768), .ZN(new_n1133));
  AOI211_X1 g708(.A(new_n1122), .B(new_n1130), .C1(new_n1103), .C2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1115), .A2(new_n1134), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g710(.A1(new_n933), .A2(new_n934), .ZN(new_n1137));
  INV_X1    g711(.A(G319), .ZN(new_n1138));
  NOR3_X1   g712(.A1(G229), .A2(new_n1138), .A3(G227), .ZN(new_n1139));
  OAI211_X1 g713(.A(new_n657), .B(new_n1139), .C1(new_n854), .C2(new_n855), .ZN(new_n1140));
  NOR2_X1   g714(.A1(new_n1137), .A2(new_n1140), .ZN(G308));
  AND2_X1   g715(.A1(new_n1139), .A2(new_n657), .ZN(new_n1142));
  OAI221_X1 g716(.A(new_n1142), .B1(new_n855), .B2(new_n854), .C1(new_n933), .C2(new_n934), .ZN(G225));
endmodule


