//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT22), .B(G137), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(G221), .A3(G234), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n191), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G140), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G125), .ZN(new_n197));
  INV_X1    g011(.A(G125), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G140), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n197), .A2(new_n199), .A3(KEYINPUT16), .ZN(new_n200));
  OR3_X1    g014(.A1(new_n198), .A2(KEYINPUT16), .A3(G140), .ZN(new_n201));
  AND3_X1   g015(.A1(new_n200), .A2(G146), .A3(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(G146), .B1(new_n200), .B2(new_n201), .ZN(new_n203));
  INV_X1    g017(.A(G119), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G128), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G119), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT24), .B(G110), .ZN(new_n209));
  OAI22_X1  g023(.A1(new_n202), .A2(new_n203), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT78), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n205), .A2(KEYINPUT23), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT77), .B1(new_n204), .B2(G128), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n212), .B(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G110), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n211), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n212), .A2(KEYINPUT77), .A3(new_n207), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n213), .A2(KEYINPUT23), .A3(new_n205), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(KEYINPUT78), .A3(G110), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n210), .B1(new_n216), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n200), .A2(new_n201), .A3(G146), .ZN(new_n222));
  XNOR2_X1  g036(.A(G125), .B(G140), .ZN(new_n223));
  INV_X1    g037(.A(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n208), .A2(new_n209), .ZN(new_n227));
  XNOR2_X1  g041(.A(new_n227), .B(KEYINPUT79), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n214), .A2(new_n215), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n226), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n195), .B1(new_n221), .B2(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n208), .A2(new_n209), .ZN(new_n232));
  INV_X1    g046(.A(new_n203), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n232), .B1(new_n233), .B2(new_n222), .ZN(new_n234));
  AOI21_X1  g048(.A(KEYINPUT78), .B1(new_n219), .B2(G110), .ZN(new_n235));
  AOI211_X1 g049(.A(new_n211), .B(new_n215), .C1(new_n217), .C2(new_n218), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n234), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n226), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT79), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n227), .B(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n219), .A2(G110), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n238), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n237), .A2(new_n242), .A3(new_n194), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n231), .A2(new_n188), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT25), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n231), .A2(KEYINPUT25), .A3(new_n243), .A4(new_n188), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n190), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n231), .A2(new_n243), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n189), .A2(G902), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(G214), .B1(G237), .B2(G902), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n192), .A2(G952), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n256), .B1(G234), .B2(G237), .ZN(new_n257));
  INV_X1    g071(.A(G234), .ZN(new_n258));
  INV_X1    g072(.A(G237), .ZN(new_n259));
  OAI21_X1  g073(.A(G902), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(new_n192), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT21), .B(G898), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n257), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(G210), .B1(G237), .B2(G902), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT82), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n266), .A2(KEYINPUT3), .ZN(new_n267));
  INV_X1    g081(.A(G104), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n268), .A2(G107), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n266), .A2(KEYINPUT3), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n267), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n268), .A2(G107), .ZN(new_n272));
  INV_X1    g086(.A(G107), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G104), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT3), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(KEYINPUT82), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n272), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(G101), .B1(new_n271), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n273), .A2(G104), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n279), .B1(new_n269), .B2(new_n267), .ZN(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT83), .B(G101), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n275), .A2(KEYINPUT82), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n276), .B1(new_n282), .B2(new_n274), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n280), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n278), .A2(KEYINPUT4), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G116), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n286), .A2(G119), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT68), .B1(new_n204), .B2(G116), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT68), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(new_n286), .A3(G119), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n287), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  XOR2_X1   g105(.A(KEYINPUT2), .B(G113), .Z(new_n292));
  XNOR2_X1  g106(.A(new_n291), .B(new_n292), .ZN(new_n293));
  XNOR2_X1  g107(.A(KEYINPUT84), .B(KEYINPUT4), .ZN(new_n294));
  OAI211_X1 g108(.A(G101), .B(new_n294), .C1(new_n271), .C2(new_n277), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n285), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n291), .A2(new_n292), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n204), .A2(G116), .ZN(new_n298));
  OAI21_X1  g112(.A(G113), .B1(new_n298), .B2(KEYINPUT5), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n299), .B1(new_n291), .B2(KEYINPUT5), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(G101), .B1(new_n279), .B2(new_n269), .ZN(new_n302));
  AND2_X1   g116(.A1(new_n284), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n296), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(G110), .B(G122), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n296), .A2(new_n304), .A3(new_n306), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(KEYINPUT6), .A3(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT65), .B1(new_n224), .B2(G143), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT65), .ZN(new_n312));
  INV_X1    g126(.A(G143), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n313), .A3(G146), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n311), .A2(new_n314), .B1(G143), .B2(new_n224), .ZN(new_n315));
  NAND2_X1  g129(.A1(KEYINPUT0), .A2(G128), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT64), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n316), .B(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(KEYINPUT0), .A2(G128), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n224), .A2(G143), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n313), .A2(G146), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AOI22_X1  g137(.A1(new_n315), .A2(new_n317), .B1(new_n319), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G125), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n311), .A2(new_n314), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n206), .A2(KEYINPUT1), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(new_n321), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n321), .A2(new_n322), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT1), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n331), .B1(G143), .B2(new_n224), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n330), .B1(new_n332), .B2(new_n206), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n329), .A2(new_n198), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n326), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n192), .A2(G224), .ZN(new_n336));
  XOR2_X1   g150(.A(new_n336), .B(KEYINPUT87), .Z(new_n337));
  XNOR2_X1  g151(.A(new_n335), .B(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT6), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n305), .A2(new_n339), .A3(new_n307), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n310), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n306), .B(KEYINPUT8), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n284), .A2(new_n302), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n344), .B1(new_n297), .B2(new_n300), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT88), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n346), .B1(new_n304), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n301), .A2(new_n303), .A3(KEYINPUT88), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n343), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT89), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT7), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n337), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n326), .A2(new_n351), .A3(new_n334), .A4(new_n353), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n353), .B(new_n334), .C1(new_n198), .C2(new_n324), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT89), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n324), .A2(new_n198), .ZN(new_n357));
  INV_X1    g171(.A(new_n334), .ZN(new_n358));
  OAI22_X1  g172(.A1(new_n357), .A2(new_n358), .B1(new_n352), .B2(new_n337), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n309), .A2(new_n354), .A3(new_n356), .A4(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n188), .B1(new_n350), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n265), .B1(new_n341), .B2(new_n361), .ZN(new_n362));
  AND4_X1   g176(.A1(new_n309), .A2(new_n354), .A3(new_n359), .A4(new_n356), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n304), .A2(new_n347), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n364), .A2(new_n349), .A3(new_n345), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n342), .ZN(new_n366));
  AOI21_X1  g180(.A(G902), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n310), .A2(new_n338), .A3(new_n340), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n264), .A3(new_n368), .ZN(new_n369));
  AOI211_X1 g183(.A(new_n255), .B(new_n263), .C1(new_n362), .C2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n329), .A2(new_n333), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n303), .A2(KEYINPUT10), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n285), .A2(new_n324), .A3(new_n295), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT10), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT85), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n329), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n332), .A2(new_n206), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n315), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n327), .A2(KEYINPUT85), .A3(new_n321), .A4(new_n328), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n284), .A2(new_n302), .A3(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n375), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n383), .A2(KEYINPUT86), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT86), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n329), .B(new_n376), .C1(new_n315), .C2(new_n378), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n386), .A2(new_n302), .A3(new_n284), .A4(new_n381), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n385), .B1(new_n387), .B2(new_n375), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n374), .B1(new_n384), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT11), .ZN(new_n390));
  INV_X1    g204(.A(G134), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n390), .B1(new_n391), .B2(G137), .ZN(new_n392));
  INV_X1    g206(.A(G137), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(KEYINPUT11), .A3(G134), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n393), .A2(G134), .ZN(new_n396));
  OAI21_X1  g210(.A(G131), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT67), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n393), .A2(KEYINPUT11), .A3(G134), .ZN(new_n399));
  AOI21_X1  g213(.A(KEYINPUT11), .B1(new_n393), .B2(G134), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AND2_X1   g215(.A1(KEYINPUT66), .A2(G131), .ZN(new_n402));
  NOR2_X1   g216(.A1(KEYINPUT66), .A2(G131), .ZN(new_n403));
  NOR3_X1   g217(.A1(new_n396), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n398), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  OR2_X1    g219(.A1(KEYINPUT66), .A2(G131), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n391), .A2(G137), .ZN(new_n407));
  NAND2_X1  g221(.A1(KEYINPUT66), .A2(G131), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n395), .A2(new_n409), .A3(KEYINPUT67), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n397), .B1(new_n405), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n389), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n192), .A2(G227), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n413), .B(KEYINPUT81), .ZN(new_n414));
  XNOR2_X1  g228(.A(G110), .B(G140), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n414), .B(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n372), .A2(new_n373), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n383), .A2(KEYINPUT86), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n387), .A2(new_n385), .A3(new_n375), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G131), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n421), .B1(new_n401), .B2(new_n407), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n401), .A2(new_n404), .A3(new_n398), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT67), .B1(new_n395), .B2(new_n409), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n416), .B1(new_n420), .B2(new_n425), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n374), .B(new_n425), .C1(new_n384), .C2(new_n388), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT12), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n284), .A2(new_n302), .A3(new_n381), .ZN(new_n429));
  INV_X1    g243(.A(new_n371), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n429), .A2(new_n386), .B1(new_n430), .B2(new_n344), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n428), .B1(new_n431), .B2(new_n425), .ZN(new_n432));
  OAI22_X1  g246(.A1(new_n380), .A2(new_n382), .B1(new_n303), .B2(new_n371), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(KEYINPUT12), .A3(new_n411), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n427), .A2(new_n435), .ZN(new_n436));
  AOI22_X1  g250(.A1(new_n412), .A2(new_n426), .B1(new_n436), .B2(new_n416), .ZN(new_n437));
  OAI21_X1  g251(.A(G469), .B1(new_n437), .B2(G902), .ZN(new_n438));
  INV_X1    g252(.A(G469), .ZN(new_n439));
  INV_X1    g253(.A(new_n416), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n440), .B1(new_n412), .B2(new_n427), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n427), .A2(new_n440), .A3(new_n435), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n439), .B(new_n188), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT9), .B(G234), .ZN(new_n445));
  OAI21_X1  g259(.A(G221), .B1(new_n445), .B2(G902), .ZN(new_n446));
  XOR2_X1   g260(.A(new_n446), .B(KEYINPUT80), .Z(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(G113), .B(G122), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(new_n268), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT90), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n197), .A2(new_n199), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT19), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n223), .A2(KEYINPUT19), .ZN(new_n455));
  AOI21_X1  g269(.A(G146), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n451), .B1(new_n456), .B2(new_n202), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n452), .A2(new_n453), .ZN(new_n458));
  AOI21_X1  g272(.A(KEYINPUT19), .B1(new_n197), .B2(new_n199), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n224), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(KEYINPUT90), .A3(new_n222), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n406), .A2(new_n408), .ZN(new_n462));
  NOR2_X1   g276(.A1(G237), .A2(G953), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n463), .A2(G143), .A3(G214), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(G143), .B1(new_n463), .B2(G214), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n259), .A2(new_n192), .A3(G214), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n313), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n469), .A2(new_n406), .A3(new_n408), .A4(new_n464), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n457), .A2(new_n461), .A3(new_n471), .ZN(new_n472));
  OAI211_X1 g286(.A(KEYINPUT18), .B(G131), .C1(new_n465), .C2(new_n466), .ZN(new_n473));
  NAND2_X1  g287(.A1(KEYINPUT18), .A2(G131), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n469), .A2(new_n464), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n452), .A2(G146), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n225), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n473), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n450), .B1(new_n472), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n478), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT17), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n467), .A2(new_n481), .A3(new_n470), .ZN(new_n482));
  OAI211_X1 g296(.A(KEYINPUT17), .B(new_n462), .C1(new_n465), .C2(new_n466), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n233), .A2(new_n483), .A3(new_n222), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n482), .B1(KEYINPUT91), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT91), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n233), .A2(new_n483), .A3(new_n486), .A4(new_n222), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n480), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n479), .B1(new_n488), .B2(new_n450), .ZN(new_n489));
  NOR2_X1   g303(.A1(G475), .A2(G902), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(KEYINPUT20), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT20), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n484), .A2(KEYINPUT91), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n494), .B(new_n487), .C1(KEYINPUT17), .C2(new_n471), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n495), .A2(new_n450), .A3(new_n478), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n493), .B(new_n490), .C1(new_n496), .C2(new_n479), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n450), .B1(new_n495), .B2(new_n478), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n188), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(G475), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(KEYINPUT92), .B1(new_n286), .B2(G122), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT92), .ZN(new_n504));
  INV_X1    g318(.A(G122), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n504), .A2(new_n505), .A3(G116), .ZN(new_n506));
  AND2_X1   g320(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(KEYINPUT14), .B1(new_n505), .B2(G116), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT14), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(new_n286), .A3(G122), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(G107), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n503), .A2(new_n506), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n286), .A2(G122), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n273), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n313), .A2(G128), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n206), .A2(G143), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n517), .A3(new_n391), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n391), .B1(new_n516), .B2(new_n517), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n512), .B(new_n515), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n206), .A2(G143), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT13), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n391), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT13), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n524), .A2(new_n525), .B1(new_n518), .B2(KEYINPUT93), .ZN(new_n526));
  OR2_X1    g340(.A1(new_n518), .A2(KEYINPUT93), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n513), .A2(new_n273), .A3(new_n514), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n273), .B1(new_n513), .B2(new_n514), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n526), .B(new_n527), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT94), .ZN(new_n531));
  INV_X1    g345(.A(new_n445), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n187), .A2(G953), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR4_X1   g348(.A1(new_n445), .A2(KEYINPUT94), .A3(new_n187), .A4(G953), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n521), .A2(new_n530), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n536), .B1(new_n521), .B2(new_n530), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n537), .A2(new_n538), .A3(G902), .ZN(new_n539));
  INV_X1    g353(.A(G478), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n540), .A2(KEYINPUT15), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n539), .B(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n502), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n370), .A2(new_n444), .A3(new_n448), .A4(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT72), .ZN(new_n546));
  INV_X1    g360(.A(new_n293), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n393), .A2(G134), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n421), .B1(new_n548), .B2(new_n407), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n371), .B(new_n550), .C1(new_n405), .C2(new_n410), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n551), .B1(new_n425), .B2(new_n325), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT30), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n411), .A2(new_n324), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT30), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(new_n555), .A3(new_n551), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n547), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n551), .B(new_n547), .C1(new_n425), .C2(new_n325), .ZN(new_n558));
  XNOR2_X1  g372(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT26), .B(G101), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT70), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n463), .A2(G210), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n561), .A2(KEYINPUT70), .ZN(new_n566));
  NOR3_X1   g380(.A1(new_n563), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  OR2_X1    g381(.A1(new_n561), .A2(KEYINPUT70), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n564), .B1(new_n568), .B2(new_n562), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n560), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n565), .B1(new_n563), .B2(new_n566), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n568), .A2(new_n564), .A3(new_n562), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(new_n559), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n558), .A2(new_n574), .A3(KEYINPUT71), .ZN(new_n575));
  AOI21_X1  g389(.A(KEYINPUT71), .B1(new_n558), .B2(new_n574), .ZN(new_n576));
  NOR3_X1   g390(.A1(new_n557), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT31), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n546), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n558), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(KEYINPUT28), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n549), .B1(new_n423), .B2(new_n424), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n411), .A2(new_n324), .B1(new_n583), .B2(new_n371), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT73), .B1(new_n584), .B2(new_n547), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT73), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n552), .A2(new_n586), .A3(new_n293), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n580), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT28), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n582), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n574), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n577), .A2(new_n578), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n552), .A2(KEYINPUT30), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n555), .B1(new_n554), .B2(new_n551), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n293), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n576), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n558), .A2(new_n574), .A3(KEYINPUT71), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n599), .A2(KEYINPUT72), .A3(KEYINPUT31), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n579), .A2(new_n592), .A3(new_n593), .A4(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(G472), .A2(G902), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT74), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT74), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n601), .A2(new_n605), .A3(new_n602), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT75), .B(KEYINPUT32), .Z(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n604), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n601), .A2(KEYINPUT32), .A3(new_n602), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n591), .B1(new_n557), .B2(new_n580), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT29), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n590), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n613), .B1(new_n614), .B2(new_n574), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT76), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n552), .A2(new_n293), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n589), .B1(new_n617), .B2(new_n558), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(new_n581), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n574), .A2(KEYINPUT29), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n616), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  NOR4_X1   g436(.A1(new_n618), .A2(new_n581), .A3(KEYINPUT76), .A4(new_n620), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n188), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(G472), .B1(new_n615), .B2(new_n624), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n610), .A2(new_n625), .ZN(new_n626));
  AOI211_X1 g440(.A(new_n253), .B(new_n545), .C1(new_n609), .C2(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(new_n281), .ZN(G3));
  NAND2_X1  g442(.A1(new_n601), .A2(new_n188), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(G472), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n447), .B1(new_n438), .B2(new_n443), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n604), .A2(new_n630), .A3(new_n606), .A4(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n253), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT95), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT97), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n540), .A2(G902), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT96), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n637), .B1(new_n536), .B2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n537), .A2(new_n640), .A3(new_n538), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n521), .A2(new_n530), .ZN(new_n642));
  INV_X1    g456(.A(new_n536), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n521), .A2(new_n530), .A3(new_n536), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n639), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n635), .B(new_n636), .C1(new_n641), .C2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n636), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n640), .B1(new_n537), .B2(new_n538), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n644), .A2(new_n645), .A3(new_n639), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(KEYINPUT97), .B1(new_n539), .B2(G478), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n647), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(KEYINPUT98), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT98), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n647), .B(new_n655), .C1(new_n651), .C2(new_n652), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n370), .A2(new_n502), .A3(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n634), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT34), .B(G104), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G6));
  NOR3_X1   g476(.A1(new_n489), .A2(KEYINPUT20), .A3(new_n491), .ZN(new_n663));
  AOI22_X1  g477(.A1(new_n663), .A2(KEYINPUT99), .B1(new_n500), .B2(G475), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT99), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n492), .A2(new_n497), .A3(new_n665), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n664), .A2(new_n543), .A3(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n634), .A2(new_n370), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT35), .B(G107), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G9));
  INV_X1    g484(.A(new_n632), .ZN(new_n671));
  INV_X1    g485(.A(new_n370), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT101), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n195), .A2(KEYINPUT36), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n221), .A2(new_n230), .A3(KEYINPUT100), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT100), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n677), .B1(new_n237), .B2(new_n242), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n675), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g493(.A(KEYINPUT100), .B1(new_n221), .B2(new_n230), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n237), .A2(new_n242), .A3(new_n677), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n680), .A2(new_n674), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n673), .B1(new_n683), .B2(new_n251), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n251), .ZN(new_n686));
  AOI211_X1 g500(.A(KEYINPUT101), .B(new_n686), .C1(new_n679), .C2(new_n682), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n685), .A2(new_n688), .A3(new_n249), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n544), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n672), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n671), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT37), .B(G110), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G12));
  AND3_X1   g508(.A1(new_n367), .A2(new_n264), .A3(new_n368), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n264), .B1(new_n367), .B2(new_n368), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n254), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n684), .A2(new_n687), .A3(new_n248), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n260), .A2(G900), .A3(new_n192), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT102), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n257), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n700), .A2(new_n701), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  AND4_X1   g519(.A1(new_n543), .A2(new_n664), .A3(new_n666), .A4(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n699), .A2(new_n631), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n707), .B1(new_n609), .B2(new_n626), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(new_n206), .ZN(G30));
  AND3_X1   g523(.A1(new_n502), .A2(new_n254), .A3(new_n543), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n698), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT103), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n695), .A2(new_n696), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(KEYINPUT38), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g529(.A(new_n705), .B(KEYINPUT39), .Z(new_n716));
  AOI211_X1 g530(.A(new_n447), .B(new_n716), .C1(new_n438), .C2(new_n443), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  OR2_X1    g532(.A1(new_n718), .A2(KEYINPUT40), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n574), .B1(new_n617), .B2(new_n558), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n188), .B1(new_n577), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(G472), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n610), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n609), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n718), .A2(KEYINPUT40), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n715), .A2(new_n719), .A3(new_n724), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G143), .ZN(G45));
  INV_X1    g541(.A(new_n705), .ZN(new_n728));
  AOI221_X4 g542(.A(new_n728), .B1(new_n498), .B2(new_n501), .C1(new_n654), .C2(new_n656), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n699), .A3(new_n631), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n601), .A2(new_n605), .A3(new_n602), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n605), .B1(new_n601), .B2(new_n602), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n732), .A2(new_n733), .A3(new_n607), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n610), .A2(new_n625), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n731), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT104), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n609), .A2(new_n626), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(KEYINPUT104), .A3(new_n731), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G146), .ZN(G48));
  INV_X1    g556(.A(new_n253), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n412), .A2(new_n427), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n416), .ZN(new_n745));
  INV_X1    g559(.A(new_n442), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n188), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(G469), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(new_n446), .A3(new_n443), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n739), .A2(new_n743), .A3(new_n659), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(KEYINPUT41), .B(G113), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n752), .B(new_n753), .ZN(G15));
  NAND2_X1  g568(.A1(new_n370), .A2(new_n667), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n750), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n739), .A2(new_n743), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(KEYINPUT105), .B(G116), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(G18));
  NOR2_X1   g573(.A1(new_n750), .A2(new_n697), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n690), .A2(new_n263), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n760), .B(new_n761), .C1(new_n734), .C2(new_n735), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G119), .ZN(G21));
  NAND2_X1  g577(.A1(new_n362), .A2(new_n369), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n710), .A2(new_n764), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n750), .A2(new_n765), .A3(new_n263), .ZN(new_n766));
  INV_X1    g580(.A(G472), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n767), .B1(new_n601), .B2(new_n188), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n599), .A2(KEYINPUT31), .ZN(new_n769));
  OAI21_X1  g583(.A(KEYINPUT106), .B1(new_n618), .B2(new_n581), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n591), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n618), .A2(KEYINPUT106), .A3(new_n581), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n593), .B(new_n769), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n768), .B1(new_n602), .B2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT107), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n253), .B(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n766), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G122), .ZN(G24));
  AOI21_X1  g592(.A(new_n439), .B1(new_n747), .B2(new_n188), .ZN(new_n779));
  INV_X1    g593(.A(new_n443), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n697), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n781), .A2(new_n729), .A3(new_n446), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n773), .A2(new_n602), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n630), .A2(new_n689), .A3(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(new_n198), .ZN(G27));
  AOI21_X1  g601(.A(KEYINPUT32), .B1(new_n601), .B2(new_n602), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n776), .B1(new_n735), .B2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT108), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n776), .B(KEYINPUT108), .C1(new_n735), .C2(new_n788), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n446), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n764), .A2(new_n794), .A3(new_n255), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n729), .A2(new_n795), .A3(new_n444), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT42), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n796), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n739), .A2(new_n743), .A3(new_n799), .ZN(new_n800));
  AOI22_X1  g614(.A1(new_n793), .A2(new_n798), .B1(new_n800), .B2(new_n797), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(new_n421), .ZN(G33));
  AND3_X1   g616(.A1(new_n795), .A2(new_n706), .A3(new_n444), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n743), .B(new_n803), .C1(new_n734), .C2(new_n735), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G134), .ZN(G36));
  NOR3_X1   g619(.A1(new_n695), .A2(new_n696), .A3(new_n255), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n426), .A2(new_n412), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n436), .A2(new_n416), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT45), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n439), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n812), .B1(new_n811), .B2(new_n810), .ZN(new_n813));
  NAND2_X1  g627(.A1(G469), .A2(G902), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT46), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(new_n443), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n815), .A2(new_n816), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n446), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n820), .A2(new_n716), .ZN(new_n821));
  INV_X1    g635(.A(new_n657), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n822), .A2(new_n502), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(KEYINPUT43), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n732), .A2(new_n733), .A3(new_n768), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n824), .A2(new_n826), .A3(new_n689), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT44), .ZN(new_n828));
  AOI211_X1 g642(.A(new_n807), .B(new_n821), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n827), .A2(new_n828), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(KEYINPUT109), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(G137), .ZN(G39));
  XOR2_X1   g647(.A(new_n820), .B(KEYINPUT47), .Z(new_n834));
  INV_X1    g648(.A(new_n739), .ZN(new_n835));
  AND4_X1   g649(.A1(new_n835), .A2(new_n253), .A3(new_n729), .A4(new_n806), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(new_n196), .ZN(G42));
  INV_X1    g652(.A(KEYINPUT113), .ZN(new_n839));
  AOI211_X1 g653(.A(new_n737), .B(new_n730), .C1(new_n626), .C2(new_n609), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT104), .B1(new_n739), .B2(new_n731), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n708), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n705), .A2(new_n446), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n689), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(new_n444), .A3(new_n710), .A4(new_n764), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n724), .A2(new_n847), .ZN(new_n848));
  OR2_X1    g662(.A1(new_n783), .A2(new_n785), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n843), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n842), .A2(new_n850), .A3(KEYINPUT52), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT52), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n846), .B1(new_n609), .B2(new_n723), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n708), .A2(new_n853), .A3(new_n786), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n852), .B1(new_n741), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n839), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT52), .B1(new_n842), .B2(new_n850), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n741), .A2(new_n854), .A3(new_n852), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n857), .A2(new_n858), .A3(KEYINPUT113), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n785), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n799), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n444), .A2(new_n448), .A3(new_n689), .A4(new_n806), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n543), .A2(new_n728), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n664), .A2(new_n666), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT112), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n664), .A2(KEYINPUT112), .A3(new_n666), .A4(new_n864), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n863), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n870), .B1(new_n734), .B2(new_n735), .ZN(new_n871));
  AND4_X1   g685(.A1(KEYINPUT53), .A2(new_n804), .A3(new_n862), .A4(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n671), .A2(new_n743), .A3(new_n659), .ZN(new_n873));
  INV_X1    g687(.A(new_n545), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n739), .A2(new_n743), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n873), .A2(new_n875), .A3(KEYINPUT110), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT110), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n632), .A2(new_n253), .A3(new_n658), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n877), .B1(new_n627), .B2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n502), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(new_n543), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT111), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n882), .A2(new_n672), .ZN(new_n883));
  AOI22_X1  g697(.A1(new_n633), .A2(new_n883), .B1(new_n671), .B2(new_n691), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n872), .A2(new_n876), .A3(new_n879), .A4(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n752), .A2(new_n757), .A3(new_n777), .A4(new_n762), .ZN(new_n886));
  OAI21_X1  g700(.A(KEYINPUT115), .B1(new_n801), .B2(new_n886), .ZN(new_n887));
  AND4_X1   g701(.A1(new_n752), .A2(new_n757), .A3(new_n762), .A4(new_n777), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n800), .A2(new_n797), .ZN(new_n889));
  INV_X1    g703(.A(new_n792), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT32), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n603), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n892), .A2(new_n625), .A3(new_n610), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT108), .B1(new_n893), .B2(new_n776), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n798), .B1(new_n890), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n889), .A2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT115), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n888), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n885), .B1(new_n887), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n804), .A2(new_n871), .A3(new_n862), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n801), .A2(new_n886), .A3(new_n900), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n879), .A2(new_n876), .A3(new_n884), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n901), .A2(new_n902), .A3(new_n858), .A4(new_n857), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT53), .ZN(new_n904));
  AOI22_X1  g718(.A1(new_n860), .A2(new_n899), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT54), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n901), .A2(new_n902), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n909), .B1(new_n859), .B2(new_n856), .ZN(new_n910));
  OAI21_X1  g724(.A(KEYINPUT114), .B1(new_n910), .B2(KEYINPUT53), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT114), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n857), .A2(KEYINPUT113), .A3(new_n858), .ZN(new_n913));
  AOI21_X1  g727(.A(KEYINPUT113), .B1(new_n857), .B2(new_n858), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n912), .B(new_n904), .C1(new_n915), .C2(new_n909), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n903), .A2(new_n904), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n911), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n908), .B1(new_n918), .B2(KEYINPUT54), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT51), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n779), .A2(new_n780), .A3(new_n448), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n834), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n774), .A2(new_n776), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n824), .A2(new_n257), .ZN(new_n924));
  OR2_X1    g738(.A1(new_n924), .A2(KEYINPUT116), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(KEYINPUT116), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n922), .A2(new_n806), .A3(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n781), .A2(new_n795), .ZN(new_n930));
  OR4_X1    g744(.A1(new_n253), .A2(new_n724), .A3(new_n703), .A4(new_n930), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n931), .A2(new_n502), .A3(new_n657), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n930), .B1(new_n925), .B2(new_n926), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n932), .B1(new_n933), .B2(new_n861), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n751), .A2(new_n714), .A3(new_n255), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n927), .A2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT50), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT50), .B1(new_n927), .B2(new_n935), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n934), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n920), .B1(new_n929), .B2(new_n940), .ZN(new_n941));
  OR2_X1    g755(.A1(new_n938), .A2(new_n939), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n942), .A2(KEYINPUT51), .A3(new_n928), .A4(new_n934), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n927), .A2(new_n760), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n256), .B(KEYINPUT117), .Z(new_n945));
  NAND2_X1  g759(.A1(new_n657), .A2(new_n502), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n944), .B(new_n945), .C1(new_n946), .C2(new_n931), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n933), .A2(new_n793), .ZN(new_n948));
  OR2_X1    g762(.A1(new_n948), .A2(KEYINPUT48), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(KEYINPUT48), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n941), .A2(new_n943), .A3(new_n951), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n919), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(G952), .A2(G953), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n781), .B(KEYINPUT49), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n776), .A2(new_n448), .A3(new_n254), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n955), .A2(new_n714), .A3(new_n956), .A4(new_n823), .ZN(new_n957));
  OAI22_X1  g771(.A1(new_n953), .A2(new_n954), .B1(new_n724), .B2(new_n957), .ZN(G75));
  NOR2_X1   g772(.A1(new_n905), .A2(new_n188), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n959), .A2(G210), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n960), .A2(KEYINPUT56), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n310), .A2(new_n340), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(new_n338), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT55), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  XOR2_X1   g779(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n966));
  NAND2_X1  g780(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  OAI22_X1  g781(.A1(new_n960), .A2(new_n967), .B1(G952), .B2(new_n192), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n965), .A2(new_n968), .ZN(G51));
  NOR2_X1   g783(.A1(new_n192), .A2(G952), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n899), .B1(new_n913), .B2(new_n914), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n903), .A2(new_n904), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(KEYINPUT54), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n907), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n814), .B(KEYINPUT57), .Z(new_n976));
  AND2_X1   g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n747), .ZN(new_n978));
  OAI21_X1  g792(.A(KEYINPUT119), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n905), .A2(new_n188), .A3(new_n813), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n978), .B1(new_n975), .B2(new_n976), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT119), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n970), .B1(new_n979), .B2(new_n983), .ZN(G54));
  AND3_X1   g798(.A1(new_n959), .A2(KEYINPUT58), .A3(G475), .ZN(new_n985));
  INV_X1    g799(.A(new_n489), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n985), .A2(new_n986), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n987), .A2(new_n988), .A3(new_n970), .ZN(G60));
  NOR2_X1   g803(.A1(new_n641), .A2(new_n646), .ZN(new_n990));
  NAND2_X1  g804(.A1(G478), .A2(G902), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT59), .Z(new_n992));
  OAI21_X1  g806(.A(new_n990), .B1(new_n919), .B2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT120), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n990), .A2(new_n992), .ZN(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n996), .B1(new_n974), .B2(new_n907), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n994), .B1(new_n997), .B2(new_n970), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n970), .B1(new_n975), .B2(new_n995), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(KEYINPUT120), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n993), .A2(new_n998), .A3(new_n1000), .ZN(G63));
  INV_X1    g815(.A(KEYINPUT61), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n1002), .A2(KEYINPUT122), .ZN(new_n1003));
  NAND2_X1  g817(.A1(G217), .A2(G902), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(KEYINPUT60), .ZN(new_n1005));
  OAI21_X1  g819(.A(KEYINPUT121), .B1(new_n905), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT121), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1005), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n973), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(new_n250), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1006), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n970), .B1(KEYINPUT122), .B2(new_n1002), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AOI22_X1  g827(.A1(new_n1006), .A2(new_n1009), .B1(new_n682), .B2(new_n679), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1003), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n683), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1003), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n1017), .A2(new_n1018), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1019));
  AND2_X1   g833(.A1(new_n1015), .A2(new_n1019), .ZN(G66));
  INV_X1    g834(.A(new_n262), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n192), .B1(new_n1021), .B2(G224), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n902), .A2(new_n888), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1022), .B1(new_n1023), .B2(new_n192), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n962), .B1(G898), .B2(new_n192), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1025), .B(KEYINPUT123), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n1024), .B(new_n1026), .ZN(G69));
  AOI21_X1  g841(.A(new_n837), .B1(new_n831), .B2(new_n829), .ZN(new_n1028));
  AND2_X1   g842(.A1(new_n896), .A2(new_n804), .ZN(new_n1029));
  NOR3_X1   g843(.A1(new_n842), .A2(new_n708), .A3(new_n786), .ZN(new_n1030));
  INV_X1    g844(.A(new_n793), .ZN(new_n1031));
  OR3_X1    g845(.A1(new_n821), .A2(new_n1031), .A3(new_n765), .ZN(new_n1032));
  NAND4_X1  g846(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .A4(new_n1032), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1033), .A2(new_n192), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n594), .A2(new_n595), .ZN(new_n1035));
  NOR2_X1   g849(.A1(new_n458), .A2(new_n459), .ZN(new_n1036));
  XNOR2_X1  g850(.A(new_n1036), .B(KEYINPUT124), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n1035), .B(new_n1037), .Z(new_n1038));
  INV_X1    g852(.A(new_n1038), .ZN(new_n1039));
  OAI211_X1 g853(.A(new_n1034), .B(new_n1039), .C1(G900), .C2(new_n192), .ZN(new_n1040));
  INV_X1    g854(.A(KEYINPUT126), .ZN(new_n1041));
  NAND2_X1  g855(.A1(G227), .A2(G900), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1042), .A2(G953), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1030), .A2(new_n726), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1044), .A2(KEYINPUT62), .ZN(new_n1045));
  OR2_X1    g859(.A1(new_n1044), .A2(KEYINPUT62), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n882), .A2(new_n946), .ZN(new_n1047));
  AOI211_X1 g861(.A(new_n807), .B(new_n718), .C1(new_n1047), .C2(KEYINPUT125), .ZN(new_n1048));
  NOR2_X1   g862(.A1(new_n835), .A2(new_n253), .ZN(new_n1049));
  OAI211_X1 g863(.A(new_n1048), .B(new_n1049), .C1(KEYINPUT125), .C2(new_n1047), .ZN(new_n1050));
  NAND4_X1  g864(.A1(new_n1028), .A2(new_n1045), .A3(new_n1046), .A4(new_n1050), .ZN(new_n1051));
  NOR2_X1   g865(.A1(new_n1039), .A2(G953), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND4_X1  g867(.A1(new_n1040), .A2(new_n1041), .A3(new_n1043), .A4(new_n1053), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n1043), .A2(new_n1041), .ZN(new_n1055));
  NAND3_X1  g869(.A1(new_n1042), .A2(KEYINPUT126), .A3(G953), .ZN(new_n1056));
  NOR2_X1   g870(.A1(new_n192), .A2(G900), .ZN(new_n1057));
  AOI211_X1 g871(.A(new_n1057), .B(new_n1038), .C1(new_n1033), .C2(new_n192), .ZN(new_n1058));
  INV_X1    g872(.A(new_n1053), .ZN(new_n1059));
  OAI211_X1 g873(.A(new_n1055), .B(new_n1056), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  AND2_X1   g874(.A1(new_n1054), .A2(new_n1060), .ZN(G72));
  NAND2_X1  g875(.A1(G472), .A2(G902), .ZN(new_n1062));
  XOR2_X1   g876(.A(new_n1062), .B(KEYINPUT63), .Z(new_n1063));
  OAI21_X1  g877(.A(new_n1063), .B1(new_n1033), .B2(new_n1023), .ZN(new_n1064));
  NOR2_X1   g878(.A1(new_n557), .A2(new_n580), .ZN(new_n1065));
  XNOR2_X1  g879(.A(new_n1065), .B(KEYINPUT127), .ZN(new_n1066));
  AND2_X1   g880(.A1(new_n1066), .A2(new_n591), .ZN(new_n1067));
  AOI21_X1  g881(.A(new_n970), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g882(.A(new_n1063), .B1(new_n1051), .B2(new_n1023), .ZN(new_n1069));
  NOR2_X1   g883(.A1(new_n1066), .A2(new_n591), .ZN(new_n1070));
  NAND2_X1  g884(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g885(.A1(new_n1068), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g886(.A(new_n1063), .ZN(new_n1073));
  AOI21_X1  g887(.A(new_n1073), .B1(new_n599), .B2(new_n611), .ZN(new_n1074));
  AOI21_X1  g888(.A(new_n1072), .B1(new_n918), .B2(new_n1074), .ZN(G57));
endmodule


