//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1246, new_n1247, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n202), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0003(.A(G1), .ZN(new_n204));
  INV_X1    g0004(.A(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  OAI21_X1  g0010(.A(G50), .B1(G58), .B2(G68), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n205), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT65), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n207), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n210), .B(new_n215), .C1(KEYINPUT1), .C2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XNOR2_X1  g0024(.A(G238), .B(G244), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(G232), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT2), .B(G226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G264), .B(G270), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n228), .B(new_n231), .Z(G358));
  XOR2_X1   g0032(.A(G68), .B(G77), .Z(new_n233));
  XNOR2_X1  g0033(.A(G50), .B(G58), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G351));
  NAND2_X1  g0039(.A1(G33), .A2(G41), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(KEYINPUT66), .ZN(new_n241));
  INV_X1    g0041(.A(KEYINPUT66), .ZN(new_n242));
  NAND3_X1  g0042(.A1(new_n242), .A2(G33), .A3(G41), .ZN(new_n243));
  INV_X1    g0043(.A(new_n213), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n241), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(G41), .ZN(new_n246));
  INV_X1    g0046(.A(G45), .ZN(new_n247));
  AOI21_X1  g0047(.A(G1), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n245), .A2(G274), .A3(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(new_n248), .ZN(new_n250));
  AND2_X1   g0050(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G226), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT3), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G1698), .ZN(new_n258));
  INV_X1    g0058(.A(G223), .ZN(new_n259));
  INV_X1    g0059(.A(G77), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n258), .A2(new_n259), .B1(new_n260), .B2(new_n257), .ZN(new_n261));
  AOI21_X1  g0061(.A(G1698), .B1(new_n255), .B2(new_n256), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n261), .B1(G222), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n244), .A2(new_n240), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n249), .B(new_n252), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  OR2_X1    g0065(.A1(new_n265), .A2(G179), .ZN(new_n266));
  NAND3_X1  g0066(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(new_n213), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n268), .B1(new_n204), .B2(G20), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G50), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n204), .A2(G13), .A3(G20), .ZN(new_n271));
  NOR3_X1   g0071(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n205), .A2(new_n254), .ZN(new_n273));
  INV_X1    g0073(.A(G150), .ZN(new_n274));
  OAI22_X1  g0074(.A1(new_n272), .A2(new_n205), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT68), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT67), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT8), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n276), .B(G58), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G58), .ZN(new_n280));
  OAI211_X1 g0080(.A(KEYINPUT67), .B(KEYINPUT8), .C1(new_n280), .C2(KEYINPUT68), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n277), .B1(new_n278), .B2(G58), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n279), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n254), .A2(G20), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n275), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n268), .ZN(new_n286));
  OAI221_X1 g0086(.A(new_n270), .B1(G50), .B2(new_n271), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G169), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n265), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n266), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G190), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n265), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n293), .B(KEYINPUT71), .ZN(new_n294));
  XOR2_X1   g0094(.A(new_n287), .B(KEYINPUT9), .Z(new_n295));
  AOI21_X1  g0095(.A(new_n295), .B1(G200), .B2(new_n265), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT10), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n295), .B(KEYINPUT70), .ZN(new_n299));
  AOI21_X1  g0099(.A(KEYINPUT10), .B1(new_n265), .B2(G200), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n299), .A2(new_n294), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n291), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G1698), .ZN(new_n303));
  AND2_X1   g0103(.A1(KEYINPUT3), .A2(G33), .ZN(new_n304));
  NOR2_X1   g0104(.A1(KEYINPUT3), .A2(G33), .ZN(new_n305));
  OAI211_X1 g0105(.A(G226), .B(new_n303), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  OAI211_X1 g0106(.A(G232), .B(G1698), .C1(new_n304), .C2(new_n305), .ZN(new_n307));
  NAND2_X1  g0107(.A1(G33), .A2(G97), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n264), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n245), .A2(G238), .A3(new_n250), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n249), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(KEYINPUT13), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n249), .A2(new_n313), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT13), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(new_n317), .A3(new_n311), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n315), .A2(G190), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n271), .ZN(new_n320));
  INV_X1    g0120(.A(G68), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n322), .B(KEYINPUT12), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n284), .A2(G77), .B1(G20), .B2(new_n321), .ZN(new_n324));
  INV_X1    g0124(.A(G50), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n324), .B1(new_n325), .B2(new_n273), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n326), .A2(KEYINPUT11), .A3(new_n268), .ZN(new_n327));
  INV_X1    g0127(.A(new_n269), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n323), .B(new_n327), .C1(new_n321), .C2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT11), .B1(new_n326), .B2(new_n268), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n319), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G200), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(new_n315), .B2(new_n318), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n288), .B1(new_n315), .B2(new_n318), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT14), .ZN(new_n337));
  OAI21_X1  g0137(.A(KEYINPUT72), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NOR3_X1   g0138(.A1(new_n312), .A2(new_n314), .A3(KEYINPUT13), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n317), .B1(new_n316), .B2(new_n311), .ZN(new_n340));
  OAI21_X1  g0140(.A(G169), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT72), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n341), .A2(new_n342), .A3(KEYINPUT14), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n315), .A2(G179), .A3(new_n318), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n336), .A2(new_n337), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n338), .A2(new_n343), .A3(new_n344), .A4(new_n345), .ZN(new_n346));
  XNOR2_X1  g0146(.A(new_n331), .B(KEYINPUT73), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n335), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n304), .A2(new_n305), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n262), .A2(G232), .B1(new_n349), .B2(G107), .ZN(new_n350));
  INV_X1    g0150(.A(G238), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n350), .B1(new_n351), .B2(new_n258), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n310), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n251), .A2(G244), .ZN(new_n354));
  AND3_X1   g0154(.A1(new_n353), .A2(new_n249), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(G190), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n353), .A2(new_n249), .A3(new_n354), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(G200), .ZN(new_n358));
  XNOR2_X1  g0158(.A(KEYINPUT15), .B(G87), .ZN(new_n359));
  INV_X1    g0159(.A(new_n284), .ZN(new_n360));
  OAI22_X1  g0160(.A1(new_n359), .A2(new_n360), .B1(new_n205), .B2(new_n260), .ZN(new_n361));
  XNOR2_X1  g0161(.A(KEYINPUT8), .B(G58), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n362), .A2(new_n273), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n268), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  XOR2_X1   g0164(.A(new_n364), .B(KEYINPUT69), .Z(new_n365));
  NOR2_X1   g0165(.A1(new_n271), .A2(G77), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(new_n269), .B2(G77), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n356), .A2(new_n358), .A3(new_n365), .A4(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n365), .A2(new_n367), .ZN(new_n369));
  INV_X1    g0169(.A(G179), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n355), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n357), .A2(new_n288), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n369), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n302), .A2(new_n348), .A3(new_n368), .A4(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n328), .A2(new_n283), .ZN(new_n375));
  OR2_X1    g0175(.A1(new_n283), .A2(new_n320), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT7), .B1(new_n349), .B2(new_n205), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n255), .A2(KEYINPUT7), .A3(new_n205), .A4(new_n256), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(G68), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n280), .A2(new_n321), .ZN(new_n382));
  NOR2_X1   g0182(.A1(G58), .A2(G68), .ZN(new_n383));
  OAI21_X1  g0183(.A(G20), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n273), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(G159), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(KEYINPUT16), .B1(new_n381), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n255), .A2(new_n205), .A3(new_n256), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT7), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n321), .B1(new_n392), .B2(new_n379), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n384), .A2(new_n386), .A3(KEYINPUT16), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n268), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT74), .ZN(new_n396));
  NOR3_X1   g0196(.A1(new_n389), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  AND3_X1   g0197(.A1(new_n384), .A2(new_n386), .A3(KEYINPUT16), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n286), .B1(new_n381), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT16), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n400), .B1(new_n393), .B2(new_n387), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT74), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n377), .B1(new_n397), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n245), .A2(G232), .A3(new_n250), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n249), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(G226), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(G1698), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(G223), .B2(G1698), .ZN(new_n408));
  INV_X1    g0208(.A(G87), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n408), .A2(new_n349), .B1(new_n254), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT75), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n264), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(G223), .A2(G1698), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n413), .B1(new_n406), .B2(G1698), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n414), .A2(new_n257), .B1(G33), .B2(G87), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT75), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n405), .B1(new_n412), .B2(new_n416), .ZN(new_n417));
  OR2_X1    g0217(.A1(new_n417), .A2(new_n288), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(G179), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT76), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n403), .A2(new_n420), .A3(new_n421), .A4(KEYINPUT18), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n396), .B1(new_n389), .B2(new_n395), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n399), .A2(KEYINPUT74), .A3(new_n401), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n405), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n310), .B1(new_n415), .B2(KEYINPUT75), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n410), .A2(new_n411), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n426), .B(new_n292), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(new_n417), .B2(G200), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n425), .A2(new_n377), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT17), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n425), .A2(KEYINPUT17), .A3(new_n377), .A4(new_n430), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n422), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n403), .A2(new_n420), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT18), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n425), .A2(new_n377), .B1(new_n418), .B2(new_n419), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT18), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n438), .A2(new_n440), .A3(KEYINPUT76), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n435), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n374), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n204), .A2(G45), .ZN(new_n445));
  OR2_X1    g0245(.A1(KEYINPUT5), .A2(G41), .ZN(new_n446));
  NAND2_X1  g0246(.A1(KEYINPUT5), .A2(G41), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n448), .A2(new_n245), .A3(G274), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n247), .A2(G1), .ZN(new_n450));
  AND2_X1   g0250(.A1(KEYINPUT5), .A2(G41), .ZN(new_n451));
  NOR2_X1   g0251(.A1(KEYINPUT5), .A2(G41), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n245), .A2(new_n453), .A3(G264), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(G257), .B(G1698), .C1(new_n304), .C2(new_n305), .ZN(new_n456));
  OAI211_X1 g0256(.A(G250), .B(new_n303), .C1(new_n304), .C2(new_n305), .ZN(new_n457));
  INV_X1    g0257(.A(G294), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n254), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n456), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n461), .A2(KEYINPUT84), .A3(new_n310), .ZN(new_n462));
  AOI21_X1  g0262(.A(KEYINPUT84), .B1(new_n461), .B2(new_n310), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n292), .B(new_n455), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n461), .A2(new_n310), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n455), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n333), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n205), .B(G87), .C1(new_n304), .C2(new_n305), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT22), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT22), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n257), .A2(new_n471), .A3(new_n205), .A4(G87), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT24), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT23), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n475), .B1(new_n205), .B2(G107), .ZN(new_n476));
  INV_X1    g0276(.A(G107), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n477), .A2(KEYINPUT23), .A3(G20), .ZN(new_n478));
  INV_X1    g0278(.A(G116), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n254), .A2(new_n479), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n476), .A2(new_n478), .B1(new_n480), .B2(new_n205), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n473), .A2(new_n474), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n474), .B1(new_n473), .B2(new_n481), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n268), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  XOR2_X1   g0284(.A(KEYINPUT83), .B(KEYINPUT25), .Z(new_n485));
  NOR2_X1   g0285(.A1(new_n271), .A2(G107), .ZN(new_n486));
  XNOR2_X1  g0286(.A(new_n485), .B(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n204), .A2(G33), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n271), .A2(new_n488), .A3(new_n213), .A4(new_n267), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n487), .B1(G107), .B2(new_n490), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n468), .A2(new_n484), .A3(new_n491), .ZN(new_n492));
  OR2_X1    g0292(.A1(new_n445), .A2(G274), .ZN(new_n493));
  INV_X1    g0293(.A(G250), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n445), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n493), .A2(new_n245), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(G244), .B1(new_n304), .B2(new_n305), .ZN(new_n497));
  OAI22_X1  g0297(.A1(new_n497), .A2(new_n303), .B1(new_n254), .B2(new_n479), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT80), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n257), .A2(new_n499), .A3(G238), .A4(new_n303), .ZN(new_n500));
  OAI211_X1 g0300(.A(G238), .B(new_n303), .C1(new_n304), .C2(new_n305), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT80), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n498), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(G190), .B(new_n496), .C1(new_n503), .C2(new_n264), .ZN(new_n504));
  INV_X1    g0304(.A(new_n359), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(new_n271), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n489), .A2(new_n409), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT19), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n284), .A2(new_n508), .A3(G97), .ZN(new_n509));
  NOR2_X1   g0309(.A1(G97), .A2(G107), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n510), .A2(new_n409), .B1(new_n308), .B2(new_n205), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n509), .B1(new_n511), .B2(new_n508), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n257), .A2(KEYINPUT81), .A3(new_n205), .A4(G68), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n205), .B(G68), .C1(new_n304), .C2(new_n305), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT81), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n512), .A2(new_n513), .A3(new_n516), .ZN(new_n517));
  AOI211_X1 g0317(.A(new_n506), .B(new_n507), .C1(new_n517), .C2(new_n268), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n502), .A2(new_n500), .ZN(new_n519));
  INV_X1    g0319(.A(G244), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n520), .B1(new_n255), .B2(new_n256), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n480), .B1(new_n521), .B2(G1698), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n264), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n496), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n504), .B(new_n518), .C1(new_n525), .C2(new_n333), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n288), .B1(new_n523), .B2(new_n524), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n506), .B1(new_n517), .B2(new_n268), .ZN(new_n528));
  OR2_X1    g0328(.A1(new_n489), .A2(new_n359), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n370), .B(new_n496), .C1(new_n503), .C2(new_n264), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n527), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n526), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n455), .B1(new_n462), .B2(new_n463), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G169), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n455), .A2(G179), .A3(new_n465), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n535), .A2(new_n536), .B1(new_n484), .B2(new_n491), .ZN(new_n537));
  NOR3_X1   g0337(.A1(new_n492), .A2(new_n533), .A3(new_n537), .ZN(new_n538));
  OAI211_X1 g0338(.A(G264), .B(G1698), .C1(new_n304), .C2(new_n305), .ZN(new_n539));
  OAI211_X1 g0339(.A(G257), .B(new_n303), .C1(new_n304), .C2(new_n305), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n255), .A2(G303), .A3(new_n256), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n310), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n245), .A2(new_n453), .A3(G270), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n543), .A2(new_n449), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G200), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n320), .A2(new_n479), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(new_n489), .B2(new_n479), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n267), .A2(new_n213), .B1(G20), .B2(new_n479), .ZN(new_n549));
  NAND2_X1  g0349(.A1(G33), .A2(G283), .ZN(new_n550));
  INV_X1    g0350(.A(G97), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n550), .B(new_n205), .C1(G33), .C2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT20), .B1(new_n549), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n549), .A2(KEYINPUT20), .A3(new_n552), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n548), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n543), .A2(G190), .A3(new_n449), .A4(new_n544), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n546), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT82), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n546), .A2(KEYINPUT82), .A3(new_n556), .A4(new_n557), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n245), .A2(new_n453), .ZN(new_n563));
  AOI22_X1  g0363(.A1(G270), .A2(new_n563), .B1(new_n542), .B2(new_n310), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n564), .A2(G179), .A3(new_n449), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n565), .A2(new_n556), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n545), .A2(G169), .ZN(new_n567));
  OAI21_X1  g0367(.A(KEYINPUT21), .B1(new_n567), .B2(new_n556), .ZN(new_n568));
  INV_X1    g0368(.A(new_n555), .ZN(new_n569));
  OAI221_X1 g0369(.A(new_n547), .B1(new_n479), .B2(new_n489), .C1(new_n569), .C2(new_n553), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT21), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n570), .A2(new_n571), .A3(new_n545), .A4(G169), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n566), .B1(new_n568), .B2(new_n572), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n562), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n245), .A2(new_n453), .A3(G257), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n449), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n494), .B1(new_n255), .B2(new_n256), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT4), .ZN(new_n579));
  OAI21_X1  g0379(.A(G1698), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n497), .A2(new_n579), .B1(G33), .B2(G283), .ZN(new_n581));
  AND2_X1   g0381(.A1(KEYINPUT4), .A2(G244), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n303), .B(new_n582), .C1(new_n304), .C2(new_n305), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(KEYINPUT78), .B1(new_n584), .B2(new_n310), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n583), .B(new_n550), .C1(new_n521), .C2(KEYINPUT4), .ZN(new_n586));
  OAI21_X1  g0386(.A(G250), .B1(new_n304), .B2(new_n305), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n303), .B1(new_n587), .B2(KEYINPUT4), .ZN(new_n588));
  OAI211_X1 g0388(.A(KEYINPUT78), .B(new_n310), .C1(new_n586), .C2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n370), .B(new_n577), .C1(new_n585), .C2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT77), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n273), .A2(new_n260), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  XNOR2_X1  g0394(.A(G97), .B(G107), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT6), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n596), .A2(new_n551), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n595), .A2(new_n596), .B1(new_n477), .B2(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n592), .B(new_n594), .C1(new_n598), .C2(new_n205), .ZN(new_n599));
  AND2_X1   g0399(.A1(G97), .A2(G107), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n596), .B1(new_n600), .B2(new_n510), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n477), .A2(KEYINPUT6), .A3(G97), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n205), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(KEYINPUT77), .B1(new_n603), .B2(new_n593), .ZN(new_n604));
  OAI21_X1  g0404(.A(G107), .B1(new_n378), .B2(new_n380), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n599), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n268), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n320), .A2(new_n551), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n489), .B2(new_n551), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n310), .B1(new_n586), .B2(new_n588), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n577), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n288), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n591), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n609), .B1(new_n606), .B2(new_n268), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n576), .B1(new_n584), .B2(new_n310), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(G190), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT78), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n612), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n576), .B1(new_n620), .B2(new_n589), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n616), .B(new_n618), .C1(new_n621), .C2(new_n333), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n615), .A2(new_n622), .A3(KEYINPUT79), .ZN(new_n623));
  AOI21_X1  g0423(.A(KEYINPUT79), .B1(new_n615), .B2(new_n622), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n538), .B(new_n574), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n444), .A2(new_n625), .ZN(G372));
  NAND2_X1  g0426(.A1(new_n438), .A2(new_n440), .ZN(new_n627));
  INV_X1    g0427(.A(new_n335), .ZN(new_n628));
  INV_X1    g0428(.A(new_n373), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n347), .A2(new_n346), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n433), .A2(new_n434), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n627), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n298), .A2(new_n301), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n291), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n591), .A2(new_n614), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n636), .A2(KEYINPUT86), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT86), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n638), .B1(new_n591), .B2(new_n614), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n637), .A2(new_n616), .A3(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n532), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n518), .B1(new_n525), .B2(new_n333), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n642), .A2(KEYINPUT85), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n642), .A2(KEYINPUT85), .B1(G190), .B2(new_n525), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n640), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(KEYINPUT26), .B1(new_n615), .B2(new_n533), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n643), .A2(new_n644), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n468), .A2(new_n484), .A3(new_n491), .ZN(new_n651));
  INV_X1    g0451(.A(new_n573), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n650), .B(new_n651), .C1(new_n652), .C2(new_n537), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n615), .A2(new_n622), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n532), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n649), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n635), .B1(new_n444), .B2(new_n656), .ZN(G369));
  NAND3_X1  g0457(.A1(new_n204), .A2(new_n205), .A3(G13), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(G213), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(G343), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(new_n556), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n652), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n562), .A2(new_n573), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n666), .B1(new_n667), .B2(new_n665), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(G330), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n492), .A2(new_n537), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n484), .A2(new_n491), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n663), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n535), .A2(new_n536), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n672), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n674), .B1(new_n676), .B2(new_n664), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n670), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n573), .A2(new_n663), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n671), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n537), .A2(new_n664), .ZN(new_n681));
  AOI21_X1  g0481(.A(KEYINPUT87), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  AND3_X1   g0482(.A1(new_n680), .A2(KEYINPUT87), .A3(new_n681), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n678), .B1(new_n682), .B2(new_n683), .ZN(G399));
  INV_X1    g0484(.A(KEYINPUT88), .ZN(new_n685));
  INV_X1    g0485(.A(new_n208), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n685), .B1(new_n686), .B2(G41), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n208), .A2(KEYINPUT88), .A3(new_n246), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n510), .A2(new_n409), .A3(new_n479), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n690), .A2(new_n204), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n692), .B1(new_n212), .B2(new_n690), .ZN(new_n693));
  XOR2_X1   g0493(.A(new_n693), .B(KEYINPUT28), .Z(new_n694));
  OAI21_X1  g0494(.A(new_n664), .B1(new_n649), .B2(new_n655), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT29), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT90), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OR3_X1    g0499(.A1(new_n615), .A2(new_n533), .A3(KEYINPUT26), .ZN(new_n700));
  OAI211_X1 g0500(.A(new_n700), .B(new_n532), .C1(new_n653), .C2(new_n654), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n646), .B1(new_n640), .B2(new_n645), .ZN(new_n702));
  OAI211_X1 g0502(.A(KEYINPUT29), .B(new_n664), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n695), .A2(KEYINPUT90), .A3(new_n696), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n466), .A2(new_n370), .A3(new_n545), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n577), .B1(new_n585), .B2(new_n590), .ZN(new_n709));
  INV_X1    g0509(.A(new_n525), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT89), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n613), .A2(new_n536), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n543), .A2(new_n544), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n523), .A2(new_n714), .A3(new_n524), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n712), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT30), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n711), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n459), .B1(new_n262), .B2(G250), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n264), .B1(new_n719), .B2(new_n456), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n449), .A2(new_n454), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n617), .A2(new_n722), .A3(G179), .ZN(new_n723));
  OAI211_X1 g0523(.A(new_n564), .B(new_n496), .C1(new_n264), .C2(new_n503), .ZN(new_n724));
  OAI21_X1  g0524(.A(KEYINPUT89), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(KEYINPUT30), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n663), .B1(new_n718), .B2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT31), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n707), .A2(new_n525), .ZN(new_n730));
  AOI22_X1  g0530(.A1(new_n725), .A2(KEYINPUT30), .B1(new_n709), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n716), .A2(new_n717), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n664), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(KEYINPUT31), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n729), .B(new_n734), .C1(new_n625), .C2(new_n663), .ZN(new_n735));
  AOI22_X1  g0535(.A1(new_n705), .A2(new_n706), .B1(G330), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n694), .B1(new_n736), .B2(G1), .ZN(G364));
  INV_X1    g0537(.A(G13), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G20), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n204), .B1(new_n739), .B2(G45), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n690), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n670), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(G330), .B2(new_n668), .ZN(new_n744));
  INV_X1    g0544(.A(new_n742), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n213), .B1(G20), .B2(new_n288), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n205), .A2(new_n370), .A3(new_n333), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT94), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G190), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G68), .ZN(new_n751));
  XOR2_X1   g0551(.A(KEYINPUT95), .B(KEYINPUT32), .Z(new_n752));
  NOR2_X1   g0552(.A1(new_n205), .A2(G190), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G179), .A2(G200), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(G159), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n752), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n205), .B1(new_n754), .B2(G190), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n551), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  OR3_X1    g0560(.A1(new_n752), .A2(new_n755), .A3(new_n756), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n751), .A2(new_n757), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n749), .A2(new_n292), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n762), .B1(G50), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n205), .A2(new_n292), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n370), .A2(G200), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n753), .A2(new_n766), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n767), .A2(new_n280), .B1(new_n768), .B2(new_n260), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(KEYINPUT93), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n769), .A2(KEYINPUT93), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n333), .A2(G179), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n753), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n477), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n765), .A2(new_n772), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI211_X1 g0576(.A(new_n349), .B(new_n774), .C1(G87), .C2(new_n776), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n764), .A2(new_n770), .A3(new_n771), .A4(new_n777), .ZN(new_n778));
  XNOR2_X1  g0578(.A(KEYINPUT33), .B(G317), .ZN(new_n779));
  AOI22_X1  g0579(.A1(G326), .A2(new_n763), .B1(new_n750), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n755), .B(KEYINPUT96), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G329), .ZN(new_n782));
  INV_X1    g0582(.A(G322), .ZN(new_n783));
  INV_X1    g0583(.A(G311), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n767), .A2(new_n783), .B1(new_n768), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n773), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n785), .B1(G283), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G303), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n349), .B1(new_n775), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n758), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n789), .B1(G294), .B2(new_n790), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n780), .A2(new_n782), .A3(new_n787), .A4(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n747), .B1(new_n778), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(G13), .A2(G33), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(G20), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n746), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n208), .A2(new_n257), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n798), .B(KEYINPUT91), .Z(new_n799));
  AOI22_X1  g0599(.A1(new_n799), .A2(G355), .B1(new_n479), .B2(new_n686), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n686), .A2(new_n257), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(new_n247), .B2(new_n212), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT92), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n803), .A2(new_n804), .B1(new_n247), .B2(new_n235), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n800), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n745), .B(new_n793), .C1(new_n797), .C2(new_n807), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n796), .B(KEYINPUT97), .Z(new_n809));
  OAI21_X1  g0609(.A(new_n808), .B1(new_n668), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n744), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(G396));
  NAND2_X1  g0612(.A1(new_n369), .A2(new_n663), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n368), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n373), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n629), .A2(new_n664), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n794), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n746), .A2(new_n794), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT98), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n742), .B1(G77), .B2(new_n820), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT99), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G283), .A2(new_n750), .B1(new_n763), .B2(G303), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n781), .A2(G311), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n767), .A2(new_n458), .B1(new_n768), .B2(new_n479), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(G107), .B2(new_n776), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n257), .B(new_n759), .C1(G87), .C2(new_n786), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n823), .A2(new_n824), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n767), .ZN(new_n829));
  INV_X1    g0629(.A(new_n768), .ZN(new_n830));
  AOI22_X1  g0630(.A1(G143), .A2(new_n829), .B1(new_n830), .B2(G159), .ZN(new_n831));
  INV_X1    g0631(.A(new_n763), .ZN(new_n832));
  INV_X1    g0632(.A(G137), .ZN(new_n833));
  INV_X1    g0633(.A(new_n750), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n831), .B1(new_n832), .B2(new_n833), .C1(new_n274), .C2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT34), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n349), .B1(new_n786), .B2(G68), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n838), .B1(new_n325), .B2(new_n775), .C1(new_n280), .C2(new_n758), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(G132), .B2(new_n781), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n835), .A2(new_n836), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n828), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n822), .B1(new_n843), .B2(new_n746), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n818), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n695), .A2(new_n817), .ZN(new_n846));
  INV_X1    g0646(.A(new_n817), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n664), .B(new_n847), .C1(new_n649), .C2(new_n655), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n735), .A2(G330), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT100), .Z(new_n852));
  AOI21_X1  g0652(.A(new_n742), .B1(new_n849), .B2(new_n850), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n845), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(G384));
  NOR2_X1   g0655(.A1(new_n739), .A2(new_n204), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n848), .A2(new_n816), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT37), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n377), .B1(new_n389), .B2(new_n395), .ZN(new_n860));
  INV_X1    g0660(.A(new_n661), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n860), .B1(new_n420), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n859), .B1(new_n862), .B2(new_n431), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n403), .A2(new_n861), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n436), .A2(new_n865), .A3(new_n859), .A4(new_n431), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT101), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n866), .A2(new_n867), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n864), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n860), .A2(new_n861), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n442), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT38), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n425), .A2(new_n377), .A3(new_n430), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n875), .A2(new_n439), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n876), .A2(KEYINPUT101), .A3(new_n859), .A4(new_n865), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n866), .A2(new_n867), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n863), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n871), .B1(new_n435), .B2(new_n441), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT38), .ZN(new_n881));
  NOR3_X1   g0681(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n874), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n346), .A2(new_n347), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n347), .A2(new_n663), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n884), .A2(new_n885), .A3(new_n628), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n347), .B(new_n663), .C1(new_n346), .C2(new_n335), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NOR3_X1   g0689(.A1(new_n858), .A2(new_n883), .A3(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n627), .A2(new_n861), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n870), .A2(KEYINPUT38), .A3(new_n873), .ZN(new_n893));
  XNOR2_X1  g0693(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n876), .A2(new_n865), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n877), .A2(new_n878), .B1(new_n895), .B2(KEYINPUT37), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n865), .B1(new_n631), .B2(new_n627), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT39), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n893), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n881), .B1(new_n879), .B2(new_n880), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n899), .B1(new_n893), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT103), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT39), .B1(new_n874), .B2(new_n882), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT103), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n893), .A2(new_n898), .A3(new_n899), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n884), .A2(new_n663), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n903), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n892), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n699), .A2(new_n443), .A3(new_n706), .A4(new_n703), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n635), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n910), .B(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT40), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT79), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n654), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n615), .A2(new_n622), .A3(KEYINPUT79), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n676), .A2(new_n651), .A3(new_n526), .A4(new_n532), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n919), .A2(new_n667), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n918), .A2(new_n920), .A3(new_n664), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT104), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n733), .B2(KEYINPUT31), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n727), .A2(KEYINPUT104), .A3(new_n728), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n921), .A2(new_n923), .A3(new_n734), .A4(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n817), .B1(new_n886), .B2(new_n887), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n914), .B1(new_n883), .B2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT105), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n893), .A2(new_n898), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n925), .A2(KEYINPUT105), .A3(new_n926), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n930), .A2(new_n931), .A3(KEYINPUT40), .A4(new_n932), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n928), .A2(new_n933), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n443), .A2(new_n925), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n936), .A2(G330), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n856), .B1(new_n913), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n913), .B2(new_n938), .ZN(new_n940));
  INV_X1    g0740(.A(new_n598), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n941), .A2(KEYINPUT35), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(KEYINPUT35), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n942), .A2(new_n943), .A3(G116), .A4(new_n214), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT36), .ZN(new_n945));
  NOR3_X1   g0745(.A1(new_n382), .A2(new_n211), .A3(new_n260), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n321), .A2(G50), .ZN(new_n947));
  OAI211_X1 g0747(.A(G1), .B(new_n738), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n940), .A2(new_n945), .A3(new_n948), .ZN(G367));
  NAND2_X1  g0749(.A1(new_n801), .A2(new_n231), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n950), .B(new_n797), .C1(new_n208), .C2(new_n359), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n951), .A2(KEYINPUT108), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(KEYINPUT108), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n952), .A2(new_n745), .A3(new_n953), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n518), .A2(new_n664), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n955), .A2(new_n532), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(new_n645), .B2(new_n955), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n773), .A2(new_n551), .ZN(new_n959));
  INV_X1    g0759(.A(new_n755), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n959), .B1(G317), .B2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(G283), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n961), .B1(new_n962), .B2(new_n768), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n775), .A2(new_n479), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(KEYINPUT46), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n965), .B(new_n349), .C1(new_n788), .C2(new_n767), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n964), .A2(KEYINPUT46), .B1(new_n477), .B2(new_n758), .ZN(new_n967));
  NOR3_X1   g0767(.A1(new_n963), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n968), .B1(new_n458), .B2(new_n834), .C1(new_n784), .C2(new_n832), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT109), .Z(new_n970));
  OAI221_X1 g0770(.A(new_n257), .B1(new_n758), .B2(new_n321), .C1(new_n325), .C2(new_n768), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n775), .A2(new_n280), .B1(new_n755), .B2(new_n833), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n767), .A2(new_n274), .B1(new_n773), .B2(new_n260), .ZN(new_n973));
  NOR3_X1   g0773(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(G143), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n974), .B1(new_n832), .B2(new_n975), .C1(new_n756), .C2(new_n834), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n970), .A2(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT47), .Z(new_n978));
  OAI221_X1 g0778(.A(new_n954), .B1(new_n809), .B2(new_n958), .C1(new_n978), .C2(new_n747), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n640), .A2(new_n663), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n615), .B(new_n622), .C1(new_n616), .C2(new_n664), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OR3_X1    g0782(.A1(new_n982), .A2(new_n683), .A3(new_n682), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT44), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n982), .B1(new_n683), .B2(new_n682), .ZN(new_n985));
  XOR2_X1   g0785(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n986));
  XNOR2_X1  g0786(.A(new_n985), .B(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n670), .B(new_n677), .C1(new_n984), .C2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT44), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n983), .B(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n991), .A2(new_n678), .A3(new_n987), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT107), .ZN(new_n994));
  OR3_X1    g0794(.A1(new_n677), .A2(new_n994), .A3(new_n679), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n994), .B1(new_n677), .B2(new_n679), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n995), .A2(new_n680), .A3(new_n996), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(new_n670), .ZN(new_n998));
  INV_X1    g0798(.A(new_n706), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n998), .B(new_n850), .C1(new_n999), .C2(new_n704), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n736), .B1(new_n993), .B2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n689), .B(KEYINPUT41), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n741), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n982), .A2(new_n671), .A3(new_n679), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT42), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n982), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n615), .B1(new_n1008), .B2(new_n676), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n664), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n1007), .A2(new_n1010), .B1(KEYINPUT43), .B2(new_n958), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT43), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n957), .A2(new_n1012), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n678), .B2(new_n1008), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n678), .A2(new_n1008), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1014), .A2(new_n1018), .A3(new_n1015), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n979), .B1(new_n1004), .B2(new_n1020), .ZN(G387));
  OR2_X1    g0821(.A1(new_n677), .A2(new_n809), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n801), .B1(new_n228), .B2(new_n247), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n799), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n691), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1023), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n362), .A2(G50), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT50), .ZN(new_n1028));
  AOI21_X1  g0828(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1028), .A2(new_n1025), .A3(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n1026), .A2(new_n1030), .B1(new_n477), .B2(new_n686), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n797), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n742), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n776), .A2(G77), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n274), .B2(new_n755), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n349), .B(new_n959), .C1(new_n1035), .C2(KEYINPUT110), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(KEYINPUT110), .B2(new_n1035), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT111), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n758), .A2(new_n359), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n767), .A2(new_n325), .B1(new_n768), .B2(new_n321), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1039), .B(new_n1040), .C1(new_n750), .C2(new_n283), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1038), .B(new_n1041), .C1(new_n756), .C2(new_n832), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n257), .B1(new_n960), .B2(G326), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n775), .A2(new_n458), .B1(new_n758), .B2(new_n962), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(G317), .A2(new_n829), .B1(new_n830), .B2(G303), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n832), .B2(new_n783), .C1(new_n784), .C2(new_n834), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT48), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1044), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n1047), .B2(new_n1046), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT49), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1043), .B1(new_n479), .B2(new_n773), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  AND2_X1   g0851(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1042), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1033), .B1(new_n1053), .B2(new_n746), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n998), .A2(new_n741), .B1(new_n1022), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n736), .A2(new_n998), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1000), .A2(new_n690), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1055), .B1(new_n1056), .B2(new_n1057), .ZN(G393));
  NAND2_X1  g0858(.A1(new_n1008), .A2(new_n796), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n763), .A2(G317), .B1(G311), .B2(new_n829), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT52), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n768), .A2(new_n458), .B1(new_n755), .B2(new_n783), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(G283), .B2(new_n776), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n257), .B(new_n774), .C1(G116), .C2(new_n790), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1063), .B(new_n1064), .C1(new_n834), .C2(new_n788), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n763), .A2(G150), .B1(G159), .B2(new_n829), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT51), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n768), .A2(new_n362), .B1(new_n755), .B2(new_n975), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(G68), .B2(new_n776), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n257), .B1(new_n773), .B2(new_n409), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(G77), .B2(new_n790), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1069), .B(new_n1071), .C1(new_n834), .C2(new_n325), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n1061), .A2(new_n1065), .B1(new_n1067), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n746), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n797), .B1(new_n551), .B2(new_n208), .C1(new_n802), .C2(new_n238), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1059), .A2(new_n742), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n993), .B2(new_n740), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n993), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1000), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n689), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n993), .A2(new_n1000), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1077), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(G390));
  NAND3_X1  g0883(.A1(new_n925), .A2(G330), .A3(new_n926), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n908), .B1(new_n857), .B2(new_n888), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n903), .B2(new_n907), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n664), .B(new_n815), .C1(new_n701), .C2(new_n702), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n816), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n888), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n908), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1090), .A2(new_n1091), .A3(new_n931), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1085), .B1(new_n1087), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1086), .ZN(new_n1095));
  NOR3_X1   g0895(.A1(new_n900), .A2(new_n902), .A3(KEYINPUT103), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n905), .B1(new_n904), .B2(new_n906), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1095), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n926), .A2(new_n735), .A3(G330), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1098), .A2(new_n1099), .A3(new_n1092), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1094), .A2(new_n1100), .A3(new_n741), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n794), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n742), .B1(new_n283), .B2(new_n820), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n767), .A2(new_n479), .B1(new_n758), .B2(new_n260), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT116), .Z(new_n1105));
  OAI21_X1  g0905(.A(new_n349), .B1(new_n775), .B2(new_n409), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n321), .A2(new_n773), .B1(new_n768), .B2(new_n551), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1106), .B(new_n1107), .C1(new_n781), .C2(G294), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n763), .A2(G283), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n750), .A2(G107), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1105), .A2(new_n1108), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(KEYINPUT54), .B(G143), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n830), .A2(new_n1113), .B1(new_n790), .B2(G159), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n834), .B2(new_n833), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n763), .A2(G128), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n781), .A2(G125), .ZN(new_n1118));
  INV_X1    g0918(.A(G132), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n257), .B1(new_n767), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(G50), .B2(new_n786), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n775), .A2(new_n274), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT53), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1117), .A2(new_n1118), .A3(new_n1121), .A4(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1111), .B1(new_n1116), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1103), .B1(new_n1125), .B2(new_n746), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1102), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1101), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n925), .A2(G330), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n735), .A2(G330), .A3(new_n847), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1130), .A2(new_n926), .B1(new_n889), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(KEYINPUT112), .B1(new_n1132), .B2(new_n858), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1131), .A2(new_n889), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n1084), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT112), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1135), .A2(new_n1136), .A3(new_n857), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n925), .A2(G330), .A3(new_n847), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n1138), .A2(new_n889), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1099), .A2(new_n816), .A3(new_n1088), .ZN(new_n1140));
  NOR3_X1   g0940(.A1(new_n1139), .A2(KEYINPUT113), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT113), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n1099), .A2(new_n816), .A3(new_n1088), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1138), .A2(new_n889), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1133), .B(new_n1137), .C1(new_n1141), .C2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n443), .A2(new_n1130), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n911), .A2(new_n635), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1146), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(KEYINPUT114), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1094), .A2(new_n1100), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT114), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1146), .A2(new_n1153), .A3(new_n1149), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n1151), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(KEYINPUT113), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1143), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1135), .A2(new_n857), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n1156), .A2(new_n1157), .B1(new_n1158), .B2(KEYINPUT112), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1148), .B1(new_n1159), .B2(new_n1137), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1160), .A2(new_n1094), .A3(new_n1100), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n690), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1129), .B1(new_n1155), .B2(new_n1162), .ZN(G378));
  AOI21_X1  g0963(.A(new_n745), .B1(new_n325), .B2(new_n819), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT119), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n634), .A2(new_n290), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n287), .A2(new_n861), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n302), .A2(new_n1167), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1169), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1176), .A2(new_n795), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1034), .B1(new_n321), .B2(new_n758), .C1(new_n477), .C2(new_n767), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n349), .A2(new_n246), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n773), .A2(new_n280), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n768), .A2(new_n359), .ZN(new_n1181));
  NOR4_X1   g0981(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .A4(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n781), .A2(G283), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(G97), .A2(new_n750), .B1(new_n763), .B2(G116), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT58), .ZN(new_n1186));
  AOI21_X1  g0986(.A(G50), .B1(new_n254), .B2(new_n246), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n1185), .A2(new_n1186), .B1(new_n1179), .B2(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT117), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(G128), .A2(new_n829), .B1(new_n776), .B2(new_n1113), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT118), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n768), .A2(new_n833), .B1(new_n758), .B2(new_n274), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n763), .B2(G125), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1191), .B(new_n1193), .C1(new_n1119), .C2(new_n834), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n786), .A2(G159), .ZN(new_n1197));
  AOI211_X1 g0997(.A(G33), .B(G41), .C1(new_n960), .C2(G124), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1189), .B1(new_n1186), .B2(new_n1185), .C1(new_n1195), .C2(new_n1199), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1165), .B(new_n1177), .C1(new_n746), .C2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n928), .A2(new_n933), .A3(G330), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1176), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1176), .A2(G330), .A3(new_n928), .A4(new_n933), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(new_n910), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1204), .A2(new_n909), .A3(new_n892), .A4(new_n1205), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1201), .B1(new_n1209), .B2(new_n741), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1161), .A2(new_n1149), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT57), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1211), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n690), .ZN(new_n1215));
  AOI21_X1  g1015(.A(KEYINPUT57), .B1(new_n1211), .B2(new_n1209), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1210), .B1(new_n1215), .B2(new_n1216), .ZN(G375));
  NAND3_X1  g1017(.A1(new_n1159), .A2(new_n1148), .A3(new_n1137), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1151), .A2(new_n1003), .A3(new_n1154), .A4(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n889), .A2(new_n794), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n742), .B1(G68), .B2(new_n820), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n257), .B(new_n1039), .C1(G77), .C2(new_n786), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n781), .A2(G303), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n551), .A2(new_n775), .B1(new_n767), .B2(new_n962), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(G107), .B2(new_n830), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1222), .A2(new_n1223), .A3(new_n1225), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n479), .A2(new_n834), .B1(new_n832), .B2(new_n458), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n1119), .A2(new_n832), .B1(new_n834), .B2(new_n1112), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n349), .B(new_n1180), .C1(G50), .C2(new_n790), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n781), .A2(G128), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n833), .A2(new_n767), .B1(new_n775), .B2(new_n756), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(G150), .B2(new_n830), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1229), .A2(new_n1230), .A3(new_n1232), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n1226), .A2(new_n1227), .B1(new_n1228), .B2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1221), .B1(new_n1234), .B2(new_n746), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1146), .A2(new_n741), .B1(new_n1220), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1219), .A2(new_n1236), .ZN(G381));
  NOR4_X1   g1037(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1162), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1151), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1128), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1082), .B(new_n979), .C1(new_n1004), .C2(new_n1020), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1238), .A2(new_n1241), .A3(new_n1243), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1244), .A2(G375), .ZN(G407));
  NAND2_X1  g1045(.A1(new_n1241), .A2(new_n662), .ZN(new_n1246));
  OAI211_X1 g1046(.A(G407), .B(G213), .C1(G375), .C2(new_n1246), .ZN(new_n1247));
  XOR2_X1   g1047(.A(new_n1247), .B(KEYINPUT120), .Z(G409));
  INV_X1    g1048(.A(KEYINPUT123), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(G387), .A2(G390), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(G393), .B(G396), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n1250), .A2(new_n1242), .A3(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1251), .B1(new_n1250), .B2(new_n1242), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1249), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1250), .A2(new_n1242), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1251), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1250), .A2(new_n1242), .A3(new_n1251), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1257), .A2(KEYINPUT123), .A3(new_n1258), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1254), .A2(new_n1259), .A3(KEYINPUT124), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT124), .B1(new_n1254), .B2(new_n1259), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  OAI211_X1 g1062(.A(G378), .B(new_n1210), .C1(new_n1215), .C2(new_n1216), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1211), .A2(new_n1209), .A3(new_n1003), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n1210), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1241), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1263), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT60), .ZN(new_n1268));
  OR2_X1    g1068(.A1(new_n1218), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1218), .A2(new_n1268), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1269), .A2(new_n690), .A3(new_n1150), .A4(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1236), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n854), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1271), .A2(G384), .A3(new_n1236), .ZN(new_n1274));
  AND2_X1   g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n662), .A2(G213), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1267), .A2(new_n1275), .A3(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT121), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1267), .A2(KEYINPUT121), .A3(new_n1275), .A4(new_n1276), .ZN(new_n1280));
  AOI21_X1  g1080(.A(KEYINPUT62), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1267), .A2(new_n1276), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT122), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1273), .A2(new_n1283), .A3(new_n1274), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1283), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n662), .A2(G213), .A3(G2897), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1284), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1275), .A2(new_n1283), .A3(new_n1286), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1282), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1277), .A2(KEYINPUT62), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT61), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1290), .A2(new_n1291), .A3(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1262), .B1(new_n1281), .B2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT63), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1277), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1279), .A2(new_n1295), .A3(new_n1280), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1298), .A2(new_n1299), .A3(new_n1292), .A4(new_n1290), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1294), .A2(new_n1300), .ZN(G405));
  INV_X1    g1101(.A(KEYINPUT125), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT126), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1275), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1305));
  OAI21_X1  g1105(.A(KEYINPUT126), .B1(new_n1305), .B2(KEYINPUT125), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1304), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(G375), .A2(new_n1241), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1307), .A2(new_n1263), .A3(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1263), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1304), .A2(new_n1310), .A3(new_n1306), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1309), .A2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1254), .A2(new_n1259), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1309), .A2(new_n1259), .A3(new_n1254), .A4(new_n1311), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(G402));
endmodule


