//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 1 1 1 1 1 1 1 1 1 1 0 1 0 1 1 1 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n557, new_n559,
    new_n560, new_n561, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n572, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n608, new_n609, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1149,
    new_n1150, new_n1151;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT67), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT68), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT70), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n462), .B(new_n463), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT69), .B(G2105), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(new_n466), .A3(G137), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n465), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n468));
  OAI211_X1 g043(.A(new_n464), .B(new_n467), .C1(new_n468), .C2(new_n466), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(G160));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT3), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT71), .ZN(new_n478));
  OAI221_X1 g053(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n466), .C2(G112), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n475), .A2(new_n466), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n478), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  AND2_X1   g058(.A1(G126), .A2(G2105), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n472), .A2(new_n474), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT72), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n465), .A2(KEYINPUT72), .A3(new_n484), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  AND2_X1   g065(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n491));
  NOR2_X1   g066(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n472), .B(new_n474), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G114), .C2(new_n461), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n465), .A2(new_n466), .A3(KEYINPUT4), .A4(G138), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n489), .A2(new_n495), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  XOR2_X1   g081(.A(KEYINPUT73), .B(G88), .Z(new_n507));
  AOI22_X1  g082(.A1(new_n506), .A2(new_n507), .B1(G50), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT6), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  OR3_X1    g088(.A1(new_n508), .A2(KEYINPUT74), .A3(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n515), .A2(new_n509), .ZN(new_n516));
  OAI21_X1  g091(.A(KEYINPUT74), .B1(new_n508), .B2(new_n513), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n514), .A2(new_n516), .A3(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  INV_X1    g094(.A(KEYINPUT75), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n513), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT6), .B(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT75), .ZN(new_n523));
  AND3_X1   g098(.A1(new_n521), .A2(new_n523), .A3(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G51), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT76), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n526), .A2(G89), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(G89), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n522), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G63), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n530), .B2(new_n509), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(new_n506), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n525), .A2(new_n532), .A3(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  NAND2_X1  g111(.A1(new_n524), .A2(G52), .ZN(new_n537));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n505), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G651), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n505), .A2(new_n513), .ZN(new_n542));
  XNOR2_X1  g117(.A(KEYINPUT77), .B(G90), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n537), .A2(new_n541), .A3(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(G171));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n505), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n542), .A2(G81), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n521), .A2(new_n523), .A3(G543), .ZN(new_n552));
  INV_X1    g127(.A(G43), .ZN(new_n553));
  OAI211_X1 g128(.A(new_n550), .B(new_n551), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT78), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n557), .A2(new_n561), .ZN(G188));
  NAND3_X1  g137(.A1(new_n524), .A2(KEYINPUT9), .A3(G53), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n505), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(G651), .A2(new_n566), .B1(new_n542), .B2(G91), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n552), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n563), .A2(new_n567), .A3(new_n570), .ZN(G299));
  XNOR2_X1  g146(.A(new_n545), .B(KEYINPUT79), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G301));
  NAND4_X1  g148(.A1(new_n521), .A2(new_n523), .A3(G49), .A4(G543), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n542), .A2(G87), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n505), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G651), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT80), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(G48), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G86), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n505), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(new_n522), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n580), .A2(KEYINPUT80), .A3(G651), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n583), .A2(new_n587), .A3(new_n588), .ZN(G305));
  NAND2_X1  g164(.A1(new_n542), .A2(G85), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G47), .ZN(new_n592));
  OAI221_X1 g167(.A(new_n590), .B1(new_n591), .B2(new_n509), .C1(new_n592), .C2(new_n552), .ZN(G290));
  NAND2_X1  g168(.A1(new_n542), .A2(G92), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n594), .B(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n524), .A2(G54), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n506), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n598), .A2(new_n509), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n596), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(new_n572), .B2(new_n601), .ZN(G284));
  OAI21_X1  g178(.A(new_n602), .B1(new_n572), .B2(new_n601), .ZN(G321));
  NAND2_X1  g179(.A1(G299), .A2(new_n601), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(new_n601), .B2(G168), .ZN(G297));
  OAI21_X1  g181(.A(new_n605), .B1(new_n601), .B2(G168), .ZN(G280));
  INV_X1    g182(.A(new_n600), .ZN(new_n608));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G860), .ZN(G148));
  NAND2_X1  g185(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g189(.A1(G123), .A2(new_n480), .B1(new_n476), .B2(G135), .ZN(new_n615));
  OAI221_X1 g190(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n466), .C2(G111), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(KEYINPUT81), .B(G2096), .Z(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT13), .B(G2100), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n619), .A2(new_n623), .ZN(G156));
  INV_X1    g199(.A(G14), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2427), .B(G2438), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2430), .ZN(new_n629));
  INV_X1    g204(.A(KEYINPUT15), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(G2435), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n629), .A2(new_n630), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n629), .A2(new_n630), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(G2435), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n633), .A2(KEYINPUT14), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT83), .B(G2446), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2451), .B(G2454), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2443), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  NAND4_X1  g218(.A1(new_n633), .A2(KEYINPUT14), .A3(new_n636), .A4(new_n638), .ZN(new_n644));
  AND3_X1   g219(.A1(new_n640), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n643), .B1(new_n640), .B2(new_n644), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n627), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n640), .A2(new_n644), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(new_n642), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n640), .A2(new_n643), .A3(new_n644), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(new_n626), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G1341), .B(G1348), .Z(new_n653));
  AOI21_X1  g228(.A(new_n625), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n647), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(KEYINPUT84), .ZN(new_n657));
  INV_X1    g232(.A(KEYINPUT84), .ZN(new_n658));
  NAND4_X1  g233(.A1(new_n647), .A2(new_n651), .A3(new_n658), .A4(new_n655), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n654), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(KEYINPUT85), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT85), .ZN(new_n662));
  NAND4_X1  g237(.A1(new_n654), .A2(new_n657), .A3(new_n662), .A4(new_n659), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(G401));
  XOR2_X1   g240(.A(G2072), .B(G2078), .Z(new_n666));
  XOR2_X1   g241(.A(G2067), .B(G2678), .Z(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n666), .B1(new_n670), .B2(KEYINPUT18), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2096), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G2100), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n670), .A2(KEYINPUT17), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n668), .A2(new_n669), .ZN(new_n675));
  AOI21_X1  g250(.A(KEYINPUT18), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n673), .B(new_n676), .Z(G227));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT86), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT20), .Z(new_n685));
  NOR2_X1   g260(.A1(new_n680), .A2(new_n681), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n687), .A2(new_n679), .A3(new_n682), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n685), .B(new_n688), .C1(new_n679), .C2(new_n687), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G1991), .B(G1996), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(G1981), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1986), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n691), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(G229));
  NAND2_X1  g271(.A1(G299), .A2(G16), .ZN(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G20), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT103), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT23), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT104), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G1956), .ZN(new_n704));
  INV_X1    g279(.A(G2090), .ZN(new_n705));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G35), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G162), .B2(new_n706), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT29), .Z(new_n709));
  OAI21_X1  g284(.A(new_n704), .B1(new_n705), .B2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT105), .ZN(new_n711));
  OR2_X1    g286(.A1(G29), .A2(G32), .ZN(new_n712));
  AOI22_X1  g287(.A1(G129), .A2(new_n480), .B1(new_n476), .B2(G141), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n714));
  NAND3_X1  g289(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT26), .Z(new_n716));
  NAND3_X1  g291(.A1(new_n713), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(KEYINPUT96), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n717), .A2(KEYINPUT96), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n712), .B1(new_n721), .B2(new_n706), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT27), .B(G1996), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT97), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n722), .B(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT99), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G5), .B2(G16), .ZN(new_n727));
  OR3_X1    g302(.A1(new_n726), .A2(G5), .A3(G16), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n727), .B(new_n728), .C1(new_n545), .C2(new_n698), .ZN(new_n729));
  INV_X1    g304(.A(G1961), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT100), .Z(new_n732));
  AND2_X1   g307(.A1(KEYINPUT24), .A2(G34), .ZN(new_n733));
  NOR2_X1   g308(.A1(KEYINPUT24), .A2(G34), .ZN(new_n734));
  NOR3_X1   g309(.A1(new_n733), .A2(new_n734), .A3(G29), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(new_n469), .B2(G29), .ZN(new_n736));
  INV_X1    g311(.A(G2084), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT30), .B(G28), .Z(new_n738));
  OAI22_X1  g313(.A1(new_n736), .A2(new_n737), .B1(G29), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n737), .B2(new_n736), .ZN(new_n740));
  AND3_X1   g315(.A1(new_n725), .A2(new_n732), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(G168), .A2(G16), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G16), .B2(G21), .ZN(new_n743));
  INV_X1    g318(.A(G1966), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n743), .B1(KEYINPUT98), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(KEYINPUT98), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n745), .B(new_n746), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n706), .A2(G33), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT95), .B(KEYINPUT25), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n476), .A2(G139), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n466), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n748), .B1(new_n755), .B2(new_n706), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n756), .A2(G2072), .ZN(new_n757));
  NOR2_X1   g332(.A1(G27), .A2(G29), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G164), .B2(G29), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT101), .ZN(new_n760));
  INV_X1    g335(.A(G2078), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT31), .ZN(new_n763));
  OAI22_X1  g338(.A1(new_n617), .A2(new_n706), .B1(new_n763), .B2(G11), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n763), .B2(G11), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n729), .A2(new_n730), .B1(new_n756), .B2(G2072), .ZN(new_n766));
  AND3_X1   g341(.A1(new_n762), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n741), .A2(new_n747), .A3(new_n757), .A4(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT102), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n767), .A2(new_n757), .ZN(new_n771));
  NAND4_X1  g346(.A1(new_n771), .A2(KEYINPUT102), .A3(new_n747), .A4(new_n741), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n706), .A2(G26), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT28), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n466), .A2(G116), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n775), .A2(new_n471), .ZN(new_n776));
  NOR2_X1   g351(.A1(G104), .A2(G2105), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT93), .Z(new_n778));
  AOI22_X1  g353(.A1(new_n776), .A2(new_n778), .B1(G140), .B2(new_n476), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT92), .ZN(new_n780));
  INV_X1    g355(.A(new_n480), .ZN(new_n781));
  INV_X1    g356(.A(G128), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n480), .A2(KEYINPUT92), .A3(G128), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n779), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(G29), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n786), .A2(KEYINPUT94), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n786), .A2(KEYINPUT94), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n774), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G2067), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n705), .B2(new_n709), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n711), .A2(new_n770), .A3(new_n772), .A4(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT91), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n793), .A2(KEYINPUT36), .ZN(new_n794));
  NOR2_X1   g369(.A1(G16), .A2(G23), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT89), .ZN(new_n796));
  NAND2_X1  g371(.A1(G288), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n574), .A2(new_n575), .A3(KEYINPUT89), .A4(new_n576), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n795), .B1(new_n799), .B2(G16), .ZN(new_n800));
  INV_X1    g375(.A(G1976), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT90), .B(KEYINPUT33), .Z(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n802), .A2(new_n804), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n698), .A2(G22), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G166), .B2(new_n698), .ZN(new_n808));
  INV_X1    g383(.A(G1971), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  MUX2_X1   g385(.A(G6), .B(G305), .S(G16), .Z(new_n811));
  XOR2_X1   g386(.A(KEYINPUT32), .B(G1981), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n805), .A2(new_n806), .A3(new_n810), .A4(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT34), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  MUX2_X1   g391(.A(G24), .B(G290), .S(G16), .Z(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT88), .B(G1986), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n817), .B(new_n818), .Z(new_n819));
  NAND2_X1  g394(.A1(new_n706), .A2(G25), .ZN(new_n820));
  OAI221_X1 g395(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n466), .C2(G107), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT87), .Z(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(G131), .B2(new_n476), .ZN(new_n823));
  INV_X1    g398(.A(G119), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n824), .B2(new_n781), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n820), .B1(new_n826), .B2(new_n706), .ZN(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT35), .B(G1991), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(new_n793), .B2(KEYINPUT36), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n816), .A2(new_n819), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n792), .B1(new_n794), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(G16), .A2(G19), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(new_n555), .B2(G16), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(G1341), .Z(new_n835));
  NAND2_X1  g410(.A1(new_n698), .A2(G4), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n608), .B2(new_n698), .ZN(new_n837));
  INV_X1    g412(.A(G1348), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n831), .A2(new_n794), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n832), .A2(new_n835), .A3(new_n839), .A4(new_n840), .ZN(G150));
  INV_X1    g416(.A(G150), .ZN(G311));
  NAND2_X1  g417(.A1(G80), .A2(G543), .ZN(new_n843));
  INV_X1    g418(.A(G67), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n843), .B1(new_n505), .B2(new_n844), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n845), .A2(G651), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT106), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n524), .A2(G55), .B1(G93), .B2(new_n542), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(G860), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT37), .Z(new_n851));
  NAND2_X1  g426(.A1(new_n608), .A2(G559), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT38), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT39), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n849), .A2(KEYINPUT107), .A3(new_n554), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n554), .A2(KEYINPUT107), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n554), .A2(KEYINPUT107), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n856), .A2(new_n847), .A3(new_n857), .A4(new_n848), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n854), .B(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n851), .B1(new_n860), .B2(G860), .ZN(G145));
  XOR2_X1   g436(.A(new_n621), .B(KEYINPUT109), .Z(new_n862));
  XNOR2_X1  g437(.A(new_n785), .B(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n755), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT108), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n866), .B1(new_n719), .B2(new_n720), .ZN(new_n867));
  OR2_X1    g442(.A1(new_n717), .A2(KEYINPUT96), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n868), .A2(new_n718), .A3(KEYINPUT108), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n865), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n755), .A2(new_n717), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n826), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NOR3_X1   g447(.A1(new_n719), .A2(new_n866), .A3(new_n720), .ZN(new_n873));
  AOI21_X1  g448(.A(KEYINPUT108), .B1(new_n868), .B2(new_n718), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n755), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n871), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(new_n825), .A3(new_n876), .ZN(new_n877));
  AOI22_X1  g452(.A1(G130), .A2(new_n480), .B1(new_n476), .B2(G142), .ZN(new_n878));
  OAI221_X1 g453(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n466), .C2(G118), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n499), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n872), .A2(new_n877), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n882), .B1(new_n872), .B2(new_n877), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n864), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n872), .A2(new_n877), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(new_n881), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n872), .A2(new_n877), .A3(new_n882), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n887), .A2(new_n863), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n617), .B(G160), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(G162), .ZN(new_n892));
  AOI21_X1  g467(.A(G37), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n892), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n885), .A2(new_n889), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(KEYINPUT110), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT110), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n885), .A2(new_n889), .A3(new_n897), .A4(new_n894), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n893), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(KEYINPUT111), .B(KEYINPUT40), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n899), .B(new_n900), .ZN(G395));
  NAND2_X1  g476(.A1(new_n849), .A2(new_n601), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n600), .B(G299), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT41), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n903), .B(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n903), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n855), .A2(new_n858), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(new_n611), .ZN(new_n909));
  MUX2_X1   g484(.A(new_n906), .B(new_n907), .S(new_n909), .Z(new_n910));
  XOR2_X1   g485(.A(G303), .B(G290), .Z(new_n911));
  XNOR2_X1  g486(.A(new_n799), .B(G305), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n911), .B(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(KEYINPUT42), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n910), .B(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n902), .B1(new_n915), .B2(new_n601), .ZN(G295));
  OAI21_X1  g491(.A(new_n902), .B1(new_n915), .B2(new_n601), .ZN(G331));
  NOR2_X1   g492(.A1(G168), .A2(new_n545), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n919), .B1(new_n572), .B2(G286), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT112), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(new_n922), .A3(new_n908), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n859), .A2(new_n920), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT112), .B1(new_n859), .B2(new_n920), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n903), .B1(new_n920), .B2(new_n859), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n921), .A2(new_n908), .ZN(new_n928));
  AOI22_X1  g503(.A1(new_n926), .A2(new_n906), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(G37), .B1(new_n929), .B2(new_n913), .ZN(new_n930));
  INV_X1    g505(.A(new_n913), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n905), .B1(new_n924), .B2(new_n928), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n923), .A2(new_n927), .A3(new_n925), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n930), .A2(KEYINPUT43), .A3(new_n934), .ZN(new_n935));
  OR2_X1    g510(.A1(new_n929), .A2(new_n913), .ZN(new_n936));
  AOI21_X1  g511(.A(KEYINPUT43), .B1(new_n936), .B2(new_n930), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT44), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT43), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n930), .A2(new_n939), .A3(new_n934), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n939), .B1(new_n936), .B2(new_n930), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n938), .B1(new_n942), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g518(.A(G1384), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n495), .A2(new_n497), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT72), .B1(new_n465), .B2(new_n484), .ZN(new_n946));
  AND4_X1   g521(.A1(KEYINPUT72), .A2(new_n472), .A3(new_n474), .A4(new_n484), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n498), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n944), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT45), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(G160), .A2(G40), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n953), .A2(G1996), .A3(new_n717), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT113), .ZN(new_n955));
  OR2_X1    g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n721), .A2(G1996), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n785), .B(G2067), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n953), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n954), .A2(new_n955), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n956), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n953), .ZN(new_n962));
  INV_X1    g537(.A(new_n828), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n825), .B(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n961), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(G290), .B(G1986), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n965), .B1(new_n953), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(G8), .B1(new_n952), .B2(new_n949), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n801), .B1(new_n797), .B2(new_n798), .ZN(new_n969));
  INV_X1    g544(.A(G288), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n970), .A2(G1976), .ZN(new_n971));
  OR4_X1    g546(.A1(KEYINPUT52), .A2(new_n968), .A3(new_n969), .A4(new_n971), .ZN(new_n972));
  OR2_X1    g547(.A1(G305), .A2(G1981), .ZN(new_n973));
  NAND2_X1  g548(.A1(G305), .A2(G1981), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT49), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G8), .ZN(new_n978));
  INV_X1    g553(.A(new_n949), .ZN(new_n979));
  INV_X1    g554(.A(G40), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n469), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n978), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n973), .A2(KEYINPUT49), .A3(new_n974), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n977), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT117), .ZN(new_n985));
  INV_X1    g560(.A(new_n969), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n982), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n985), .B1(new_n987), .B2(KEYINPUT52), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n985), .B(KEYINPUT52), .C1(new_n968), .C2(new_n969), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n972), .B(new_n984), .C1(new_n988), .C2(new_n990), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n944), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT45), .B1(new_n499), .B2(new_n944), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n994), .A2(new_n995), .A3(new_n981), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n944), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n951), .A2(new_n981), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT114), .ZN(new_n999));
  AOI21_X1  g574(.A(G1971), .B1(new_n996), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n949), .A2(KEYINPUT50), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT50), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n499), .A2(new_n1002), .A3(new_n944), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1001), .A2(new_n981), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT115), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n1004), .A2(new_n1005), .A3(G2090), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1000), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1005), .B1(new_n1004), .B2(G2090), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n978), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT116), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1012), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT116), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1014), .A2(new_n1015), .A3(new_n1010), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n991), .B1(new_n1009), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1004), .A2(G2090), .ZN(new_n1019));
  OAI21_X1  g594(.A(G8), .B1(new_n1000), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1018), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1024), .A2(KEYINPUT124), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(G286), .A2(G8), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT119), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n998), .A2(new_n1028), .A3(new_n744), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1028), .B1(new_n998), .B2(new_n744), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1004), .A2(G2084), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1026), .B(new_n1027), .C1(new_n1032), .C2(new_n978), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1024), .A2(KEYINPUT124), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n992), .A2(new_n993), .A3(new_n952), .ZN(new_n1035));
  OAI21_X1  g610(.A(KEYINPUT119), .B1(new_n1035), .B2(G1966), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1004), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n737), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n998), .A2(new_n1028), .A3(new_n744), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1036), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  OAI211_X1 g615(.A(G8), .B(new_n1025), .C1(new_n1040), .C2(G286), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1033), .A2(new_n1034), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT125), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1040), .A2(G8), .A3(G286), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1043), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT62), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT125), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT62), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n998), .A2(new_n1053), .A3(G2078), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1037), .A2(G1961), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n996), .A2(new_n999), .A3(new_n761), .ZN(new_n1056));
  AOI211_X1 g631(.A(new_n1054), .B(new_n1055), .C1(new_n1056), .C2(new_n1053), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1057), .A2(G301), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1047), .A2(new_n1052), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1057), .A2(G301), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1061), .B1(new_n1063), .B2(new_n1058), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1062), .B(KEYINPUT54), .C1(new_n545), .C2(new_n1057), .ZN(new_n1065));
  XNOR2_X1  g640(.A(KEYINPUT56), .B(G2072), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1035), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT57), .B1(new_n567), .B2(KEYINPUT122), .ZN(new_n1068));
  XOR2_X1   g643(.A(G299), .B(new_n1068), .Z(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G1956), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1004), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1067), .A2(new_n1070), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1067), .A2(new_n1072), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n1069), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT61), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1073), .A2(KEYINPUT61), .A3(new_n1075), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n952), .A2(new_n949), .ZN(new_n1080));
  INV_X1    g655(.A(G2067), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1004), .A2(new_n838), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1082), .A2(new_n600), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1082), .A2(new_n600), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT60), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT60), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1082), .A2(new_n1086), .A3(new_n608), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1078), .A2(new_n1079), .A3(new_n1085), .A4(new_n1087), .ZN(new_n1088));
  NOR4_X1   g663(.A1(new_n992), .A2(new_n993), .A3(new_n952), .A4(G1996), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT58), .B(G1341), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1080), .A2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n555), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  XOR2_X1   g667(.A(new_n1092), .B(KEYINPUT59), .Z(new_n1093));
  NAND2_X1  g668(.A1(new_n1073), .A2(new_n1084), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT123), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1094), .A2(new_n1095), .A3(new_n1075), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1095), .B1(new_n1094), .B2(new_n1075), .ZN(new_n1097));
  OAI22_X1  g672(.A1(new_n1088), .A2(new_n1093), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1060), .A2(new_n1064), .A3(new_n1065), .A4(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1023), .B1(new_n1059), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT63), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n995), .B1(new_n994), .B2(new_n981), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n998), .A2(KEYINPUT114), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n809), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1019), .A2(KEYINPUT115), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1104), .A2(new_n1008), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(G8), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1101), .B1(new_n1107), .B2(new_n1021), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n1032), .A2(new_n978), .A3(G286), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1018), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1106), .A2(new_n1017), .A3(G8), .ZN(new_n1111));
  INV_X1    g686(.A(new_n991), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1111), .A2(new_n1112), .A3(new_n1109), .A4(new_n1022), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT120), .B(KEYINPUT63), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1110), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1009), .A2(new_n1112), .A3(new_n1017), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n984), .A2(new_n801), .A3(new_n970), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n973), .B(KEYINPUT118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n982), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1116), .A2(new_n1117), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1116), .A2(KEYINPUT121), .A3(new_n1117), .A4(new_n1120), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n967), .B1(new_n1100), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n961), .A2(new_n963), .A3(new_n826), .ZN(new_n1127));
  OR2_X1    g702(.A1(new_n785), .A2(G2067), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n962), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n962), .A2(G1986), .A3(G290), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1130), .B(KEYINPUT48), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n965), .A2(new_n1131), .ZN(new_n1132));
  OR3_X1    g707(.A1(new_n962), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT46), .B1(new_n962), .B2(G1996), .ZN(new_n1134));
  OR2_X1    g709(.A1(new_n958), .A2(new_n717), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n1133), .A2(new_n1134), .B1(new_n1135), .B2(new_n953), .ZN(new_n1136));
  XOR2_X1   g711(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n1137));
  XNOR2_X1  g712(.A(new_n1136), .B(new_n1137), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1129), .A2(new_n1132), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1126), .A2(new_n1139), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g715(.A1(new_n899), .A2(new_n695), .ZN(new_n1142));
  INV_X1    g716(.A(G227), .ZN(new_n1143));
  NAND3_X1  g717(.A1(new_n664), .A2(G319), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g718(.A1(new_n1144), .A2(KEYINPUT127), .ZN(new_n1145));
  INV_X1    g719(.A(KEYINPUT127), .ZN(new_n1146));
  NAND4_X1  g720(.A1(new_n664), .A2(new_n1146), .A3(G319), .A4(new_n1143), .ZN(new_n1147));
  AOI211_X1 g721(.A(new_n942), .B(new_n1142), .C1(new_n1145), .C2(new_n1147), .ZN(G308));
  NAND2_X1  g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1149));
  INV_X1    g723(.A(new_n942), .ZN(new_n1150));
  INV_X1    g724(.A(new_n1142), .ZN(new_n1151));
  NAND3_X1  g725(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(G225));
endmodule


