

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596;

  XOR2_X1 U322 ( .A(n388), .B(n387), .Z(n528) );
  XOR2_X1 U323 ( .A(n433), .B(n432), .Z(n290) );
  XNOR2_X1 U324 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U325 ( .A(n375), .B(n374), .ZN(n378) );
  XNOR2_X1 U326 ( .A(n478), .B(KEYINPUT48), .ZN(n535) );
  XNOR2_X1 U327 ( .A(n440), .B(n439), .ZN(n441) );
  INV_X1 U328 ( .A(n535), .ZN(n537) );
  XNOR2_X1 U329 ( .A(n442), .B(n441), .ZN(n473) );
  XNOR2_X1 U330 ( .A(n483), .B(KEYINPUT125), .ZN(n484) );
  INV_X1 U331 ( .A(G43GAT), .ZN(n463) );
  XNOR2_X1 U332 ( .A(n485), .B(n484), .ZN(n487) );
  XNOR2_X1 U333 ( .A(n463), .B(KEYINPUT40), .ZN(n464) );
  XNOR2_X1 U334 ( .A(n465), .B(n464), .ZN(G1330GAT) );
  XOR2_X1 U335 ( .A(KEYINPUT66), .B(G71GAT), .Z(n292) );
  XNOR2_X1 U336 ( .A(G99GAT), .B(G43GAT), .ZN(n291) );
  XNOR2_X1 U337 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U338 ( .A(G127GAT), .B(G15GAT), .Z(n418) );
  XOR2_X1 U339 ( .A(n293), .B(n418), .Z(n295) );
  XNOR2_X1 U340 ( .A(G134GAT), .B(G190GAT), .ZN(n294) );
  XNOR2_X1 U341 ( .A(n295), .B(n294), .ZN(n300) );
  XNOR2_X1 U342 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n296) );
  XNOR2_X1 U343 ( .A(n296), .B(G120GAT), .ZN(n348) );
  XOR2_X1 U344 ( .A(n348), .B(G176GAT), .Z(n298) );
  NAND2_X1 U345 ( .A1(G227GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U346 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U347 ( .A(n300), .B(n299), .Z(n308) );
  XOR2_X1 U348 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n302) );
  XNOR2_X1 U349 ( .A(KEYINPUT18), .B(G169GAT), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U351 ( .A(KEYINPUT84), .B(n303), .ZN(n386) );
  XOR2_X1 U352 ( .A(KEYINPUT83), .B(KEYINPUT20), .Z(n305) );
  XNOR2_X1 U353 ( .A(G183GAT), .B(KEYINPUT85), .ZN(n304) );
  XNOR2_X1 U354 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U355 ( .A(n386), .B(n306), .Z(n307) );
  XNOR2_X1 U356 ( .A(n308), .B(n307), .ZN(n571) );
  INV_X1 U357 ( .A(KEYINPUT8), .ZN(n309) );
  NAND2_X1 U358 ( .A1(G43GAT), .A2(n309), .ZN(n311) );
  NAND2_X1 U359 ( .A1(n463), .A2(KEYINPUT8), .ZN(n310) );
  NAND2_X1 U360 ( .A1(n311), .A2(n310), .ZN(n313) );
  XNOR2_X1 U361 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n312) );
  XNOR2_X1 U362 ( .A(n313), .B(n312), .ZN(n445) );
  XOR2_X1 U363 ( .A(KEYINPUT77), .B(G134GAT), .Z(n342) );
  XOR2_X1 U364 ( .A(n445), .B(n342), .Z(n315) );
  NAND2_X1 U365 ( .A1(G232GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U366 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U367 ( .A(G85GAT), .B(G99GAT), .Z(n435) );
  XOR2_X1 U368 ( .A(n316), .B(n435), .Z(n318) );
  XNOR2_X1 U369 ( .A(KEYINPUT10), .B(KEYINPUT65), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U371 ( .A(G92GAT), .B(G106GAT), .Z(n320) );
  XNOR2_X1 U372 ( .A(KEYINPUT9), .B(KEYINPUT11), .ZN(n319) );
  XNOR2_X1 U373 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U374 ( .A(n322), .B(n321), .Z(n327) );
  XOR2_X1 U375 ( .A(G50GAT), .B(KEYINPUT76), .Z(n324) );
  XNOR2_X1 U376 ( .A(G162GAT), .B(G218GAT), .ZN(n323) );
  XNOR2_X1 U377 ( .A(n324), .B(n323), .ZN(n356) );
  XNOR2_X1 U378 ( .A(G36GAT), .B(KEYINPUT78), .ZN(n325) );
  XNOR2_X1 U379 ( .A(n325), .B(G190GAT), .ZN(n376) );
  XNOR2_X1 U380 ( .A(n356), .B(n376), .ZN(n326) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n549) );
  XOR2_X1 U382 ( .A(KEYINPUT36), .B(n549), .Z(n594) );
  INV_X1 U383 ( .A(KEYINPUT101), .ZN(n426) );
  XOR2_X1 U384 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n329) );
  XNOR2_X1 U385 ( .A(G57GAT), .B(G1GAT), .ZN(n328) );
  XNOR2_X1 U386 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U387 ( .A(KEYINPUT4), .B(KEYINPUT92), .Z(n331) );
  XNOR2_X1 U388 ( .A(KEYINPUT91), .B(KEYINPUT6), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U390 ( .A(n333), .B(n332), .Z(n338) );
  XOR2_X1 U391 ( .A(KEYINPUT88), .B(KEYINPUT1), .Z(n335) );
  NAND2_X1 U392 ( .A1(G225GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U393 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U394 ( .A(KEYINPUT5), .B(n336), .ZN(n337) );
  XNOR2_X1 U395 ( .A(n338), .B(n337), .ZN(n346) );
  XOR2_X1 U396 ( .A(G127GAT), .B(G148GAT), .Z(n340) );
  XNOR2_X1 U397 ( .A(G162GAT), .B(G85GAT), .ZN(n339) );
  XNOR2_X1 U398 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U399 ( .A(n341), .B(G155GAT), .Z(n344) );
  XNOR2_X1 U400 ( .A(G29GAT), .B(n342), .ZN(n343) );
  XNOR2_X1 U401 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U402 ( .A(n346), .B(n345), .Z(n350) );
  XNOR2_X1 U403 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n347) );
  XNOR2_X1 U404 ( .A(n347), .B(KEYINPUT2), .ZN(n357) );
  XNOR2_X1 U405 ( .A(n357), .B(n348), .ZN(n349) );
  XNOR2_X1 U406 ( .A(n350), .B(n349), .ZN(n524) );
  XOR2_X1 U407 ( .A(KEYINPUT86), .B(KEYINPUT23), .Z(n352) );
  XNOR2_X1 U408 ( .A(G78GAT), .B(G211GAT), .ZN(n351) );
  XNOR2_X1 U409 ( .A(n352), .B(n351), .ZN(n365) );
  XOR2_X1 U410 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n354) );
  NAND2_X1 U411 ( .A1(G228GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U412 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U413 ( .A(n355), .B(KEYINPUT87), .Z(n359) );
  XNOR2_X1 U414 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U415 ( .A(n359), .B(n358), .ZN(n361) );
  XNOR2_X1 U416 ( .A(G148GAT), .B(G106GAT), .ZN(n360) );
  XNOR2_X1 U417 ( .A(n360), .B(G204GAT), .ZN(n432) );
  XOR2_X1 U418 ( .A(n361), .B(n432), .Z(n363) );
  XOR2_X1 U419 ( .A(G155GAT), .B(G22GAT), .Z(n416) );
  XOR2_X1 U420 ( .A(KEYINPUT21), .B(G197GAT), .Z(n368) );
  XNOR2_X1 U421 ( .A(n416), .B(n368), .ZN(n362) );
  XNOR2_X1 U422 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U423 ( .A(n365), .B(n364), .ZN(n568) );
  XNOR2_X1 U424 ( .A(G211GAT), .B(G183GAT), .ZN(n366) );
  XNOR2_X1 U425 ( .A(n366), .B(G8GAT), .ZN(n413) );
  INV_X1 U426 ( .A(n413), .ZN(n367) );
  NAND2_X1 U427 ( .A1(n368), .A2(n367), .ZN(n371) );
  INV_X1 U428 ( .A(n368), .ZN(n369) );
  NAND2_X1 U429 ( .A1(n369), .A2(n413), .ZN(n370) );
  NAND2_X1 U430 ( .A1(n371), .A2(n370), .ZN(n375) );
  NAND2_X1 U431 ( .A1(G226GAT), .A2(G233GAT), .ZN(n373) );
  INV_X1 U432 ( .A(KEYINPUT93), .ZN(n372) );
  XNOR2_X1 U433 ( .A(n376), .B(G64GAT), .ZN(n377) );
  XNOR2_X1 U434 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U435 ( .A(G92GAT), .B(G176GAT), .Z(n434) );
  XNOR2_X1 U436 ( .A(n379), .B(n434), .ZN(n380) );
  XOR2_X1 U437 ( .A(G218GAT), .B(G204GAT), .Z(n381) );
  NAND2_X1 U438 ( .A1(n380), .A2(n381), .ZN(n385) );
  INV_X1 U439 ( .A(n380), .ZN(n383) );
  INV_X1 U440 ( .A(n381), .ZN(n382) );
  NAND2_X1 U441 ( .A1(n383), .A2(n382), .ZN(n384) );
  NAND2_X1 U442 ( .A1(n385), .A2(n384), .ZN(n388) );
  INV_X1 U443 ( .A(n386), .ZN(n387) );
  NOR2_X1 U444 ( .A1(n571), .A2(n528), .ZN(n389) );
  XOR2_X1 U445 ( .A(KEYINPUT97), .B(n389), .Z(n390) );
  NOR2_X1 U446 ( .A1(n568), .A2(n390), .ZN(n391) );
  XNOR2_X1 U447 ( .A(KEYINPUT25), .B(n391), .ZN(n395) );
  NAND2_X1 U448 ( .A1(n568), .A2(n571), .ZN(n392) );
  XNOR2_X1 U449 ( .A(n392), .B(KEYINPUT26), .ZN(n555) );
  XNOR2_X1 U450 ( .A(n528), .B(KEYINPUT27), .ZN(n398) );
  NOR2_X1 U451 ( .A1(n555), .A2(n398), .ZN(n393) );
  XOR2_X1 U452 ( .A(KEYINPUT96), .B(n393), .Z(n394) );
  NAND2_X1 U453 ( .A1(n395), .A2(n394), .ZN(n396) );
  NAND2_X1 U454 ( .A1(n524), .A2(n396), .ZN(n397) );
  XNOR2_X1 U455 ( .A(n397), .B(KEYINPUT98), .ZN(n404) );
  NOR2_X1 U456 ( .A1(n398), .A2(n524), .ZN(n399) );
  XNOR2_X1 U457 ( .A(n399), .B(KEYINPUT94), .ZN(n536) );
  XOR2_X1 U458 ( .A(KEYINPUT28), .B(KEYINPUT67), .Z(n400) );
  XOR2_X1 U459 ( .A(n568), .B(n400), .Z(n539) );
  NAND2_X1 U460 ( .A1(n536), .A2(n539), .ZN(n401) );
  XNOR2_X1 U461 ( .A(KEYINPUT95), .B(n401), .ZN(n402) );
  NAND2_X1 U462 ( .A1(n402), .A2(n571), .ZN(n403) );
  NAND2_X1 U463 ( .A1(n404), .A2(n403), .ZN(n490) );
  XOR2_X1 U464 ( .A(KEYINPUT71), .B(KEYINPUT72), .Z(n406) );
  XNOR2_X1 U465 ( .A(G64GAT), .B(KEYINPUT13), .ZN(n405) );
  XNOR2_X1 U466 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U467 ( .A(n407), .B(G71GAT), .Z(n409) );
  XNOR2_X1 U468 ( .A(G57GAT), .B(G78GAT), .ZN(n408) );
  XNOR2_X1 U469 ( .A(n409), .B(n408), .ZN(n429) );
  XOR2_X1 U470 ( .A(KEYINPUT79), .B(KEYINPUT14), .Z(n411) );
  XNOR2_X1 U471 ( .A(KEYINPUT15), .B(KEYINPUT82), .ZN(n410) );
  XNOR2_X1 U472 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U473 ( .A(n429), .B(n412), .ZN(n424) );
  XOR2_X1 U474 ( .A(n413), .B(KEYINPUT80), .Z(n415) );
  NAND2_X1 U475 ( .A1(G231GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U476 ( .A(n415), .B(n414), .ZN(n417) );
  XNOR2_X1 U477 ( .A(n417), .B(n416), .ZN(n422) );
  XOR2_X1 U478 ( .A(KEYINPUT81), .B(KEYINPUT12), .Z(n420) );
  XOR2_X1 U479 ( .A(G1GAT), .B(KEYINPUT69), .Z(n446) );
  XNOR2_X1 U480 ( .A(n418), .B(n446), .ZN(n419) );
  XNOR2_X1 U481 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U482 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U483 ( .A(n424), .B(n423), .Z(n591) );
  INV_X1 U484 ( .A(n591), .ZN(n488) );
  NAND2_X1 U485 ( .A1(n490), .A2(n488), .ZN(n425) );
  XNOR2_X1 U486 ( .A(n426), .B(n425), .ZN(n427) );
  NOR2_X1 U487 ( .A1(n594), .A2(n427), .ZN(n428) );
  XNOR2_X1 U488 ( .A(n428), .B(KEYINPUT37), .ZN(n523) );
  XNOR2_X1 U489 ( .A(n429), .B(KEYINPUT31), .ZN(n442) );
  XOR2_X1 U490 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n431) );
  XNOR2_X1 U491 ( .A(G120GAT), .B(KEYINPUT75), .ZN(n430) );
  XNOR2_X1 U492 ( .A(n431), .B(n430), .ZN(n433) );
  XNOR2_X1 U493 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U494 ( .A(n290), .B(n436), .ZN(n440) );
  XOR2_X1 U495 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n438) );
  NAND2_X1 U496 ( .A1(G230GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U497 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U498 ( .A(G197GAT), .B(G169GAT), .Z(n444) );
  XNOR2_X1 U499 ( .A(G141GAT), .B(G22GAT), .ZN(n443) );
  XNOR2_X1 U500 ( .A(n444), .B(n443), .ZN(n459) );
  XOR2_X1 U501 ( .A(n446), .B(n445), .Z(n448) );
  XNOR2_X1 U502 ( .A(G50GAT), .B(G36GAT), .ZN(n447) );
  XNOR2_X1 U503 ( .A(n448), .B(n447), .ZN(n452) );
  XOR2_X1 U504 ( .A(KEYINPUT70), .B(KEYINPUT68), .Z(n450) );
  NAND2_X1 U505 ( .A1(G229GAT), .A2(G233GAT), .ZN(n449) );
  XNOR2_X1 U506 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U507 ( .A(n452), .B(n451), .Z(n457) );
  XOR2_X1 U508 ( .A(KEYINPUT29), .B(G15GAT), .Z(n454) );
  XNOR2_X1 U509 ( .A(G113GAT), .B(G8GAT), .ZN(n453) );
  XNOR2_X1 U510 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U511 ( .A(n455), .B(KEYINPUT30), .ZN(n456) );
  XNOR2_X1 U512 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U513 ( .A(n459), .B(n458), .ZN(n509) );
  NOR2_X1 U514 ( .A1(n473), .A2(n509), .ZN(n493) );
  INV_X1 U515 ( .A(n493), .ZN(n460) );
  NOR2_X1 U516 ( .A1(n523), .A2(n460), .ZN(n462) );
  XOR2_X1 U517 ( .A(KEYINPUT102), .B(KEYINPUT38), .Z(n461) );
  XNOR2_X1 U518 ( .A(n462), .B(n461), .ZN(n505) );
  NOR2_X1 U519 ( .A1(n571), .A2(n505), .ZN(n465) );
  INV_X1 U520 ( .A(n509), .ZN(n585) );
  XOR2_X1 U521 ( .A(n473), .B(KEYINPUT41), .Z(n466) );
  XNOR2_X1 U522 ( .A(n466), .B(KEYINPUT64), .ZN(n508) );
  AND2_X1 U523 ( .A1(n585), .A2(n508), .ZN(n467) );
  XNOR2_X1 U524 ( .A(n467), .B(KEYINPUT46), .ZN(n468) );
  NOR2_X1 U525 ( .A1(n549), .A2(n468), .ZN(n469) );
  XNOR2_X1 U526 ( .A(n591), .B(KEYINPUT111), .ZN(n579) );
  NAND2_X1 U527 ( .A1(n469), .A2(n579), .ZN(n470) );
  XNOR2_X1 U528 ( .A(n470), .B(KEYINPUT47), .ZN(n477) );
  INV_X1 U529 ( .A(KEYINPUT45), .ZN(n472) );
  NOR2_X1 U530 ( .A1(n594), .A2(n488), .ZN(n471) );
  XNOR2_X1 U531 ( .A(n472), .B(n471), .ZN(n475) );
  INV_X1 U532 ( .A(n473), .ZN(n482) );
  NAND2_X1 U533 ( .A1(n482), .A2(n509), .ZN(n474) );
  NOR2_X1 U534 ( .A1(n475), .A2(n474), .ZN(n476) );
  NOR2_X1 U535 ( .A1(n477), .A2(n476), .ZN(n478) );
  NOR2_X1 U536 ( .A1(n535), .A2(n528), .ZN(n479) );
  XNOR2_X1 U537 ( .A(n479), .B(KEYINPUT54), .ZN(n480) );
  NAND2_X1 U538 ( .A1(n480), .A2(n524), .ZN(n567) );
  NOR2_X1 U539 ( .A1(n567), .A2(n555), .ZN(n481) );
  XOR2_X1 U540 ( .A(n481), .B(KEYINPUT122), .Z(n593) );
  OR2_X1 U541 ( .A1(n593), .A2(n482), .ZN(n485) );
  XOR2_X1 U542 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n483) );
  XOR2_X1 U543 ( .A(G204GAT), .B(KEYINPUT124), .Z(n486) );
  XNOR2_X1 U544 ( .A(n487), .B(n486), .ZN(G1353GAT) );
  NOR2_X1 U545 ( .A1(n549), .A2(n488), .ZN(n489) );
  XNOR2_X1 U546 ( .A(KEYINPUT16), .B(n489), .ZN(n491) );
  NAND2_X1 U547 ( .A1(n491), .A2(n490), .ZN(n492) );
  XNOR2_X1 U548 ( .A(n492), .B(KEYINPUT99), .ZN(n510) );
  NAND2_X1 U549 ( .A1(n493), .A2(n510), .ZN(n500) );
  NOR2_X1 U550 ( .A1(n524), .A2(n500), .ZN(n494) );
  XOR2_X1 U551 ( .A(n494), .B(KEYINPUT34), .Z(n495) );
  XNOR2_X1 U552 ( .A(G1GAT), .B(n495), .ZN(G1324GAT) );
  NOR2_X1 U553 ( .A1(n528), .A2(n500), .ZN(n496) );
  XOR2_X1 U554 ( .A(G8GAT), .B(n496), .Z(G1325GAT) );
  NOR2_X1 U555 ( .A1(n571), .A2(n500), .ZN(n498) );
  XNOR2_X1 U556 ( .A(KEYINPUT35), .B(KEYINPUT100), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U558 ( .A(G15GAT), .B(n499), .ZN(G1326GAT) );
  NOR2_X1 U559 ( .A1(n539), .A2(n500), .ZN(n501) );
  XOR2_X1 U560 ( .A(G22GAT), .B(n501), .Z(G1327GAT) );
  NOR2_X1 U561 ( .A1(n524), .A2(n505), .ZN(n503) );
  XNOR2_X1 U562 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n503), .B(n502), .ZN(G1328GAT) );
  NOR2_X1 U564 ( .A1(n528), .A2(n505), .ZN(n504) );
  XOR2_X1 U565 ( .A(G36GAT), .B(n504), .Z(G1329GAT) );
  NOR2_X1 U566 ( .A1(n539), .A2(n505), .ZN(n507) );
  XNOR2_X1 U567 ( .A(G50GAT), .B(KEYINPUT103), .ZN(n506) );
  XNOR2_X1 U568 ( .A(n507), .B(n506), .ZN(G1331GAT) );
  XOR2_X1 U569 ( .A(n508), .B(KEYINPUT105), .Z(n573) );
  NAND2_X1 U570 ( .A1(n573), .A2(n509), .ZN(n522) );
  INV_X1 U571 ( .A(n522), .ZN(n511) );
  NAND2_X1 U572 ( .A1(n511), .A2(n510), .ZN(n518) );
  NOR2_X1 U573 ( .A1(n524), .A2(n518), .ZN(n513) );
  XNOR2_X1 U574 ( .A(KEYINPUT104), .B(KEYINPUT42), .ZN(n512) );
  XNOR2_X1 U575 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U576 ( .A(G57GAT), .B(n514), .Z(G1332GAT) );
  NOR2_X1 U577 ( .A1(n528), .A2(n518), .ZN(n515) );
  XOR2_X1 U578 ( .A(G64GAT), .B(n515), .Z(G1333GAT) );
  NOR2_X1 U579 ( .A1(n571), .A2(n518), .ZN(n516) );
  XOR2_X1 U580 ( .A(KEYINPUT106), .B(n516), .Z(n517) );
  XNOR2_X1 U581 ( .A(G71GAT), .B(n517), .ZN(G1334GAT) );
  NOR2_X1 U582 ( .A1(n539), .A2(n518), .ZN(n520) );
  XNOR2_X1 U583 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U585 ( .A(G78GAT), .B(n521), .Z(G1335GAT) );
  OR2_X1 U586 ( .A1(n523), .A2(n522), .ZN(n532) );
  NOR2_X1 U587 ( .A1(n524), .A2(n532), .ZN(n526) );
  XNOR2_X1 U588 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n525) );
  XNOR2_X1 U589 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U590 ( .A(G85GAT), .B(n527), .ZN(G1336GAT) );
  NOR2_X1 U591 ( .A1(n528), .A2(n532), .ZN(n529) );
  XOR2_X1 U592 ( .A(G92GAT), .B(n529), .Z(G1337GAT) );
  NOR2_X1 U593 ( .A1(n571), .A2(n532), .ZN(n530) );
  XOR2_X1 U594 ( .A(KEYINPUT110), .B(n530), .Z(n531) );
  XNOR2_X1 U595 ( .A(G99GAT), .B(n531), .ZN(G1338GAT) );
  NOR2_X1 U596 ( .A1(n539), .A2(n532), .ZN(n533) );
  XOR2_X1 U597 ( .A(KEYINPUT44), .B(n533), .Z(n534) );
  XNOR2_X1 U598 ( .A(G106GAT), .B(n534), .ZN(G1339GAT) );
  NAND2_X1 U599 ( .A1(n537), .A2(n536), .ZN(n554) );
  NOR2_X1 U600 ( .A1(n571), .A2(n554), .ZN(n538) );
  XNOR2_X1 U601 ( .A(KEYINPUT112), .B(n538), .ZN(n540) );
  NAND2_X1 U602 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U603 ( .A(n541), .B(KEYINPUT113), .Z(n546) );
  INV_X1 U604 ( .A(n546), .ZN(n550) );
  NAND2_X1 U605 ( .A1(n585), .A2(n550), .ZN(n542) );
  XNOR2_X1 U606 ( .A(G113GAT), .B(n542), .ZN(G1340GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n544) );
  NAND2_X1 U608 ( .A1(n550), .A2(n573), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U610 ( .A(G120GAT), .B(n545), .ZN(G1341GAT) );
  NOR2_X1 U611 ( .A1(n579), .A2(n546), .ZN(n547) );
  XOR2_X1 U612 ( .A(KEYINPUT50), .B(n547), .Z(n548) );
  XNOR2_X1 U613 ( .A(G127GAT), .B(n548), .ZN(G1342GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT51), .B(KEYINPUT115), .Z(n552) );
  NAND2_X1 U615 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U616 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U617 ( .A(G134GAT), .B(n553), .Z(G1343GAT) );
  XNOR2_X1 U618 ( .A(G141GAT), .B(KEYINPUT116), .ZN(n557) );
  NOR2_X1 U619 ( .A1(n555), .A2(n554), .ZN(n563) );
  NAND2_X1 U620 ( .A1(n585), .A2(n563), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n557), .B(n556), .ZN(G1344GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n559) );
  NAND2_X1 U623 ( .A1(n563), .A2(n508), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U625 ( .A(G148GAT), .B(n560), .ZN(G1345GAT) );
  XOR2_X1 U626 ( .A(G155GAT), .B(KEYINPUT117), .Z(n562) );
  NAND2_X1 U627 ( .A1(n563), .A2(n591), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1346GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n565) );
  NAND2_X1 U630 ( .A1(n563), .A2(n549), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(G162GAT), .B(n566), .ZN(G1347GAT) );
  NOR2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n569), .B(KEYINPUT55), .ZN(n570) );
  NOR2_X1 U635 ( .A1(n571), .A2(n570), .ZN(n581) );
  NAND2_X1 U636 ( .A1(n581), .A2(n585), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n572), .B(G169GAT), .ZN(G1348GAT) );
  XNOR2_X1 U638 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n577) );
  XOR2_X1 U639 ( .A(G176GAT), .B(KEYINPUT120), .Z(n575) );
  NAND2_X1 U640 ( .A1(n573), .A2(n581), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1349GAT) );
  INV_X1 U643 ( .A(n581), .ZN(n578) );
  NOR2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U645 ( .A(G183GAT), .B(n580), .Z(G1350GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT58), .B(KEYINPUT121), .Z(n583) );
  NAND2_X1 U647 ( .A1(n581), .A2(n549), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(G190GAT), .B(n584), .ZN(G1351GAT) );
  XOR2_X1 U650 ( .A(G197GAT), .B(KEYINPUT60), .Z(n587) );
  INV_X1 U651 ( .A(n593), .ZN(n590) );
  NAND2_X1 U652 ( .A1(n585), .A2(n590), .ZN(n586) );
  XNOR2_X1 U653 ( .A(n587), .B(n586), .ZN(n589) );
  XOR2_X1 U654 ( .A(KEYINPUT123), .B(KEYINPUT59), .Z(n588) );
  XNOR2_X1 U655 ( .A(n589), .B(n588), .ZN(G1352GAT) );
  NAND2_X1 U656 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U657 ( .A(G211GAT), .B(n592), .ZN(G1354GAT) );
  NOR2_X1 U658 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U659 ( .A(KEYINPUT62), .B(n595), .Z(n596) );
  XNOR2_X1 U660 ( .A(G218GAT), .B(n596), .ZN(G1355GAT) );
endmodule

