//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 0 1 1 1 0 1 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n575, new_n576, new_n577, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n593, new_n594, new_n595,
    new_n596, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n453), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n454), .A2(new_n448), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  AOI22_X1  g038(.A1(new_n463), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n467), .B1(new_n468), .B2(G2105), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n465), .A2(KEYINPUT68), .A3(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n465), .A2(G137), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n463), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n466), .A2(new_n475), .ZN(G160));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  AND2_X1   g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(new_n468), .ZN(new_n482));
  NAND2_X1  g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n482), .A2(KEYINPUT69), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(G2105), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n465), .B1(new_n480), .B2(new_n484), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n486), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n493), .A2(new_n495), .A3(G2104), .ZN(new_n496));
  AND2_X1   g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n478), .B2(new_n479), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n501), .B1(new_n478), .B2(new_n479), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n501), .B(new_n504), .C1(new_n479), .C2(new_n478), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n499), .B1(new_n503), .B2(new_n505), .ZN(G164));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n507), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT5), .B(G543), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT70), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n514), .A2(G88), .A3(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  INV_X1    g094(.A(new_n512), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G50), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  OAI21_X1  g099(.A(G62), .B1(new_n508), .B2(new_n509), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n525), .A2(KEYINPUT71), .B1(G75), .B2(G543), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n515), .A2(new_n527), .A3(G62), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n524), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n518), .B(new_n523), .C1(new_n529), .C2(KEYINPUT72), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n525), .A2(KEYINPUT71), .ZN(new_n531));
  NAND2_X1  g106(.A1(G75), .A2(G543), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n528), .ZN(new_n534));
  OAI21_X1  g109(.A(G651), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT72), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n530), .A2(new_n537), .ZN(G166));
  AND2_X1   g113(.A1(new_n514), .A2(new_n517), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G89), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n516), .A2(G543), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(KEYINPUT73), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT73), .ZN(new_n543));
  OAI211_X1 g118(.A(new_n543), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G51), .ZN(new_n546));
  NAND3_X1  g121(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(KEYINPUT7), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(KEYINPUT7), .ZN(new_n549));
  AND2_X1   g124(.A1(G63), .A2(G651), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n548), .A2(new_n549), .B1(new_n515), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n540), .A2(new_n546), .A3(new_n551), .ZN(G286));
  INV_X1    g127(.A(G286), .ZN(G168));
  AOI22_X1  g128(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(new_n524), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  XNOR2_X1  g131(.A(KEYINPUT74), .B(G52), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n543), .B1(new_n516), .B2(G543), .ZN(new_n558));
  INV_X1    g133(.A(new_n544), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n514), .A2(G90), .A3(new_n517), .ZN(new_n561));
  AND3_X1   g136(.A1(new_n560), .A2(new_n561), .A3(KEYINPUT75), .ZN(new_n562));
  AOI21_X1  g137(.A(KEYINPUT75), .B1(new_n560), .B2(new_n561), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n556), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(G171));
  NAND2_X1  g140(.A1(new_n539), .A2(G81), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(new_n524), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n545), .A2(G43), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(G860), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT76), .ZN(G153));
  NAND4_X1  g148(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g149(.A1(G1), .A2(G3), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT8), .ZN(new_n576));
  NAND4_X1  g151(.A1(G319), .A2(G483), .A3(G661), .A4(new_n576), .ZN(new_n577));
  XOR2_X1   g152(.A(new_n577), .B(KEYINPUT77), .Z(G188));
  INV_X1    g153(.A(KEYINPUT9), .ZN(new_n579));
  INV_X1    g154(.A(G53), .ZN(new_n580));
  OAI211_X1 g155(.A(KEYINPUT78), .B(new_n579), .C1(new_n541), .C2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(G78), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G65), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n510), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(G651), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT78), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n580), .B1(new_n586), .B2(KEYINPUT9), .ZN(new_n587));
  OAI211_X1 g162(.A(new_n522), .B(new_n587), .C1(new_n586), .C2(KEYINPUT9), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n581), .A2(new_n585), .A3(new_n588), .ZN(new_n589));
  AND3_X1   g164(.A1(new_n514), .A2(G91), .A3(new_n517), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G299));
  NAND2_X1  g167(.A1(new_n564), .A2(KEYINPUT79), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT79), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n594), .B(new_n556), .C1(new_n562), .C2(new_n563), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G301));
  OR2_X1    g172(.A1(new_n530), .A2(new_n537), .ZN(G303));
  NAND3_X1  g173(.A1(new_n514), .A2(G87), .A3(new_n517), .ZN(new_n599));
  INV_X1    g174(.A(G74), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n510), .A2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G651), .B1(new_n522), .B2(G49), .ZN(new_n602));
  AND2_X1   g177(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G288));
  NAND2_X1  g179(.A1(G73), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G61), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n510), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n607), .A2(G651), .B1(G48), .B2(new_n522), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n514), .A2(G86), .A3(new_n517), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(G305));
  NAND2_X1  g185(.A1(new_n539), .A2(G85), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n612), .A2(new_n524), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n545), .A2(G47), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n611), .A2(new_n613), .A3(new_n614), .ZN(G290));
  INV_X1    g190(.A(G868), .ZN(new_n616));
  NOR2_X1   g191(.A1(G301), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n514), .A2(G92), .A3(new_n517), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT10), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(G79), .A2(G543), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT80), .B(G66), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n510), .B2(new_n622), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n545), .A2(G54), .B1(G651), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT81), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n617), .B1(new_n616), .B2(new_n626), .ZN(G284));
  AOI21_X1  g202(.A(new_n617), .B1(new_n616), .B2(new_n626), .ZN(G321));
  NAND2_X1  g203(.A1(G286), .A2(G868), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(G868), .B2(new_n591), .ZN(G297));
  OAI21_X1  g205(.A(new_n629), .B1(G868), .B2(new_n591), .ZN(G280));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n626), .B1(new_n632), .B2(G860), .ZN(G148));
  NAND2_X1  g208(.A1(new_n626), .A2(new_n632), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  OR3_X1    g210(.A1(new_n635), .A2(KEYINPUT82), .A3(new_n616), .ZN(new_n636));
  OAI21_X1  g211(.A(KEYINPUT82), .B1(new_n635), .B2(new_n616), .ZN(new_n637));
  INV_X1    g212(.A(new_n570), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n636), .B(new_n637), .C1(G868), .C2(new_n638), .ZN(G323));
  XNOR2_X1  g214(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g215(.A1(new_n471), .A2(new_n463), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(KEYINPUT12), .ZN(new_n642));
  INV_X1    g217(.A(KEYINPUT12), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n471), .A2(new_n643), .A3(new_n463), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2100), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT83), .B(KEYINPUT13), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n485), .A2(G135), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n487), .A2(G123), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n465), .A2(G111), .ZN(new_n651));
  OAI21_X1  g226(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n649), .B(new_n650), .C1(new_n651), .C2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(G2096), .Z(new_n654));
  NAND2_X1  g229(.A1(new_n648), .A2(new_n654), .ZN(G156));
  XNOR2_X1  g230(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2427), .B(G2438), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2430), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT15), .B(G2435), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(KEYINPUT14), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(KEYINPUT85), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n663), .A2(KEYINPUT85), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1341), .B(G1348), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n667), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n663), .A2(KEYINPUT85), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n669), .B1(new_n670), .B2(new_n664), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2451), .B(G2454), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2443), .B(G2446), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n672), .B(new_n673), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n668), .A2(new_n671), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n667), .B1(new_n665), .B2(new_n666), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n670), .A2(new_n664), .A3(new_n669), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n674), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n657), .B1(new_n676), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n675), .B1(new_n668), .B2(new_n671), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n677), .A2(new_n674), .A3(new_n678), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n681), .A2(new_n656), .A3(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n680), .A2(G14), .A3(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(G401));
  XNOR2_X1  g260(.A(G2067), .B(G2678), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT86), .ZN(new_n687));
  XNOR2_X1  g262(.A(G2084), .B(G2090), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n689), .A2(KEYINPUT17), .A3(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT88), .B(KEYINPUT18), .Z(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(G2072), .B(G2078), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT87), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n689), .B2(new_n692), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n694), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G2096), .B(G2100), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(new_n700), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(G227));
  XOR2_X1   g278(.A(G1991), .B(G1996), .Z(new_n704));
  XOR2_X1   g279(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n705));
  XNOR2_X1  g280(.A(G1971), .B(G1976), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(G1956), .B(G2474), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1961), .B(G1966), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT20), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n708), .B(new_n709), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n708), .A2(new_n709), .ZN(new_n714));
  MUX2_X1   g289(.A(new_n713), .B(new_n714), .S(new_n707), .Z(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n712), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n716), .B1(new_n712), .B2(new_n715), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n704), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n719), .ZN(new_n721));
  INV_X1    g296(.A(new_n704), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n721), .A2(new_n722), .A3(new_n717), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(G1981), .B(G1986), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n720), .A2(new_n723), .A3(new_n725), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(G229));
  NOR2_X1   g305(.A1(G16), .A2(G24), .ZN(new_n731));
  INV_X1    g306(.A(G290), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(G16), .ZN(new_n733));
  INV_X1    g308(.A(G1986), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n736));
  INV_X1    g311(.A(G107), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n736), .B1(new_n737), .B2(G2105), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n487), .B2(G119), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n485), .A2(G131), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  MUX2_X1   g316(.A(G25), .B(new_n741), .S(G29), .Z(new_n742));
  XOR2_X1   g317(.A(KEYINPUT35), .B(G1991), .Z(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n735), .A2(new_n744), .ZN(new_n745));
  MUX2_X1   g320(.A(G6), .B(G305), .S(G16), .Z(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT32), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G1981), .ZN(new_n748));
  INV_X1    g323(.A(G16), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G23), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n603), .B2(new_n749), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT33), .B(G1976), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT91), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n749), .A2(G22), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G166), .B2(new_n749), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G1971), .ZN(new_n757));
  NOR3_X1   g332(.A1(new_n748), .A2(new_n754), .A3(new_n757), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT90), .B(KEYINPUT34), .Z(new_n759));
  AOI21_X1  g334(.A(new_n745), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n759), .B2(new_n758), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT36), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n638), .A2(new_n749), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n749), .B2(G19), .ZN(new_n764));
  INV_X1    g339(.A(G1341), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OR2_X1    g341(.A1(G104), .A2(G2105), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n767), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT92), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n485), .A2(G140), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n487), .A2(G128), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G29), .ZN(new_n774));
  INV_X1    g349(.A(G29), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n775), .A2(G26), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT28), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n766), .B1(G2067), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n749), .A2(G20), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT23), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n591), .B2(new_n749), .ZN(new_n782));
  OAI22_X1  g357(.A1(new_n782), .A2(G1956), .B1(new_n778), .B2(G2067), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT24), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n784), .A2(G34), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n784), .A2(G34), .ZN(new_n787));
  AOI21_X1  g362(.A(G29), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G160), .B2(new_n775), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(G2084), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n775), .A2(G27), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT100), .Z(new_n793));
  OAI21_X1  g368(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n463), .A2(new_n497), .B1(new_n795), .B2(new_n495), .ZN(new_n796));
  INV_X1    g371(.A(new_n505), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n504), .B1(new_n463), .B2(new_n501), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n793), .B1(new_n799), .B2(G29), .ZN(new_n800));
  INV_X1    g375(.A(G2078), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n790), .A2(G2084), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n791), .A2(new_n802), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  AOI211_X1 g380(.A(new_n783), .B(new_n805), .C1(new_n764), .C2(new_n765), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n782), .A2(G1956), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n779), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n749), .A2(G4), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n626), .B2(new_n749), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1348), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n812), .A2(new_n465), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT93), .ZN(new_n814));
  INV_X1    g389(.A(G139), .ZN(new_n815));
  AOI211_X1 g390(.A(new_n815), .B(G2105), .C1(new_n480), .C2(new_n484), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT25), .ZN(new_n817));
  NAND2_X1  g392(.A1(G103), .A2(G2104), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(G2105), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n465), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n814), .B1(new_n816), .B2(new_n821), .ZN(new_n822));
  NOR3_X1   g397(.A1(new_n478), .A2(new_n479), .A3(new_n477), .ZN(new_n823));
  AOI21_X1  g398(.A(KEYINPUT69), .B1(new_n482), .B2(new_n483), .ZN(new_n824));
  OAI211_X1 g399(.A(G139), .B(new_n465), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n821), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n825), .A2(KEYINPUT93), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n813), .B1(new_n822), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n828), .A2(new_n775), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(new_n775), .B2(G33), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n831), .A2(G2072), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n775), .A2(G35), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(G162), .B2(new_n775), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT29), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n835), .A2(G2090), .ZN(new_n836));
  NOR4_X1   g411(.A1(new_n808), .A2(new_n811), .A3(new_n832), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(G2090), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT101), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n749), .A2(G5), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(G171), .B2(new_n749), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT98), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n842), .A2(G1961), .ZN(new_n843));
  AND2_X1   g418(.A1(new_n831), .A2(G2072), .ZN(new_n844));
  NOR2_X1   g419(.A1(G29), .A2(G32), .ZN(new_n845));
  NAND3_X1  g420(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT26), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(new_n487), .B2(G129), .ZN(new_n848));
  OAI211_X1 g423(.A(G141), .B(new_n465), .C1(new_n823), .C2(new_n824), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n465), .A2(KEYINPUT68), .A3(G2104), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT68), .B1(new_n465), .B2(G2104), .ZN(new_n851));
  OAI21_X1  g426(.A(G105), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(KEYINPUT94), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT94), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n471), .A2(new_n854), .A3(G105), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  AND4_X1   g431(.A1(KEYINPUT95), .A2(new_n848), .A3(new_n849), .A4(new_n856), .ZN(new_n857));
  AOI22_X1  g432(.A1(new_n853), .A2(new_n855), .B1(new_n485), .B2(G141), .ZN(new_n858));
  AOI21_X1  g433(.A(KEYINPUT95), .B1(new_n858), .B2(new_n848), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n845), .B1(new_n860), .B2(G29), .ZN(new_n861));
  XOR2_X1   g436(.A(KEYINPUT27), .B(G1996), .Z(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT96), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n861), .B(new_n863), .ZN(new_n864));
  NOR4_X1   g439(.A1(new_n839), .A2(new_n843), .A3(new_n844), .A4(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(KEYINPUT30), .B(G28), .ZN(new_n866));
  OR2_X1    g441(.A1(KEYINPUT31), .A2(G11), .ZN(new_n867));
  NAND2_X1  g442(.A1(KEYINPUT31), .A2(G11), .ZN(new_n868));
  AOI22_X1  g443(.A1(new_n866), .A2(new_n775), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n749), .A2(G21), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n870), .B1(G168), .B2(new_n749), .ZN(new_n871));
  OAI221_X1 g446(.A(new_n869), .B1(new_n775), .B2(new_n653), .C1(new_n871), .C2(G1966), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(G1966), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(KEYINPUT97), .Z(new_n874));
  AOI211_X1 g449(.A(new_n872), .B(new_n874), .C1(G1961), .C2(new_n842), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n875), .A2(KEYINPUT99), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(KEYINPUT99), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AND4_X1   g453(.A1(new_n762), .A2(new_n837), .A3(new_n865), .A4(new_n878), .ZN(G311));
  NAND4_X1  g454(.A1(new_n762), .A2(new_n837), .A3(new_n865), .A4(new_n878), .ZN(G150));
  NAND2_X1  g455(.A1(G80), .A2(G543), .ZN(new_n881));
  INV_X1    g456(.A(G67), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n881), .B1(new_n510), .B2(new_n882), .ZN(new_n883));
  AOI22_X1  g458(.A1(new_n545), .A2(G55), .B1(G651), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n539), .A2(G93), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(G860), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n887), .B(KEYINPUT37), .Z(new_n888));
  NAND2_X1  g463(.A1(new_n626), .A2(G559), .ZN(new_n889));
  XOR2_X1   g464(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n890));
  XNOR2_X1  g465(.A(new_n889), .B(new_n890), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n570), .A2(new_n886), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n570), .A2(new_n886), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n891), .B(new_n894), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n895), .A2(KEYINPUT39), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n571), .B1(new_n895), .B2(KEYINPUT39), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n888), .B1(new_n896), .B2(new_n897), .ZN(G145));
  INV_X1    g473(.A(KEYINPUT105), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n773), .A2(G164), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n770), .A2(new_n799), .A3(new_n771), .A4(new_n772), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n813), .ZN(new_n904));
  AOI211_X1 g479(.A(new_n814), .B(new_n821), .C1(new_n485), .C2(G139), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT93), .B1(new_n825), .B2(new_n826), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n858), .A2(new_n848), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT95), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n858), .A2(KEYINPUT95), .A3(new_n848), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n907), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n828), .A2(new_n908), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n903), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT104), .ZN(new_n915));
  INV_X1    g490(.A(new_n645), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n741), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n739), .A2(new_n645), .A3(new_n740), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n487), .A2(G130), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT103), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n487), .A2(KEYINPUT103), .A3(G130), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n465), .B1(new_n823), .B2(new_n824), .ZN(new_n925));
  INV_X1    g500(.A(G142), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n465), .A2(G118), .ZN(new_n927));
  OAI21_X1  g502(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n928));
  OAI22_X1  g503(.A1(new_n925), .A2(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n924), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n919), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n929), .B1(new_n922), .B2(new_n923), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n933), .A2(new_n917), .A3(new_n918), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n915), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n828), .B1(new_n857), .B2(new_n859), .ZN(new_n936));
  INV_X1    g511(.A(new_n908), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n907), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n936), .A2(new_n902), .A3(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n914), .A2(new_n935), .A3(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n653), .B(G160), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n941), .B(G162), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n936), .A2(new_n902), .A3(new_n938), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n902), .B1(new_n936), .B2(new_n938), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n933), .A2(new_n917), .A3(new_n918), .ZN(new_n946));
  AOI22_X1  g521(.A1(new_n917), .A2(new_n918), .B1(new_n924), .B2(new_n930), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT104), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n932), .A2(new_n915), .A3(new_n934), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n940), .B(new_n942), .C1(new_n945), .C2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G37), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n948), .B(new_n949), .C1(new_n943), .C2(new_n944), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n942), .B1(new_n954), .B2(new_n940), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n899), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n954), .A2(new_n940), .ZN(new_n957));
  INV_X1    g532(.A(new_n942), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n959), .A2(KEYINPUT105), .A3(new_n952), .A4(new_n951), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n956), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(KEYINPUT40), .ZN(G395));
  AND2_X1   g537(.A1(new_n892), .A2(new_n893), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n634), .B(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT41), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n620), .A2(new_n591), .A3(new_n624), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n591), .B1(new_n620), .B2(new_n624), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n965), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n968), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n970), .A2(KEYINPUT41), .A3(new_n966), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n964), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n967), .A2(new_n968), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n973), .B1(new_n974), .B2(new_n964), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT42), .ZN(new_n976));
  XNOR2_X1  g551(.A(G166), .B(G290), .ZN(new_n977));
  XOR2_X1   g552(.A(new_n603), .B(G305), .Z(new_n978));
  XNOR2_X1  g553(.A(new_n977), .B(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT42), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n973), .B(new_n980), .C1(new_n974), .C2(new_n964), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n976), .A2(new_n979), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n979), .B1(new_n976), .B2(new_n981), .ZN(new_n983));
  OAI21_X1  g558(.A(G868), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n886), .A2(new_n616), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(G295));
  NAND2_X1  g561(.A1(new_n984), .A2(new_n985), .ZN(G331));
  NAND2_X1  g562(.A1(new_n560), .A2(new_n561), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT75), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n560), .A2(new_n561), .A3(KEYINPUT75), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n594), .B1(new_n992), .B2(new_n556), .ZN(new_n993));
  INV_X1    g568(.A(new_n595), .ZN(new_n994));
  OAI21_X1  g569(.A(G168), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n564), .A2(G286), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n995), .A2(new_n963), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT106), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n996), .B1(new_n596), .B2(G168), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1001), .A2(KEYINPUT106), .A3(new_n963), .ZN(new_n1002));
  AOI21_X1  g577(.A(G286), .B1(new_n593), .B2(new_n595), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n894), .B1(new_n1003), .B2(new_n996), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1000), .A2(new_n1002), .A3(new_n974), .A4(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n972), .B1(new_n998), .B2(new_n1004), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n979), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n998), .A2(new_n1004), .A3(new_n974), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1000), .A2(new_n1004), .A3(new_n1002), .ZN(new_n1011));
  INV_X1    g586(.A(new_n972), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1010), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n952), .B(new_n1009), .C1(new_n1013), .C2(new_n1008), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT43), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT106), .B1(new_n1001), .B2(new_n963), .ZN(new_n1017));
  NOR4_X1   g592(.A1(new_n1003), .A2(new_n894), .A3(new_n996), .A4(new_n999), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n1004), .A2(new_n974), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1006), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(G37), .B1(new_n1021), .B2(new_n1008), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1008), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT43), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT44), .B1(new_n1016), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n972), .B1(new_n1019), .B2(new_n1004), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n979), .B1(new_n1027), .B2(new_n1010), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1028), .A2(new_n1022), .A3(new_n1015), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1009), .A2(new_n952), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT43), .B1(new_n1030), .B2(new_n1023), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1026), .B1(new_n1033), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g609(.A(KEYINPUT45), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1035), .B1(G164), .B2(G1384), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n471), .A2(G101), .B1(new_n463), .B2(new_n473), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1037), .B(G40), .C1(new_n465), .C2(new_n464), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1039), .A2(G1996), .A3(new_n908), .ZN(new_n1041));
  XOR2_X1   g616(.A(new_n1041), .B(KEYINPUT108), .Z(new_n1042));
  XOR2_X1   g617(.A(new_n773), .B(G2067), .Z(new_n1043));
  INV_X1    g618(.A(new_n860), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1043), .B1(new_n1044), .B2(G1996), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1042), .B1(new_n1039), .B2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1046), .A2(new_n743), .A3(new_n740), .A4(new_n739), .ZN(new_n1047));
  OR2_X1    g622(.A1(new_n773), .A2(G2067), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1040), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT46), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1050), .B1(new_n1040), .B2(G1996), .ZN(new_n1051));
  XOR2_X1   g626(.A(new_n1051), .B(KEYINPUT125), .Z(new_n1052));
  INV_X1    g627(.A(new_n1043), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n937), .B1(new_n1050), .B2(G1996), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1039), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  XOR2_X1   g631(.A(new_n1056), .B(KEYINPUT47), .Z(new_n1057));
  XNOR2_X1  g632(.A(new_n741), .B(new_n743), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1040), .B1(new_n1059), .B2(KEYINPUT109), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1060), .B1(KEYINPUT109), .B2(new_n1059), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1046), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n732), .A2(new_n1039), .A3(new_n734), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1063), .B(KEYINPUT48), .ZN(new_n1064));
  AOI211_X1 g639(.A(new_n1049), .B(new_n1057), .C1(new_n1062), .C2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G1981), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1066), .B1(new_n608), .B2(new_n609), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n608), .A2(new_n609), .A3(new_n1066), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1068), .A2(KEYINPUT49), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT49), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1069), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1071), .B1(new_n1072), .B2(new_n1067), .ZN(new_n1073));
  INV_X1    g648(.A(G1384), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n799), .A2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1075), .A2(new_n1038), .ZN(new_n1076));
  INV_X1    g651(.A(G8), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1070), .A2(new_n1073), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT111), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n599), .A2(new_n602), .A3(new_n1080), .A4(G1976), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1081), .B(G8), .C1(new_n1075), .C2(new_n1038), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1080), .B1(new_n603), .B2(G1976), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT52), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  OR2_X1    g659(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1085));
  AOI21_X1  g660(.A(G1976), .B1(new_n599), .B2(new_n602), .ZN(new_n1086));
  OR3_X1    g661(.A1(new_n1086), .A2(KEYINPUT112), .A3(KEYINPUT52), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT112), .B1(new_n1086), .B2(KEYINPUT52), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1079), .B(new_n1084), .C1(new_n1085), .C2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n799), .A2(KEYINPUT45), .A3(new_n1074), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1038), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1036), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(G1971), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT50), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n799), .A2(new_n1097), .A3(new_n1074), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1096), .A2(new_n1092), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G2090), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1095), .A2(KEYINPUT110), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1038), .B1(new_n1075), .B2(new_n1035), .ZN(new_n1102));
  AOI21_X1  g677(.A(G1971), .B1(new_n1102), .B2(new_n1091), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT110), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1077), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT55), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(G166), .B2(new_n1077), .ZN(new_n1108));
  OAI211_X1 g683(.A(KEYINPUT55), .B(G8), .C1(new_n530), .C2(new_n537), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1090), .B1(new_n1106), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT113), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1038), .B1(new_n1075), .B2(KEYINPUT50), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1113), .A2(new_n1100), .A3(new_n1098), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1077), .B1(new_n1095), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1112), .B1(new_n1110), .B2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1096), .A2(new_n1092), .A3(new_n1098), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1117), .A2(G2090), .ZN(new_n1118));
  OAI21_X1  g693(.A(G8), .B1(new_n1118), .B2(new_n1103), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1119), .A2(KEYINPUT113), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1116), .A2(new_n1120), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n1111), .A2(new_n1121), .A3(KEYINPUT123), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT123), .B1(new_n1111), .B2(new_n1121), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT51), .ZN(new_n1125));
  INV_X1    g700(.A(G1966), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT114), .B1(new_n1093), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n1117), .A2(G2084), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1093), .A2(KEYINPUT114), .A3(new_n1126), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1077), .B1(new_n1131), .B2(G168), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(G286), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1125), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(G8), .B1(new_n1133), .B2(G286), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1136), .A2(KEYINPUT51), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT62), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1036), .A2(new_n1092), .A3(new_n1091), .A4(new_n801), .ZN(new_n1139));
  XNOR2_X1  g714(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n1140));
  XNOR2_X1  g715(.A(KEYINPUT120), .B(G1961), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1139), .A2(new_n1140), .B1(new_n1117), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1093), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n801), .A2(KEYINPUT53), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1142), .A2(new_n1145), .B1(new_n593), .B2(new_n595), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1137), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT62), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1134), .ZN(new_n1149));
  OAI21_X1  g724(.A(KEYINPUT51), .B1(new_n1149), .B2(new_n1136), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1147), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1124), .A2(new_n1138), .A3(new_n1146), .A4(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT61), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n581), .A2(new_n585), .A3(new_n588), .ZN(new_n1154));
  INV_X1    g729(.A(new_n590), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT57), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1154), .A2(new_n1155), .A3(KEYINPUT116), .A4(new_n1156), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n1156), .A2(KEYINPUT116), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1156), .A2(KEYINPUT116), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1158), .B(new_n1159), .C1(new_n589), .C2(new_n590), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(KEYINPUT115), .B1(new_n1099), .B2(G1956), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT115), .ZN(new_n1164));
  INV_X1    g739(.A(G1956), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1117), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(KEYINPUT56), .B(G2072), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1143), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1162), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  AND3_X1   g745(.A1(new_n1117), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1164), .B1(new_n1117), .B2(new_n1165), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n1169), .B(new_n1162), .C1(new_n1171), .C2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1153), .B1(new_n1170), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT60), .ZN(new_n1176));
  AOI21_X1  g751(.A(G1348), .B1(new_n1113), .B2(new_n1098), .ZN(new_n1177));
  NOR3_X1   g752(.A1(new_n1075), .A2(new_n1038), .A3(G2067), .ZN(new_n1178));
  OAI21_X1  g753(.A(KEYINPUT117), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(G1348), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1178), .B1(new_n1117), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT117), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1176), .B1(new_n1179), .B2(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g759(.A(KEYINPUT58), .B(G1341), .ZN(new_n1185));
  OAI22_X1  g760(.A1(new_n1093), .A2(G1996), .B1(new_n1076), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(new_n638), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1187), .A2(KEYINPUT59), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT59), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1186), .A2(new_n638), .A3(new_n1189), .ZN(new_n1190));
  AOI22_X1  g765(.A1(new_n1184), .A2(new_n625), .B1(new_n1188), .B2(new_n1190), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1177), .A2(KEYINPUT117), .A3(new_n1178), .ZN(new_n1193));
  OAI21_X1  g768(.A(KEYINPUT60), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(new_n625), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1179), .A2(new_n1183), .A3(new_n1176), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  AOI22_X1  g772(.A1(new_n1163), .A2(new_n1166), .B1(new_n1143), .B2(new_n1168), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT118), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n1161), .B(new_n1199), .ZN(new_n1200));
  OAI211_X1 g775(.A(KEYINPUT61), .B(new_n1173), .C1(new_n1198), .C2(new_n1200), .ZN(new_n1201));
  NAND4_X1  g776(.A1(new_n1175), .A2(new_n1191), .A3(new_n1197), .A4(new_n1201), .ZN(new_n1202));
  NAND4_X1  g777(.A1(new_n1173), .A2(new_n1195), .A3(new_n1183), .A4(new_n1179), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n1161), .B(KEYINPUT118), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1203), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT119), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1203), .A2(new_n1206), .A3(KEYINPUT119), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1202), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT54), .ZN(new_n1212));
  INV_X1    g787(.A(KEYINPUT122), .ZN(new_n1213));
  AOI21_X1  g788(.A(KEYINPUT45), .B1(new_n799), .B2(new_n1074), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1213), .B1(new_n1214), .B2(new_n1038), .ZN(new_n1215));
  NAND3_X1  g790(.A1(new_n1036), .A2(KEYINPUT122), .A3(new_n1092), .ZN(new_n1216));
  NAND4_X1  g791(.A1(new_n1215), .A2(new_n1216), .A3(new_n1091), .A4(new_n1144), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1142), .A2(new_n1217), .ZN(new_n1218));
  NOR2_X1   g793(.A1(new_n1218), .A2(new_n596), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1212), .B1(new_n1219), .B2(new_n1146), .ZN(new_n1220));
  AOI21_X1  g795(.A(new_n1212), .B1(new_n1218), .B2(G171), .ZN(new_n1221));
  NAND3_X1  g796(.A1(G301), .A2(new_n1142), .A3(new_n1145), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1220), .A2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1224), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1225));
  NAND3_X1  g800(.A1(new_n1211), .A2(new_n1124), .A3(new_n1225), .ZN(new_n1226));
  NOR2_X1   g801(.A1(G288), .A2(G1976), .ZN(new_n1227));
  AND2_X1   g802(.A1(new_n1079), .A2(new_n1227), .ZN(new_n1228));
  OAI21_X1  g803(.A(new_n1078), .B1(new_n1228), .B2(new_n1072), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1106), .A2(new_n1110), .ZN(new_n1230));
  OAI21_X1  g805(.A(new_n1229), .B1(new_n1230), .B2(new_n1090), .ZN(new_n1231));
  NOR3_X1   g806(.A1(new_n1131), .A2(new_n1077), .A3(G286), .ZN(new_n1232));
  NAND3_X1  g807(.A1(new_n1232), .A2(new_n1111), .A3(new_n1121), .ZN(new_n1233));
  INV_X1    g808(.A(KEYINPUT63), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  OR2_X1    g810(.A1(new_n1106), .A2(new_n1110), .ZN(new_n1236));
  NAND4_X1  g811(.A1(new_n1236), .A2(new_n1232), .A3(new_n1111), .A4(KEYINPUT63), .ZN(new_n1237));
  AOI21_X1  g812(.A(new_n1231), .B1(new_n1235), .B2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g813(.A1(new_n1152), .A2(new_n1226), .A3(new_n1238), .ZN(new_n1239));
  INV_X1    g814(.A(KEYINPUT124), .ZN(new_n1240));
  NAND3_X1  g815(.A1(new_n1039), .A2(G1986), .A3(G290), .ZN(new_n1241));
  NAND2_X1  g816(.A1(new_n1063), .A2(new_n1241), .ZN(new_n1242));
  XNOR2_X1  g817(.A(new_n1242), .B(KEYINPUT107), .ZN(new_n1243));
  AND2_X1   g818(.A1(new_n1062), .A2(new_n1243), .ZN(new_n1244));
  AND3_X1   g819(.A1(new_n1239), .A2(new_n1240), .A3(new_n1244), .ZN(new_n1245));
  AOI21_X1  g820(.A(new_n1240), .B1(new_n1239), .B2(new_n1244), .ZN(new_n1246));
  OAI21_X1  g821(.A(new_n1065), .B1(new_n1245), .B2(new_n1246), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g822(.A(KEYINPUT126), .ZN(new_n1249));
  AOI21_X1  g823(.A(new_n461), .B1(new_n701), .B2(new_n702), .ZN(new_n1250));
  AND3_X1   g824(.A1(new_n684), .A2(new_n729), .A3(new_n1250), .ZN(new_n1251));
  NAND2_X1  g825(.A1(new_n961), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g826(.A(new_n1252), .ZN(new_n1253));
  AOI21_X1  g827(.A(new_n1249), .B1(new_n1032), .B2(new_n1253), .ZN(new_n1254));
  AOI211_X1 g828(.A(KEYINPUT126), .B(new_n1252), .C1(new_n1029), .C2(new_n1031), .ZN(new_n1255));
  NOR2_X1   g829(.A1(new_n1254), .A2(new_n1255), .ZN(G308));
  NOR2_X1   g830(.A1(new_n1014), .A2(KEYINPUT43), .ZN(new_n1257));
  AOI21_X1  g831(.A(new_n1015), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1258));
  OAI21_X1  g832(.A(new_n1253), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g833(.A1(new_n1259), .A2(KEYINPUT126), .ZN(new_n1260));
  NAND3_X1  g834(.A1(new_n1032), .A2(new_n1249), .A3(new_n1253), .ZN(new_n1261));
  NAND2_X1  g835(.A1(new_n1260), .A2(new_n1261), .ZN(G225));
endmodule


