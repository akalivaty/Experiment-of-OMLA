//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 1 0 1 0 1 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0 1 0 1 0 1 0 0 0 0 0 0 1 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1 1 0 1 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n827, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1029, new_n1030;
  AOI21_X1  g000(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(G29gat), .ZN(new_n203));
  INV_X1    g002(.A(G36gat), .ZN(new_n204));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NOR2_X1   g004(.A1(G29gat), .A2(G36gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(KEYINPUT14), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT15), .ZN(new_n211));
  AND2_X1   g010(.A1(KEYINPUT82), .A2(G43gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(KEYINPUT82), .A2(G43gat), .ZN(new_n213));
  NOR3_X1   g012(.A1(new_n212), .A2(new_n213), .A3(G50gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT83), .ZN(new_n215));
  INV_X1    g014(.A(G50gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(G43gat), .ZN(new_n217));
  INV_X1    g016(.A(G43gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n218), .A2(KEYINPUT83), .A3(G50gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n211), .B1(new_n214), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT15), .B1(new_n216), .B2(G43gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n218), .A2(G50gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n210), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n225), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT17), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT17), .ZN(new_n230));
  XNOR2_X1  g029(.A(KEYINPUT82), .B(G43gat), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n217), .B(new_n219), .C1(new_n231), .C2(G50gat), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n224), .B1(new_n232), .B2(new_n211), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n230), .B(new_n227), .C1(new_n233), .C2(new_n210), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n229), .A2(new_n234), .ZN(new_n235));
  AND2_X1   g034(.A1(G99gat), .A2(G106gat), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT8), .ZN(new_n237));
  OAI22_X1  g036(.A1(new_n236), .A2(new_n237), .B1(G85gat), .B2(G92gat), .ZN(new_n238));
  OR2_X1    g037(.A1(KEYINPUT90), .A2(KEYINPUT7), .ZN(new_n239));
  AND2_X1   g038(.A1(G85gat), .A2(G92gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(KEYINPUT90), .A2(KEYINPUT7), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G85gat), .A2(G92gat), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT91), .B1(new_n243), .B2(KEYINPUT7), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n238), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  OR2_X1    g044(.A1(G99gat), .A2(G106gat), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT92), .ZN(new_n247));
  NAND2_X1  g046(.A1(G99gat), .A2(G106gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(G99gat), .A2(G106gat), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT92), .B1(new_n236), .B2(new_n250), .ZN(new_n251));
  AND2_X1   g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n239), .A2(new_n240), .A3(KEYINPUT91), .A4(new_n241), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n245), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G85gat), .ZN(new_n255));
  INV_X1    g054(.A(G92gat), .ZN(new_n256));
  AOI22_X1  g055(.A1(KEYINPUT8), .A2(new_n248), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AND2_X1   g056(.A1(KEYINPUT90), .A2(KEYINPUT7), .ZN(new_n258));
  NOR2_X1   g057(.A1(KEYINPUT90), .A2(KEYINPUT7), .ZN(new_n259));
  NOR3_X1   g058(.A1(new_n258), .A2(new_n259), .A3(new_n243), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT91), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT7), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n261), .B1(new_n240), .B2(new_n262), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n253), .B(new_n257), .C1(new_n260), .C2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n249), .A2(new_n251), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n254), .A2(new_n266), .A3(KEYINPUT93), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT93), .B1(new_n254), .B2(new_n266), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n235), .A2(new_n269), .A3(KEYINPUT94), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT93), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n252), .B1(new_n245), .B2(new_n253), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n264), .A2(new_n265), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n254), .A2(new_n266), .A3(KEYINPUT93), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n274), .A2(new_n229), .A3(new_n275), .A4(new_n234), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT94), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n226), .A2(new_n228), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n279), .B1(new_n267), .B2(new_n268), .ZN(new_n280));
  NAND3_X1  g079(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n270), .A2(new_n278), .A3(new_n280), .A4(new_n281), .ZN(new_n282));
  XOR2_X1   g081(.A(G190gat), .B(G218gat), .Z(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT96), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n282), .A2(KEYINPUT96), .A3(new_n284), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G162gat), .ZN(new_n290));
  AND3_X1   g089(.A1(new_n270), .A2(new_n278), .A3(new_n281), .ZN(new_n291));
  NAND4_X1  g090(.A1(new_n291), .A2(KEYINPUT95), .A3(new_n283), .A4(new_n280), .ZN(new_n292));
  INV_X1    g091(.A(new_n281), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n293), .B1(new_n276), .B2(new_n277), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n294), .A2(new_n283), .A3(new_n270), .A4(new_n280), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT95), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n289), .A2(new_n290), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n290), .B1(new_n289), .B2(new_n298), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n202), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT89), .B(G134gat), .ZN(new_n302));
  AND3_X1   g101(.A1(new_n282), .A2(KEYINPUT96), .A3(new_n284), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT96), .B1(new_n282), .B2(new_n284), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n295), .B(KEYINPUT95), .ZN(new_n306));
  OAI21_X1  g105(.A(G162gat), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n202), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n289), .A2(new_n290), .A3(new_n298), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n301), .A2(new_n302), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n302), .B1(new_n301), .B2(new_n310), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G71gat), .B(G78gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(G57gat), .A2(G64gat), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT87), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(G57gat), .A2(G64gat), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n318), .B(new_n319), .C1(new_n317), .C2(new_n316), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n314), .B1(new_n320), .B2(KEYINPUT86), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n320), .A2(KEYINPUT86), .A3(new_n314), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OR2_X1    g123(.A1(new_n324), .A2(KEYINPUT21), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(KEYINPUT21), .ZN(new_n326));
  XNOR2_X1  g125(.A(G15gat), .B(G22gat), .ZN(new_n327));
  OR2_X1    g126(.A1(new_n327), .A2(G1gat), .ZN(new_n328));
  INV_X1    g127(.A(G8gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT16), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n327), .B1(new_n330), .B2(G1gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n328), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n329), .B1(new_n328), .B2(new_n331), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n325), .A2(new_n326), .A3(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n336), .B1(new_n325), .B2(new_n335), .ZN(new_n337));
  XNOR2_X1  g136(.A(G127gat), .B(G155gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n337), .B(new_n338), .ZN(new_n339));
  AND2_X1   g138(.A1(G231gat), .A2(G233gat), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  OR2_X1    g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n339), .A2(new_n341), .ZN(new_n343));
  XNOR2_X1  g142(.A(G183gat), .B(G211gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n344), .B(KEYINPUT20), .ZN(new_n345));
  XNOR2_X1  g144(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n345), .B(new_n346), .ZN(new_n347));
  AND3_X1   g146(.A1(new_n342), .A2(new_n343), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n347), .B1(new_n342), .B2(new_n343), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G113gat), .B(G141gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n351), .B(G197gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(KEYINPUT11), .ZN(new_n353));
  INV_X1    g152(.A(G169gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n353), .B(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT12), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT84), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n358), .B1(new_n333), .B2(new_n334), .ZN(new_n359));
  INV_X1    g158(.A(new_n334), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(KEYINPUT84), .A3(new_n332), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n359), .A2(new_n361), .A3(new_n229), .A4(new_n234), .ZN(new_n362));
  NAND2_X1  g161(.A1(G229gat), .A2(G233gat), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n279), .B1(new_n334), .B2(new_n333), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT18), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT85), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n357), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n335), .B1(new_n226), .B2(new_n228), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n364), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n363), .B(KEYINPUT13), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n362), .A2(KEYINPUT18), .A3(new_n363), .A4(new_n364), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n367), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n369), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n376), .A2(new_n357), .A3(new_n368), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n254), .A2(new_n266), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n264), .A2(KEYINPUT97), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n324), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n323), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n383), .B1(new_n385), .B2(new_n321), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(new_n381), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT10), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  OAI211_X1 g187(.A(KEYINPUT10), .B(new_n324), .C1(new_n267), .C2(new_n268), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(G230gat), .ZN(new_n391));
  INV_X1    g190(.A(G233gat), .ZN(new_n392));
  OAI22_X1  g191(.A1(new_n388), .A2(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n391), .A2(new_n392), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n384), .A2(new_n387), .A3(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(G120gat), .B(G148gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n396), .B(KEYINPUT98), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(G176gat), .ZN(new_n398));
  XOR2_X1   g197(.A(new_n398), .B(G204gat), .Z(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n393), .A2(new_n395), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n400), .B1(new_n393), .B2(new_n395), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n380), .A2(new_n404), .ZN(new_n405));
  NOR3_X1   g204(.A1(new_n313), .A2(new_n350), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT25), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT24), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n408), .A2(G183gat), .A3(G190gat), .ZN(new_n409));
  NAND2_X1  g208(.A1(G169gat), .A2(G176gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(G183gat), .A2(G190gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT24), .ZN(new_n412));
  NOR2_X1   g211(.A1(G183gat), .A2(G190gat), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n409), .B(new_n410), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NOR3_X1   g215(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n407), .B1(new_n414), .B2(new_n418), .ZN(new_n419));
  OR3_X1    g218(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n415), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n409), .A2(new_n410), .ZN(new_n422));
  INV_X1    g221(.A(new_n413), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n423), .A2(KEYINPUT24), .A3(new_n411), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n421), .A2(new_n422), .A3(new_n424), .A4(KEYINPUT25), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n419), .A2(new_n425), .ZN(new_n426));
  AND2_X1   g225(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n427));
  NOR2_X1   g226(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n428));
  OR2_X1    g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT28), .ZN(new_n430));
  INV_X1    g229(.A(G190gat), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n431), .B1(new_n427), .B2(new_n428), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT28), .ZN(new_n434));
  OR3_X1    g233(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(new_n410), .A3(new_n436), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n432), .A2(new_n411), .A3(new_n434), .A4(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n426), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(G120gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(G113gat), .ZN(new_n441));
  INV_X1    g240(.A(G113gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(G120gat), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT1), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT64), .ZN(new_n445));
  INV_X1    g244(.A(G134gat), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n445), .A2(new_n446), .A3(G127gat), .ZN(new_n447));
  INV_X1    g246(.A(G127gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(G134gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT65), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT64), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n445), .A2(KEYINPUT65), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n447), .A2(new_n449), .A3(new_n452), .A4(new_n453), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n444), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(G127gat), .B(G134gat), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n444), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n439), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(G227gat), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n462), .A2(new_n392), .ZN(new_n463));
  INV_X1    g262(.A(new_n444), .ZN(new_n464));
  INV_X1    g263(.A(new_n456), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n449), .A2(new_n447), .B1(new_n452), .B2(new_n453), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n459), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n469), .A2(new_n426), .A3(new_n438), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n461), .A2(new_n463), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT33), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(G15gat), .B(G43gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(G71gat), .ZN(new_n475));
  INV_X1    g274(.A(G99gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n475), .B(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n473), .A2(KEYINPUT66), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n471), .A2(KEYINPUT32), .ZN(new_n479));
  INV_X1    g278(.A(new_n477), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT67), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n472), .B1(new_n480), .B2(new_n481), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n478), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n473), .A2(new_n477), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n479), .B1(new_n486), .B2(KEYINPUT66), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT34), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n461), .A2(new_n470), .ZN(new_n489));
  INV_X1    g288(.A(new_n463), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AOI211_X1 g290(.A(KEYINPUT34), .B(new_n463), .C1(new_n461), .C2(new_n470), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n485), .A2(new_n487), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n493), .B1(new_n485), .B2(new_n487), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(G155gat), .A2(G162gat), .ZN(new_n497));
  INV_X1    g296(.A(G155gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n290), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n497), .B1(new_n499), .B2(KEYINPUT2), .ZN(new_n500));
  INV_X1    g299(.A(G148gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(G141gat), .ZN(new_n502));
  INV_X1    g301(.A(G141gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(G148gat), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT72), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n502), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n505), .B1(new_n502), .B2(new_n504), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n500), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n502), .A2(new_n504), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT2), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n511), .A2(new_n497), .A3(new_n499), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT3), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n508), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT74), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT74), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n508), .A2(new_n512), .A3(new_n516), .A4(new_n513), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  XOR2_X1   g317(.A(KEYINPUT71), .B(KEYINPUT29), .Z(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G197gat), .B(G204gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT22), .ZN(new_n523));
  INV_X1    g322(.A(G211gat), .ZN(new_n524));
  INV_X1    g323(.A(G218gat), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n524), .A2(new_n525), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n523), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AND3_X1   g328(.A1(new_n524), .A2(new_n525), .A3(KEYINPUT22), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n522), .B1(new_n530), .B2(new_n526), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(KEYINPUT69), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT79), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n521), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n508), .A2(new_n512), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT73), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n508), .A2(new_n512), .A3(KEYINPUT73), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT29), .B1(new_n529), .B2(new_n531), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n541), .B1(KEYINPUT3), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n519), .B1(new_n515), .B2(new_n517), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT79), .B1(new_n544), .B2(new_n533), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n536), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(G228gat), .A2(G233gat), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT78), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n529), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n531), .A2(KEYINPUT77), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n531), .A2(KEYINPUT77), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n529), .A2(new_n550), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT3), .B1(new_n555), .B2(new_n520), .ZN(new_n556));
  AND2_X1   g355(.A1(G155gat), .A2(G162gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(G155gat), .A2(G162gat), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n557), .B1(new_n510), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n503), .A2(G148gat), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n501), .A2(G141gat), .ZN(new_n561));
  OAI21_X1  g360(.A(KEYINPUT72), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n502), .A2(new_n504), .A3(new_n505), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n559), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n499), .A2(new_n497), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n565), .B1(new_n510), .B2(new_n509), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  OAI221_X1 g366(.A(new_n547), .B1(new_n544), .B2(new_n533), .C1(new_n556), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n549), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G78gat), .B(G106gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G22gat), .ZN(new_n571));
  XOR2_X1   g370(.A(KEYINPUT31), .B(G50gat), .Z(new_n572));
  XOR2_X1   g371(.A(new_n571), .B(new_n572), .Z(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n549), .A2(new_n568), .A3(new_n573), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT81), .ZN(new_n578));
  NOR3_X1   g377(.A1(new_n496), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G8gat), .B(G36gat), .ZN(new_n580));
  INV_X1    g379(.A(G64gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(new_n256), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n439), .A2(KEYINPUT70), .ZN(new_n585));
  NAND2_X1  g384(.A1(G226gat), .A2(G233gat), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT70), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n426), .A2(new_n588), .A3(new_n438), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n585), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT29), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n439), .A2(new_n591), .A3(new_n586), .ZN(new_n592));
  AND3_X1   g391(.A1(new_n590), .A2(new_n533), .A3(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n519), .A2(new_n587), .ZN(new_n594));
  AND3_X1   g393(.A1(new_n426), .A2(new_n588), .A3(new_n438), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n588), .B1(new_n426), .B2(new_n438), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n439), .A2(new_n586), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n533), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n584), .B1(new_n593), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n590), .A2(new_n533), .A3(new_n592), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n589), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n598), .B1(new_n603), .B2(new_n594), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n602), .B(new_n583), .C1(new_n604), .C2(new_n533), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n601), .A2(KEYINPUT30), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT30), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n607), .B(new_n584), .C1(new_n593), .C2(new_n600), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT75), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n610), .B1(new_n469), .B2(new_n537), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n460), .A2(KEYINPUT75), .A3(new_n567), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n611), .A2(new_n612), .B1(new_n541), .B2(new_n469), .ZN(new_n613));
  NAND2_X1  g412(.A1(G225gat), .A2(G233gat), .ZN(new_n614));
  OAI21_X1  g413(.A(KEYINPUT76), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT4), .ZN(new_n616));
  NOR3_X1   g415(.A1(new_n469), .A2(new_n610), .A3(new_n537), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT75), .B1(new_n460), .B2(new_n567), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NOR3_X1   g418(.A1(new_n564), .A2(new_n538), .A3(new_n566), .ZN(new_n620));
  AOI21_X1  g419(.A(KEYINPUT73), .B1(new_n508), .B2(new_n512), .ZN(new_n621));
  OAI21_X1  g420(.A(KEYINPUT3), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n518), .A2(new_n622), .A3(new_n469), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n460), .A2(KEYINPUT4), .A3(new_n567), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n619), .A2(new_n623), .A3(new_n614), .A4(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n469), .B1(new_n620), .B2(new_n621), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n626), .B1(new_n617), .B2(new_n618), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT76), .ZN(new_n628));
  INV_X1    g427(.A(new_n614), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n615), .A2(new_n625), .A3(KEYINPUT5), .A4(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n611), .A2(KEYINPUT4), .A3(new_n612), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n616), .B1(new_n469), .B2(new_n537), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n623), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n629), .A2(KEYINPUT5), .ZN(new_n635));
  OR2_X1    g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G1gat), .B(G29gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT0), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(G57gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(new_n255), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT6), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n631), .A2(new_n641), .A3(new_n636), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n637), .A2(KEYINPUT6), .A3(new_n642), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n609), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n579), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT35), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n579), .A2(new_n648), .A3(KEYINPUT35), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT68), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT36), .ZN(new_n654));
  OAI211_X1 g453(.A(new_n653), .B(new_n654), .C1(new_n494), .C2(new_n495), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n485), .A2(new_n487), .ZN(new_n656));
  INV_X1    g455(.A(new_n493), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n485), .A2(new_n487), .A3(new_n493), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n653), .A2(new_n654), .ZN(new_n660));
  NAND2_X1  g459(.A1(KEYINPUT68), .A2(KEYINPUT36), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n658), .A2(new_n659), .A3(new_n660), .A4(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n655), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n645), .A2(new_n644), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n641), .B1(new_n631), .B2(new_n636), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT37), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n668), .B1(new_n593), .B2(new_n600), .ZN(new_n669));
  OAI211_X1 g468(.A(KEYINPUT37), .B(new_n602), .C1(new_n604), .C2(new_n533), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n669), .A2(new_n583), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(KEYINPUT38), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n604), .A2(new_n533), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n590), .A2(new_n592), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(new_n534), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n673), .A2(KEYINPUT37), .A3(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT38), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n676), .A2(new_n669), .A3(new_n677), .A4(new_n583), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n672), .A2(new_n601), .A3(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n647), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n667), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n577), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT40), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n614), .B(new_n626), .C1(new_n617), .C2(new_n618), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT39), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT80), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n634), .A2(new_n629), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n684), .A2(KEYINPUT80), .A3(KEYINPUT39), .ZN(new_n689));
  AND3_X1   g488(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT39), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n634), .A2(new_n691), .A3(new_n629), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n641), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n683), .B1(new_n690), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n609), .A2(new_n694), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n692), .A2(new_n641), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n696), .A2(KEYINPUT40), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n643), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n682), .B1(new_n695), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n664), .B1(new_n681), .B2(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n648), .A2(new_n682), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n651), .B(new_n652), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n406), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT99), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT99), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n406), .A2(new_n706), .A3(new_n703), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n646), .A2(new_n647), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(G1gat), .ZN(G1324gat));
  INV_X1    g511(.A(new_n708), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n606), .A2(new_n608), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n715), .A2(KEYINPUT100), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n708), .A2(KEYINPUT100), .A3(new_n609), .ZN(new_n717));
  OAI21_X1  g516(.A(G8gat), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(KEYINPUT16), .B(G8gat), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n715), .A2(KEYINPUT42), .A3(new_n720), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n716), .A2(new_n717), .A3(new_n719), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n718), .B(new_n721), .C1(new_n722), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g522(.A(new_n496), .ZN(new_n724));
  AOI21_X1  g523(.A(G15gat), .B1(new_n708), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n713), .A2(new_n664), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n725), .B1(new_n726), .B2(G15gat), .ZN(G1326gat));
  INV_X1    g526(.A(KEYINPUT101), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n728), .B1(new_n708), .B2(new_n577), .ZN(new_n729));
  AOI211_X1 g528(.A(KEYINPUT101), .B(new_n682), .C1(new_n705), .C2(new_n707), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT43), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT43), .B1(new_n729), .B2(new_n730), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n733), .A2(G22gat), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(G22gat), .B1(new_n733), .B2(new_n734), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n735), .A2(new_n736), .ZN(G1327gat));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n698), .A2(new_n643), .ZN(new_n739));
  AOI21_X1  g538(.A(KEYINPUT40), .B1(new_n696), .B2(new_n697), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n740), .A2(new_n714), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n577), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n678), .A2(new_n601), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n646), .A2(new_n743), .A3(new_n647), .A4(new_n672), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n663), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n709), .A2(new_n714), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n746), .A2(KEYINPUT104), .A3(new_n577), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT104), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n648), .B2(new_n682), .ZN(new_n749));
  AND3_X1   g548(.A1(new_n745), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n651), .A2(new_n652), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n738), .B(new_n313), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n738), .B1(new_n703), .B2(new_n313), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT105), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n745), .A2(new_n747), .A3(new_n749), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n756), .A2(new_n651), .A3(new_n652), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n757), .A2(KEYINPUT105), .A3(new_n738), .A4(new_n313), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n350), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n760), .A2(new_n405), .ZN(new_n761));
  XOR2_X1   g560(.A(new_n761), .B(KEYINPUT103), .Z(new_n762));
  AND2_X1   g561(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(G29gat), .B1(new_n764), .B2(new_n709), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n761), .A2(new_n703), .A3(new_n313), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n766), .A2(new_n203), .A3(new_n710), .ZN(new_n767));
  XOR2_X1   g566(.A(KEYINPUT102), .B(KEYINPUT45), .Z(new_n768));
  XNOR2_X1  g567(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n765), .A2(new_n769), .ZN(G1328gat));
  OAI21_X1  g569(.A(G36gat), .B1(new_n764), .B2(new_n714), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n766), .A2(new_n204), .A3(new_n609), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT46), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(KEYINPUT106), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n772), .A2(KEYINPUT46), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT107), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n771), .A2(new_n774), .A3(new_n776), .ZN(G1329gat));
  AOI21_X1  g576(.A(new_n231), .B1(new_n763), .B2(new_n663), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n724), .A2(new_n231), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n778), .B1(new_n766), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g580(.A(new_n216), .B1(new_n763), .B2(new_n577), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n682), .A2(G50gat), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n782), .B1(new_n766), .B2(new_n783), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g584(.A(new_n757), .ZN(new_n786));
  INV_X1    g585(.A(new_n302), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n308), .B1(new_n307), .B2(new_n309), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n301), .A2(new_n302), .A3(new_n310), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n350), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n404), .ZN(new_n793));
  INV_X1    g592(.A(new_n380), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT108), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n792), .A2(KEYINPUT108), .A3(new_n793), .A4(new_n794), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n786), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n710), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g600(.A1(new_n797), .A2(new_n798), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n757), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n803), .A2(new_n714), .ZN(new_n804));
  NOR2_X1   g603(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n805));
  AND2_X1   g604(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n807), .B1(new_n804), .B2(new_n805), .ZN(new_n808));
  XOR2_X1   g607(.A(new_n808), .B(KEYINPUT109), .Z(G1333gat));
  NAND3_X1  g608(.A1(new_n799), .A2(G71gat), .A3(new_n663), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT110), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT110), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n799), .A2(new_n812), .A3(G71gat), .A4(new_n663), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(G71gat), .B1(new_n799), .B2(new_n724), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT111), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT111), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n814), .A2(new_n819), .A3(new_n816), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n818), .A2(KEYINPUT50), .A3(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT50), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n819), .B1(new_n814), .B2(new_n816), .ZN(new_n823));
  AOI211_X1 g622(.A(KEYINPUT111), .B(new_n815), .C1(new_n811), .C2(new_n813), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n821), .A2(new_n825), .ZN(G1334gat));
  NAND2_X1  g625(.A1(new_n799), .A2(new_n577), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g627(.A1(new_n760), .A2(new_n380), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n793), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n759), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(G85gat), .B1(new_n832), .B2(new_n709), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n757), .A2(new_n313), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(KEYINPUT51), .A3(new_n829), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT51), .B1(new_n834), .B2(new_n829), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT112), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n838), .B1(KEYINPUT112), .B2(new_n837), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(new_n255), .A3(new_n710), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n833), .B1(new_n840), .B2(new_n404), .ZN(G1336gat));
  NOR3_X1   g640(.A1(new_n404), .A2(G92gat), .A3(new_n714), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n759), .A2(new_n609), .A3(new_n831), .ZN(new_n844));
  AOI21_X1  g643(.A(KEYINPUT52), .B1(new_n844), .B2(G92gat), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT113), .ZN(new_n847));
  AOI211_X1 g646(.A(new_n714), .B(new_n830), .C1(new_n755), .C2(new_n758), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n847), .B1(new_n848), .B2(new_n256), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n829), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n835), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n842), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n844), .A2(KEYINPUT113), .A3(G92gat), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n849), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT114), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n856), .A2(new_n857), .A3(KEYINPUT52), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n857), .B1(new_n856), .B2(KEYINPUT52), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n846), .B1(new_n858), .B2(new_n859), .ZN(G1337gat));
  OAI21_X1  g659(.A(G99gat), .B1(new_n832), .B2(new_n664), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n839), .A2(new_n476), .A3(new_n793), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n861), .B1(new_n862), .B2(new_n496), .ZN(G1338gat));
  OAI21_X1  g662(.A(G106gat), .B1(new_n832), .B2(new_n682), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT53), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n682), .A2(new_n404), .A3(G106gat), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n867), .B1(new_n839), .B2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT112), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n870), .B1(new_n852), .B2(new_n835), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n837), .A2(KEYINPUT112), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n867), .B(new_n868), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n866), .B1(new_n869), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n853), .A2(new_n868), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n865), .B1(new_n864), .B2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT115), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n877), .A2(new_n878), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n875), .B1(new_n879), .B2(new_n880), .ZN(G1339gat));
  OR2_X1    g680(.A1(new_n376), .A2(new_n357), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n399), .B1(new_n393), .B2(KEYINPUT54), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n384), .A2(new_n387), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT10), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n394), .A3(new_n389), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(new_n393), .A3(KEYINPUT54), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n884), .A2(KEYINPUT55), .A3(new_n889), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n890), .A2(new_n401), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n363), .B1(new_n362), .B2(new_n364), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n370), .A2(new_n364), .A3(new_n372), .ZN(new_n893));
  AOI22_X1  g692(.A1(new_n892), .A2(KEYINPUT117), .B1(KEYINPUT118), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n894), .B1(KEYINPUT117), .B2(new_n892), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n893), .A2(KEYINPUT118), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n355), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT55), .ZN(new_n898));
  AND3_X1   g697(.A1(new_n888), .A2(new_n393), .A3(KEYINPUT54), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n898), .B1(new_n899), .B2(new_n883), .ZN(new_n900));
  AND4_X1   g699(.A1(new_n882), .A2(new_n891), .A3(new_n897), .A4(new_n900), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n790), .A2(new_n901), .A3(new_n791), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n793), .A2(new_n882), .A3(new_n897), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n891), .A2(new_n380), .A3(new_n900), .ZN(new_n904));
  AOI22_X1  g703(.A1(new_n790), .A2(new_n791), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n350), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n792), .A2(new_n404), .A3(new_n794), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n496), .A2(new_n577), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n710), .A3(new_n714), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n911), .A2(new_n794), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(new_n442), .ZN(G1340gat));
  NOR2_X1   g712(.A1(new_n911), .A2(new_n404), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(new_n440), .ZN(G1341gat));
  NOR2_X1   g714(.A1(new_n911), .A2(new_n350), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(new_n448), .ZN(G1342gat));
  NAND2_X1  g716(.A1(new_n790), .A2(new_n791), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n911), .A2(new_n918), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n919), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n920));
  XOR2_X1   g719(.A(KEYINPUT56), .B(G134gat), .Z(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n919), .B2(new_n921), .ZN(G1343gat));
  INV_X1    g721(.A(KEYINPUT120), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n900), .A2(new_n923), .ZN(new_n924));
  OAI211_X1 g723(.A(KEYINPUT120), .B(new_n898), .C1(new_n899), .C2(new_n883), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n891), .A2(new_n380), .A3(new_n924), .A4(new_n925), .ZN(new_n926));
  AOI22_X1  g725(.A1(new_n790), .A2(new_n791), .B1(new_n903), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n350), .B1(new_n902), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n682), .B1(new_n928), .B2(new_n907), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT57), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n908), .A2(new_n930), .A3(new_n577), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n663), .A2(new_n709), .A3(new_n609), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT119), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n931), .A2(new_n380), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n908), .A2(new_n577), .A3(new_n933), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n794), .A2(G141gat), .ZN(new_n937));
  AOI22_X1  g736(.A1(new_n935), .A2(G141gat), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OR2_X1    g737(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n939));
  NAND2_X1  g738(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n939), .B1(new_n938), .B2(new_n940), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n941), .A2(new_n942), .ZN(G1344gat));
  INV_X1    g742(.A(KEYINPUT59), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n931), .A2(new_n932), .A3(new_n934), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n945), .B2(new_n404), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n908), .A2(KEYINPUT57), .A3(new_n577), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n947), .B1(KEYINPUT57), .B2(new_n929), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n948), .A2(KEYINPUT59), .A3(new_n793), .A4(new_n934), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n501), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(G148gat), .B1(new_n936), .B2(new_n793), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n950), .B1(KEYINPUT59), .B2(new_n951), .ZN(G1345gat));
  NOR3_X1   g751(.A1(new_n945), .A2(new_n498), .A3(new_n350), .ZN(new_n953));
  AOI21_X1  g752(.A(G155gat), .B1(new_n936), .B2(new_n760), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n953), .A2(new_n954), .ZN(G1346gat));
  NOR3_X1   g754(.A1(new_n945), .A2(new_n290), .A3(new_n918), .ZN(new_n956));
  AOI21_X1  g755(.A(G162gat), .B1(new_n936), .B2(new_n313), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n956), .A2(new_n957), .ZN(G1347gat));
  AOI21_X1  g757(.A(KEYINPUT122), .B1(new_n908), .B2(new_n709), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT122), .ZN(new_n960));
  AOI211_X1 g759(.A(new_n960), .B(new_n710), .C1(new_n906), .C2(new_n907), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n909), .A2(new_n609), .ZN(new_n963));
  XOR2_X1   g762(.A(new_n963), .B(KEYINPUT123), .Z(new_n964));
  AND2_X1   g763(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n965), .A2(new_n354), .A3(new_n380), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n710), .A2(new_n714), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n910), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(G169gat), .B1(new_n968), .B2(new_n794), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n966), .A2(new_n969), .ZN(G1348gat));
  INV_X1    g769(.A(G176gat), .ZN(new_n971));
  NOR3_X1   g770(.A1(new_n968), .A2(new_n971), .A3(new_n404), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n965), .A2(new_n793), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n972), .B1(new_n973), .B2(new_n971), .ZN(G1349gat));
  NAND4_X1  g773(.A1(new_n962), .A2(new_n429), .A3(new_n760), .A4(new_n964), .ZN(new_n975));
  OAI21_X1  g774(.A(G183gat), .B1(new_n968), .B2(new_n350), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n977), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g777(.A1(new_n910), .A2(new_n313), .A3(new_n967), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT61), .ZN(new_n980));
  AND3_X1   g779(.A1(new_n979), .A2(new_n980), .A3(G190gat), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n980), .B1(new_n979), .B2(G190gat), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n962), .A2(new_n431), .A3(new_n964), .ZN(new_n983));
  OAI22_X1  g782(.A1(new_n981), .A2(new_n982), .B1(new_n918), .B2(new_n983), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT124), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI221_X1 g785(.A(KEYINPUT124), .B1(new_n983), .B2(new_n918), .C1(new_n981), .C2(new_n982), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n986), .A2(new_n987), .ZN(G1351gat));
  NOR3_X1   g787(.A1(new_n663), .A2(new_n714), .A3(new_n682), .ZN(new_n989));
  AND2_X1   g788(.A1(new_n962), .A2(new_n989), .ZN(new_n990));
  INV_X1    g789(.A(G197gat), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n990), .A2(new_n991), .A3(new_n380), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n967), .A2(new_n664), .ZN(new_n993));
  INV_X1    g792(.A(new_n993), .ZN(new_n994));
  AND2_X1   g793(.A1(new_n948), .A2(new_n994), .ZN(new_n995));
  AND2_X1   g794(.A1(new_n995), .A2(new_n380), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n992), .B1(new_n996), .B2(new_n991), .ZN(G1352gat));
  INV_X1    g796(.A(KEYINPUT126), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n908), .A2(new_n709), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n999), .A2(new_n960), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n908), .A2(KEYINPUT122), .A3(new_n709), .ZN(new_n1001));
  NOR2_X1   g800(.A1(new_n404), .A2(G204gat), .ZN(new_n1002));
  NAND4_X1  g801(.A1(new_n1000), .A2(new_n1001), .A3(new_n989), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1003), .A2(KEYINPUT125), .ZN(new_n1004));
  INV_X1    g803(.A(KEYINPUT125), .ZN(new_n1005));
  NAND4_X1  g804(.A1(new_n962), .A2(new_n1005), .A3(new_n989), .A4(new_n1002), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n998), .B1(new_n1007), .B2(KEYINPUT62), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1007), .A2(KEYINPUT62), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n948), .A2(new_n793), .A3(new_n994), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1010), .A2(G204gat), .ZN(new_n1011));
  INV_X1    g810(.A(KEYINPUT62), .ZN(new_n1012));
  NAND4_X1  g811(.A1(new_n1004), .A2(new_n1006), .A3(KEYINPUT126), .A4(new_n1012), .ZN(new_n1013));
  NAND4_X1  g812(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .A4(new_n1013), .ZN(G1353gat));
  NAND2_X1  g813(.A1(new_n928), .A2(new_n907), .ZN(new_n1015));
  AOI21_X1  g814(.A(KEYINPUT57), .B1(new_n1015), .B2(new_n577), .ZN(new_n1016));
  AOI211_X1 g815(.A(new_n930), .B(new_n682), .C1(new_n906), .C2(new_n907), .ZN(new_n1017));
  OAI211_X1 g816(.A(new_n760), .B(new_n994), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  INV_X1    g817(.A(KEYINPUT127), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g819(.A1(new_n948), .A2(KEYINPUT127), .A3(new_n760), .A4(new_n994), .ZN(new_n1021));
  NAND3_X1  g820(.A1(new_n1020), .A2(G211gat), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g821(.A(KEYINPUT63), .ZN(new_n1023));
  NAND2_X1  g822(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND4_X1  g823(.A1(new_n1020), .A2(new_n1021), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n1025));
  NAND2_X1  g824(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g825(.A1(new_n990), .A2(new_n524), .A3(new_n760), .ZN(new_n1027));
  NAND2_X1  g826(.A1(new_n1026), .A2(new_n1027), .ZN(G1354gat));
  AOI21_X1  g827(.A(G218gat), .B1(new_n990), .B2(new_n313), .ZN(new_n1029));
  NOR2_X1   g828(.A1(new_n918), .A2(new_n525), .ZN(new_n1030));
  AOI21_X1  g829(.A(new_n1029), .B1(new_n995), .B2(new_n1030), .ZN(G1355gat));
endmodule


