//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 1 0 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005;
  XNOR2_X1  g000(.A(G110), .B(G122), .ZN(new_n187));
  XOR2_X1   g001(.A(new_n187), .B(KEYINPUT83), .Z(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  NOR3_X1   g003(.A1(new_n189), .A2(KEYINPUT3), .A3(G107), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G104), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT77), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n194), .B(KEYINPUT3), .C1(new_n189), .C2(G107), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n191), .A2(G104), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n194), .B1(new_n197), .B2(KEYINPUT3), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n193), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G101), .ZN(new_n200));
  INV_X1    g014(.A(G101), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n193), .B(new_n201), .C1(new_n196), .C2(new_n198), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n200), .A2(KEYINPUT4), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G119), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT66), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT66), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G119), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n207), .A3(G116), .ZN(new_n208));
  OR2_X1    g022(.A1(new_n204), .A2(G116), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT2), .B(G113), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(KEYINPUT67), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n211), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT67), .ZN(new_n214));
  INV_X1    g028(.A(new_n211), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(new_n208), .A3(new_n209), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n213), .A2(new_n214), .A3(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT4), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n199), .A2(new_n218), .A3(G101), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n203), .A2(new_n212), .A3(new_n217), .A4(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n210), .A2(new_n211), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n208), .A2(KEYINPUT5), .ZN(new_n222));
  INV_X1    g036(.A(G113), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n208), .A2(KEYINPUT5), .A3(new_n209), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n221), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n189), .A2(G107), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n201), .B1(new_n197), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n202), .A2(KEYINPUT80), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(KEYINPUT80), .B1(new_n202), .B2(new_n229), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n226), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n188), .B1(new_n220), .B2(new_n232), .ZN(new_n233));
  OR2_X1    g047(.A1(new_n233), .A2(KEYINPUT6), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n220), .A2(new_n232), .A3(new_n188), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT84), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n220), .A2(new_n232), .A3(KEYINPUT84), .A4(new_n188), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n233), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT6), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n234), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G143), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n242), .A2(G146), .ZN(new_n243));
  INV_X1    g057(.A(G146), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT64), .B1(new_n244), .B2(G143), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT64), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n246), .A2(new_n242), .A3(G146), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n243), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  AND2_X1   g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  NOR2_X1   g063(.A1(KEYINPUT0), .A2(G128), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n244), .A2(G143), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n242), .A2(G146), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI22_X1  g068(.A1(new_n248), .A2(new_n249), .B1(new_n251), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G125), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n257), .B(KEYINPUT85), .ZN(new_n258));
  INV_X1    g072(.A(G128), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(KEYINPUT1), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n248), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(KEYINPUT1), .B1(new_n242), .B2(G146), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT65), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n252), .A2(KEYINPUT65), .A3(KEYINPUT1), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n259), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n254), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n261), .B(new_n256), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n268), .B(KEYINPUT86), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n258), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G224), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n271), .A2(G953), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n270), .B(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n241), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT7), .B1(new_n271), .B2(G953), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n258), .A2(new_n269), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT89), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n258), .A2(new_n269), .A3(KEYINPUT89), .A4(new_n276), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT88), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n269), .A2(new_n281), .ZN(new_n282));
  OR2_X1    g096(.A1(new_n268), .A2(KEYINPUT86), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n268), .A2(KEYINPUT86), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n283), .A2(KEYINPUT88), .A3(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n282), .A2(new_n258), .A3(new_n285), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n279), .A2(new_n280), .B1(new_n286), .B2(new_n275), .ZN(new_n287));
  XOR2_X1   g101(.A(new_n188), .B(KEYINPUT8), .Z(new_n288));
  NAND2_X1  g102(.A1(new_n202), .A2(new_n229), .ZN(new_n289));
  OR2_X1    g103(.A1(new_n225), .A2(KEYINPUT87), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n225), .A2(KEYINPUT87), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(new_n224), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n289), .B1(new_n292), .B2(new_n216), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n226), .A2(new_n289), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n288), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n295), .B1(new_n237), .B2(new_n238), .ZN(new_n296));
  AOI21_X1  g110(.A(G902), .B1(new_n287), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n274), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(G210), .B1(G237), .B2(G902), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n274), .A2(new_n297), .A3(new_n299), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(G214), .B1(G237), .B2(G902), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT90), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n274), .A2(new_n299), .A3(new_n297), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n299), .B1(new_n274), .B2(new_n297), .ZN(new_n307));
  OAI211_X1 g121(.A(KEYINPUT90), .B(new_n304), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT69), .B(G953), .ZN(new_n310));
  INV_X1    g124(.A(G237), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(G214), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n242), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n310), .A2(G143), .A3(G214), .A4(new_n311), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AND2_X1   g129(.A1(KEYINPUT18), .A2(G131), .ZN(new_n316));
  OR2_X1    g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G131), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n318), .B1(new_n313), .B2(new_n314), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT18), .ZN(new_n320));
  XNOR2_X1  g134(.A(G125), .B(G140), .ZN(new_n321));
  OR2_X1    g135(.A1(new_n321), .A2(KEYINPUT72), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(KEYINPUT72), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(new_n323), .A3(new_n244), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n321), .B(KEYINPUT91), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n324), .B1(new_n325), .B2(new_n244), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n317), .A2(new_n320), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT92), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n317), .A2(new_n320), .A3(KEYINPUT92), .A4(new_n326), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n315), .A2(G131), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n313), .A2(new_n318), .A3(new_n314), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT93), .B1(new_n334), .B2(KEYINPUT17), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT93), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT17), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n332), .A2(new_n336), .A3(new_n337), .A4(new_n333), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n321), .A2(KEYINPUT16), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT16), .ZN(new_n340));
  INV_X1    g154(.A(G140), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n341), .A3(G125), .ZN(new_n342));
  AOI21_X1  g156(.A(G146), .B1(new_n339), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n339), .A2(G146), .A3(new_n342), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  AOI211_X1 g159(.A(new_n343), .B(new_n345), .C1(new_n319), .C2(KEYINPUT17), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n335), .A2(new_n338), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n331), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(G113), .B(G122), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n349), .B(new_n189), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n322), .A2(new_n323), .ZN(new_n352));
  MUX2_X1   g166(.A(new_n352), .B(new_n325), .S(KEYINPUT19), .Z(new_n353));
  AOI21_X1  g167(.A(new_n345), .B1(new_n353), .B2(new_n244), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n350), .B1(new_n354), .B2(new_n334), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n331), .A2(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(G475), .A2(G902), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n351), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT20), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n348), .A2(new_n350), .B1(new_n331), .B2(new_n355), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT20), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(new_n361), .A3(new_n357), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n350), .A2(KEYINPUT95), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n348), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G902), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n331), .A2(new_n347), .A3(new_n363), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  XOR2_X1   g182(.A(KEYINPUT94), .B(G475), .Z(new_n369));
  AOI22_X1  g183(.A1(new_n359), .A2(new_n362), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G952), .ZN(new_n371));
  AOI211_X1 g185(.A(G953), .B(new_n371), .C1(G234), .C2(G237), .ZN(new_n372));
  AOI211_X1 g186(.A(new_n366), .B(new_n310), .C1(G234), .C2(G237), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT21), .B(G898), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G122), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G116), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n191), .B1(new_n378), .B2(KEYINPUT14), .ZN(new_n379));
  XNOR2_X1  g193(.A(G116), .B(G122), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n379), .B(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n242), .A2(G128), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n259), .A2(G143), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT96), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n382), .A2(new_n383), .A3(KEYINPUT96), .ZN(new_n386));
  AOI21_X1  g200(.A(G134), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n386), .ZN(new_n388));
  INV_X1    g202(.A(G134), .ZN(new_n389));
  NOR3_X1   g203(.A1(new_n388), .A2(new_n389), .A3(new_n384), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n381), .B1(new_n387), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n389), .B1(new_n388), .B2(new_n384), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n380), .B(new_n191), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT13), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n382), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n383), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n382), .A2(new_n394), .ZN(new_n397));
  OAI21_X1  g211(.A(G134), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n392), .A2(new_n393), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n391), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(KEYINPUT9), .B(G234), .ZN(new_n401));
  INV_X1    g215(.A(G217), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n401), .A2(new_n402), .A3(G953), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n403), .B(KEYINPUT97), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n400), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n391), .A2(new_n404), .A3(new_n399), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n366), .ZN(new_n409));
  INV_X1    g223(.A(G478), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n410), .A2(KEYINPUT15), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n411), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n413), .B1(new_n408), .B2(new_n366), .ZN(new_n414));
  OR3_X1    g228(.A1(new_n412), .A2(KEYINPUT98), .A3(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(KEYINPUT98), .B1(new_n412), .B2(new_n414), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n370), .A2(new_n376), .A3(new_n417), .ZN(new_n418));
  NOR3_X1   g232(.A1(new_n305), .A2(new_n309), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G469), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT11), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n421), .B1(new_n389), .B2(G137), .ZN(new_n422));
  INV_X1    g236(.A(G137), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n423), .A2(KEYINPUT11), .A3(G134), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n389), .A2(G137), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n422), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G131), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n422), .A2(new_n424), .A3(new_n318), .A4(new_n425), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n227), .B1(new_n197), .B2(KEYINPUT3), .ZN(new_n430));
  OAI21_X1  g244(.A(KEYINPUT3), .B1(new_n189), .B2(G107), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT77), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n430), .B1(new_n195), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n228), .B1(new_n433), .B2(new_n201), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n262), .A2(KEYINPUT79), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT79), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n252), .A2(new_n436), .A3(KEYINPUT1), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n259), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n261), .B1(new_n438), .B2(new_n248), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n261), .B1(new_n266), .B2(new_n267), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n434), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n429), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT12), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI211_X1 g259(.A(KEYINPUT12), .B(new_n429), .C1(new_n440), .C2(new_n442), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n202), .A2(KEYINPUT4), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n432), .A2(new_n195), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n201), .B1(new_n449), .B2(new_n193), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n219), .A2(new_n255), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT78), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT78), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n203), .A2(new_n454), .A3(new_n255), .A4(new_n219), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT80), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n289), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n202), .A2(KEYINPUT80), .A3(new_n229), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n441), .A2(KEYINPUT10), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT10), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n434), .A2(new_n439), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n460), .A2(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n429), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n456), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n447), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n310), .A2(G227), .ZN(new_n468));
  XNOR2_X1  g282(.A(G110), .B(G140), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n468), .B(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n456), .A2(new_n464), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n429), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(new_n466), .A3(new_n470), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n420), .B1(new_n476), .B2(new_n366), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n470), .B1(new_n474), .B2(new_n466), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n447), .A2(new_n466), .A3(new_n470), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n420), .B(new_n366), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT81), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n456), .A2(new_n464), .A3(new_n465), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n465), .B1(new_n456), .B2(new_n464), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n471), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n447), .A2(new_n466), .A3(new_n470), .ZN(new_n487));
  AOI21_X1  g301(.A(G902), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(KEYINPUT81), .B1(new_n488), .B2(new_n420), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n478), .B1(new_n483), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(G221), .B1(new_n401), .B2(G902), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(KEYINPUT82), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT82), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n481), .A2(new_n482), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n488), .A2(KEYINPUT81), .A3(new_n420), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n477), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n491), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n493), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n492), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  XNOR2_X1  g314(.A(KEYINPUT66), .B(G119), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n259), .A2(KEYINPUT23), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n259), .A2(KEYINPUT23), .A3(G119), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n504), .B1(KEYINPUT23), .B2(new_n259), .ZN(new_n505));
  NOR3_X1   g319(.A1(new_n503), .A2(G110), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n204), .A2(new_n259), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n507), .B1(new_n501), .B2(new_n259), .ZN(new_n508));
  XOR2_X1   g322(.A(KEYINPUT24), .B(G110), .Z(new_n509));
  NOR2_X1   g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n344), .B(new_n324), .C1(new_n506), .C2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(G110), .B1(new_n503), .B2(new_n505), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n508), .A2(new_n509), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n512), .B(new_n513), .C1(new_n345), .C2(new_n343), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n310), .A2(G221), .A3(G234), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT22), .B(G137), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n515), .B(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n511), .A2(new_n514), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT74), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT74), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n511), .A2(new_n514), .A3(new_n520), .A4(new_n517), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n511), .A2(new_n514), .ZN(new_n523));
  INV_X1    g337(.A(new_n517), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT73), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n517), .B1(new_n511), .B2(new_n514), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT73), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n522), .A2(new_n527), .A3(new_n366), .A4(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(KEYINPUT75), .A2(KEYINPUT25), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n528), .B(new_n526), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n534), .A2(new_n366), .A3(new_n522), .A4(new_n531), .ZN(new_n535));
  AOI22_X1  g349(.A1(new_n533), .A2(new_n535), .B1(KEYINPUT75), .B2(KEYINPUT25), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n402), .B1(G234), .B2(new_n366), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n534), .A2(new_n522), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n538), .A2(G902), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(KEYINPUT76), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n217), .A2(new_n212), .ZN(new_n545));
  INV_X1    g359(.A(new_n425), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n389), .A2(G137), .ZN(new_n547));
  OAI21_X1  g361(.A(G131), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AND2_X1   g362(.A1(new_n548), .A2(new_n428), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n441), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n429), .A2(new_n255), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AND2_X1   g366(.A1(KEYINPUT68), .A2(KEYINPUT30), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n441), .A2(new_n549), .B1(new_n429), .B2(new_n255), .ZN(new_n555));
  NOR2_X1   g369(.A1(KEYINPUT68), .A2(KEYINPUT30), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n545), .B1(new_n554), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n310), .A2(G210), .A3(new_n311), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(KEYINPUT27), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT26), .B(G101), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n561), .B(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n217), .A2(new_n212), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n552), .A2(new_n565), .ZN(new_n566));
  NOR4_X1   g380(.A1(new_n559), .A2(new_n564), .A3(KEYINPUT70), .A4(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT31), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n552), .A2(new_n565), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n555), .A2(new_n545), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT28), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n572), .B1(KEYINPUT28), .B2(new_n566), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n567), .A2(new_n568), .B1(new_n573), .B2(new_n564), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n554), .A2(new_n558), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n565), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT70), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n576), .A2(new_n577), .A3(new_n570), .A4(new_n563), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT31), .ZN(new_n579));
  AOI21_X1  g393(.A(G902), .B1(new_n574), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT32), .ZN(new_n581));
  INV_X1    g395(.A(G472), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n573), .A2(new_n564), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n559), .A2(new_n566), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n585), .A2(new_n577), .A3(new_n568), .A4(new_n563), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n579), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n587), .A2(new_n582), .A3(new_n366), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(KEYINPUT32), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n583), .A2(new_n589), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n572), .B(new_n563), .C1(KEYINPUT28), .C2(new_n566), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT29), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n366), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(KEYINPUT71), .ZN(new_n594));
  INV_X1    g408(.A(new_n585), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n564), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n596), .A2(new_n592), .A3(new_n591), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n593), .A2(KEYINPUT71), .ZN(new_n599));
  OAI21_X1  g413(.A(G472), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n544), .B1(new_n590), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n419), .A2(new_n500), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(G101), .ZN(G3));
  NAND2_X1  g417(.A1(new_n587), .A2(new_n366), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(G472), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n588), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n606), .A2(new_n544), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n492), .A2(new_n498), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n368), .A2(new_n369), .ZN(new_n609));
  AND4_X1   g423(.A1(new_n361), .A2(new_n351), .A3(new_n356), .A4(new_n357), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n361), .B1(new_n360), .B2(new_n357), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n409), .A2(new_n410), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n408), .A2(KEYINPUT33), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT100), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n400), .A2(KEYINPUT99), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT99), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n391), .A2(new_n617), .A3(new_n399), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n615), .B1(new_n619), .B2(new_n404), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n404), .B1(new_n616), .B2(new_n618), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(KEYINPUT100), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n620), .A2(new_n407), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n614), .B1(new_n623), .B2(KEYINPUT33), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n410), .A2(G902), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n613), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n612), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n304), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n630), .B1(new_n301), .B2(new_n302), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n376), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n608), .A2(new_n629), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(new_n634), .B(KEYINPUT101), .Z(new_n635));
  XOR2_X1   g449(.A(KEYINPUT34), .B(G104), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G6));
  NAND2_X1  g451(.A1(new_n359), .A2(new_n362), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n638), .A2(new_n609), .A3(new_n416), .A4(new_n415), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n632), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n608), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT35), .B(G107), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G9));
  NOR2_X1   g457(.A1(new_n524), .A2(KEYINPUT36), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n523), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n542), .ZN(new_n646));
  INV_X1    g460(.A(new_n538), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n646), .B1(new_n536), .B2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n606), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n419), .A2(new_n500), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT102), .ZN(new_n652));
  XNOR2_X1  g466(.A(KEYINPUT37), .B(G110), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G12));
  OAI21_X1  g468(.A(new_n304), .B1(new_n306), .B2(new_n307), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n499), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n590), .A2(new_n600), .ZN(new_n657));
  INV_X1    g471(.A(G900), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n372), .B1(new_n373), .B2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n639), .A2(new_n659), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n657), .A2(new_n648), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G128), .ZN(G30));
  XOR2_X1   g477(.A(new_n659), .B(KEYINPUT39), .Z(new_n664));
  NAND2_X1  g478(.A1(new_n500), .A2(new_n664), .ZN(new_n665));
  OR2_X1    g479(.A1(new_n665), .A2(KEYINPUT40), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(KEYINPUT40), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n303), .A2(KEYINPUT38), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n303), .A2(KEYINPUT38), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(G472), .A2(G902), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n595), .A2(new_n564), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n571), .A2(new_n564), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(G472), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n671), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT103), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n590), .A2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n417), .B1(new_n638), .B2(new_n609), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n679), .A2(new_n304), .A3(new_n649), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n666), .A2(new_n667), .A3(new_n670), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G143), .ZN(G45));
  INV_X1    g497(.A(new_n659), .ZN(new_n684));
  AND4_X1   g498(.A1(new_n612), .A2(new_n648), .A3(new_n627), .A4(new_n684), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n657), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n656), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G146), .ZN(G48));
  NOR2_X1   g502(.A1(new_n488), .A2(new_n420), .ZN(new_n689));
  AOI211_X1 g503(.A(new_n497), .B(new_n689), .C1(new_n494), .C2(new_n495), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n633), .A2(new_n601), .A3(new_n629), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT41), .B(G113), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G15));
  NAND3_X1  g507(.A1(new_n640), .A2(new_n601), .A3(new_n690), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G116), .ZN(G18));
  AOI21_X1  g509(.A(new_n689), .B1(new_n494), .B2(new_n495), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n491), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n697), .A2(new_n655), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n418), .A2(new_n649), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n698), .A2(new_n657), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G119), .ZN(G21));
  AOI22_X1  g515(.A1(new_n537), .A2(new_n538), .B1(new_n542), .B2(new_n540), .ZN(new_n702));
  AOI21_X1  g516(.A(KEYINPUT104), .B1(new_n604), .B2(G472), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT104), .ZN(new_n704));
  AOI211_X1 g518(.A(new_n704), .B(new_n582), .C1(new_n587), .C2(new_n366), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n702), .B(new_n588), .C1(new_n703), .C2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n697), .A2(new_n375), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n303), .A2(new_n304), .A3(new_n679), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n707), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G122), .ZN(G24));
  OAI21_X1  g526(.A(new_n704), .B1(new_n580), .B2(new_n582), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n604), .A2(KEYINPUT104), .A3(G472), .ZN(new_n714));
  AOI22_X1  g528(.A1(new_n713), .A2(new_n714), .B1(new_n582), .B2(new_n580), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n715), .A2(new_n690), .A3(new_n685), .A4(new_n631), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT105), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n698), .A2(KEYINPUT105), .A3(new_n685), .A4(new_n715), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G125), .ZN(G27));
  NAND3_X1  g535(.A1(new_n301), .A2(new_n304), .A3(new_n302), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n722), .A2(new_n496), .A3(new_n497), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n628), .A2(new_n659), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n723), .A2(new_n601), .A3(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT42), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n723), .A2(new_n601), .A3(KEYINPUT42), .A4(new_n724), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G131), .ZN(G33));
  NAND3_X1  g544(.A1(new_n723), .A2(new_n601), .A3(new_n660), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G134), .ZN(G36));
  AND2_X1   g546(.A1(new_n472), .A2(new_n475), .ZN(new_n733));
  OAI21_X1  g547(.A(G469), .B1(new_n733), .B2(KEYINPUT45), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT106), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n736), .B(G469), .C1(new_n733), .C2(KEYINPUT45), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n733), .A2(KEYINPUT45), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n735), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(G469), .A2(G902), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT46), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n494), .A2(new_n495), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n739), .A2(KEYINPUT46), .A3(new_n740), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(new_n491), .A3(new_n664), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n722), .B(KEYINPUT107), .ZN(new_n748));
  INV_X1    g562(.A(new_n622), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n407), .B1(new_n621), .B2(KEYINPUT100), .ZN(new_n750));
  OAI21_X1  g564(.A(KEYINPUT33), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(KEYINPUT33), .B2(new_n408), .ZN(new_n752));
  AOI22_X1  g566(.A1(new_n752), .A2(new_n625), .B1(new_n410), .B2(new_n409), .ZN(new_n753));
  OAI21_X1  g567(.A(KEYINPUT43), .B1(new_n753), .B2(new_n612), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT43), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n370), .A2(new_n755), .A3(new_n627), .ZN(new_n756));
  AND4_X1   g570(.A1(new_n606), .A2(new_n754), .A3(new_n648), .A4(new_n756), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n757), .A2(KEYINPUT44), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n757), .A2(KEYINPUT44), .ZN(new_n759));
  NOR4_X1   g573(.A1(new_n747), .A2(new_n748), .A3(new_n758), .A4(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(new_n423), .ZN(G39));
  NAND2_X1  g575(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n745), .A2(new_n744), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT46), .B1(new_n739), .B2(new_n740), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n491), .B(new_n762), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(new_n766), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n746), .A2(new_n491), .A3(new_n762), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n722), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n724), .A2(new_n771), .A3(new_n544), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n657), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G140), .ZN(G42));
  NOR2_X1   g589(.A1(G952), .A2(G953), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n691), .A2(new_n711), .A3(new_n700), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n778), .A2(new_n729), .A3(new_n694), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n500), .B(new_n631), .C1(new_n661), .C2(new_n686), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n659), .B(KEYINPUT114), .ZN(new_n781));
  NOR4_X1   g595(.A1(new_n496), .A2(new_n497), .A3(new_n648), .A4(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n710), .A2(new_n782), .A3(new_n677), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n780), .A2(new_n720), .A3(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n780), .A2(new_n720), .A3(KEYINPUT52), .A4(new_n783), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n779), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT109), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT90), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n655), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n791), .A2(new_n376), .A3(new_n308), .A4(new_n629), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n608), .B1(new_n789), .B2(new_n792), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n792), .A2(new_n789), .ZN(new_n794));
  OAI211_X1 g608(.A(KEYINPUT110), .B(new_n602), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n305), .A2(new_n309), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n797), .A2(KEYINPUT109), .A3(new_n376), .A4(new_n629), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n792), .A2(new_n789), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n608), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT110), .B1(new_n800), .B2(new_n602), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n796), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n412), .A2(new_n414), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n612), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n791), .A2(new_n376), .A3(new_n308), .A4(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n608), .B1(KEYINPUT111), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n805), .A2(KEYINPUT111), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n651), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(KEYINPUT112), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT112), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n810), .B(new_n651), .C1(new_n806), .C2(new_n807), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  AND4_X1   g626(.A1(new_n370), .A2(new_n648), .A3(new_n803), .A4(new_n684), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n657), .A2(new_n771), .A3(new_n813), .ZN(new_n814));
  OR3_X1    g628(.A1(new_n814), .A2(new_n499), .A3(KEYINPUT113), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT113), .B1(new_n814), .B2(new_n499), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n715), .A2(new_n648), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(new_n724), .A3(new_n723), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n817), .A2(new_n731), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n788), .A2(new_n802), .A3(new_n812), .A4(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n811), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT111), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n797), .A2(new_n827), .A3(new_n376), .A4(new_n804), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n805), .A2(KEYINPUT111), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(new_n608), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n810), .B1(new_n830), .B2(new_n651), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n826), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n602), .B1(new_n793), .B2(new_n794), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT110), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n795), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n832), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT117), .B1(new_n837), .B2(new_n822), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n802), .A2(KEYINPUT117), .A3(new_n812), .A4(new_n822), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n840));
  AOI211_X1 g654(.A(new_n840), .B(new_n779), .C1(new_n786), .C2(new_n787), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n777), .B(new_n825), .C1(new_n838), .C2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT118), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n835), .B(new_n795), .C1(new_n826), .C2(new_n831), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n846), .B1(new_n847), .B2(new_n821), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n848), .A2(new_n839), .A3(new_n841), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(KEYINPUT118), .A3(new_n777), .A4(new_n825), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n847), .A2(new_n821), .ZN(new_n851));
  INV_X1    g665(.A(new_n824), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n851), .A2(KEYINPUT116), .A3(new_n788), .A4(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT116), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n854), .B1(new_n823), .B2(new_n824), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n823), .A2(new_n840), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n853), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  AOI22_X1  g671(.A1(new_n845), .A2(new_n850), .B1(KEYINPUT54), .B2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n707), .A2(new_n372), .A3(new_n754), .A4(new_n756), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n698), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n690), .A2(new_n372), .ZN(new_n862));
  NOR4_X1   g676(.A1(new_n862), .A2(new_n677), .A3(new_n544), .A4(new_n722), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(new_n629), .ZN(new_n864));
  INV_X1    g678(.A(G953), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n861), .A2(new_n864), .A3(G952), .A4(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n754), .A2(new_n756), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n862), .A2(new_n868), .A3(new_n722), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n601), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT48), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n867), .A2(new_n871), .A3(KEYINPUT120), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT120), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT48), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n870), .B(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n873), .B1(new_n875), .B2(new_n866), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n696), .A2(new_n497), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n767), .A2(new_n769), .A3(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n859), .A2(new_n748), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT51), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n668), .A2(new_n630), .A3(new_n669), .A4(new_n690), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n859), .A2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT50), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n884), .A2(KEYINPUT119), .A3(new_n885), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n885), .A2(KEYINPUT119), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n885), .A2(KEYINPUT119), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n887), .B(new_n888), .C1(new_n859), .C2(new_n883), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n612), .A2(new_n627), .ZN(new_n890));
  AOI22_X1  g704(.A1(new_n863), .A2(new_n890), .B1(new_n869), .B2(new_n819), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n886), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n881), .A2(new_n882), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n882), .B1(new_n881), .B2(new_n892), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n877), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(KEYINPUT121), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n877), .B(new_n897), .C1(new_n893), .C2(new_n894), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n776), .B1(new_n858), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n702), .A2(new_n491), .A3(new_n304), .ZN(new_n902));
  OR4_X1    g716(.A1(new_n612), .A2(new_n677), .A3(new_n753), .A4(new_n902), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n696), .B(KEYINPUT49), .Z(new_n904));
  NOR3_X1   g718(.A1(new_n903), .A2(new_n904), .A3(new_n670), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT122), .B1(new_n901), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n907));
  INV_X1    g721(.A(new_n905), .ZN(new_n908));
  AOI221_X4 g722(.A(new_n899), .B1(new_n857), .B2(KEYINPUT54), .C1(new_n845), .C2(new_n850), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n907), .B(new_n908), .C1(new_n909), .C2(new_n776), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n906), .A2(new_n910), .ZN(G75));
  AOI21_X1  g725(.A(new_n366), .B1(new_n849), .B2(new_n825), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(G210), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT56), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n241), .B(new_n273), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT55), .ZN(new_n916));
  AOI22_X1  g730(.A1(new_n915), .A2(new_n916), .B1(KEYINPUT123), .B2(new_n914), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n917), .B1(new_n916), .B2(new_n915), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n913), .A2(new_n914), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n918), .B1(new_n913), .B2(new_n914), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n310), .A2(G952), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(G51));
  NAND2_X1  g736(.A1(new_n849), .A2(new_n825), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(KEYINPUT54), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n843), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n740), .B(KEYINPUT57), .Z(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n927), .B1(new_n479), .B2(new_n480), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n912), .A2(new_n735), .A3(new_n737), .A4(new_n738), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n921), .B1(new_n928), .B2(new_n929), .ZN(G54));
  INV_X1    g744(.A(new_n921), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n912), .A2(KEYINPUT58), .A3(G475), .ZN(new_n932));
  INV_X1    g746(.A(new_n360), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n934), .B1(new_n933), .B2(new_n932), .ZN(G60));
  NAND2_X1  g749(.A1(G478), .A2(G902), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT59), .Z(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n925), .A2(new_n752), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n931), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n858), .A2(new_n937), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n940), .B1(new_n941), .B2(new_n624), .ZN(G63));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n943));
  NAND2_X1  g757(.A1(G217), .A2(G902), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT60), .Z(new_n945));
  AOI21_X1  g759(.A(new_n943), .B1(new_n923), .B2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n540), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n923), .A2(new_n943), .A3(new_n945), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n945), .ZN(new_n951));
  AOI211_X1 g765(.A(KEYINPUT124), .B(new_n951), .C1(new_n849), .C2(new_n825), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n645), .B1(new_n946), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n950), .A2(new_n953), .A3(new_n931), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT61), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n950), .A2(new_n953), .A3(KEYINPUT61), .A4(new_n931), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(G66));
  OAI21_X1  g772(.A(G953), .B1(new_n374), .B2(new_n271), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n778), .A2(new_n694), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n837), .A2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n310), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n959), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n241), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n965), .B1(G898), .B2(new_n310), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n964), .B(new_n966), .ZN(G69));
  INV_X1    g781(.A(new_n601), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n771), .B1(new_n629), .B2(new_n804), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n665), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n760), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n780), .A2(new_n720), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n682), .A2(KEYINPUT62), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(KEYINPUT62), .B1(new_n682), .B2(new_n973), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n774), .B(new_n971), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n976), .A2(new_n310), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n575), .B(new_n353), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT125), .Z(new_n979));
  OR2_X1    g793(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(G227), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n963), .B1(new_n981), .B2(new_n658), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n747), .A2(new_n968), .A3(new_n709), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n760), .A2(new_n983), .A3(new_n972), .ZN(new_n984));
  AND4_X1   g798(.A1(new_n729), .A2(new_n984), .A3(new_n731), .A4(new_n774), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n310), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n986), .B(new_n978), .C1(new_n658), .C2(new_n310), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n980), .A2(new_n982), .A3(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT126), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n988), .A2(new_n989), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n980), .A2(new_n987), .ZN(new_n992));
  OAI22_X1  g806(.A1(new_n990), .A2(new_n991), .B1(new_n982), .B2(new_n992), .ZN(G72));
  NAND2_X1  g807(.A1(new_n962), .A2(new_n985), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n671), .B(KEYINPUT63), .Z(new_n995));
  AND2_X1   g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n585), .A2(new_n564), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n995), .B1(new_n976), .B2(new_n961), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n585), .A2(new_n564), .ZN(new_n999));
  AND3_X1   g813(.A1(new_n998), .A2(KEYINPUT127), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(KEYINPUT127), .B1(new_n998), .B2(new_n999), .ZN(new_n1001));
  OAI221_X1 g815(.A(new_n931), .B1(new_n996), .B2(new_n997), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n672), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n596), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n1004), .A2(new_n995), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1002), .B1(new_n857), .B2(new_n1005), .ZN(G57));
endmodule


