//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n991, new_n992, new_n993, new_n995, new_n996, new_n997, new_n998,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1023, new_n1024, new_n1025;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT11), .ZN(new_n203));
  INV_X1    g002(.A(G169gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G197gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(KEYINPUT92), .B(KEYINPUT12), .Z(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT14), .ZN(new_n211));
  INV_X1    g010(.A(G29gat), .ZN(new_n212));
  INV_X1    g011(.A(G36gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n215));
  AOI22_X1  g014(.A1(new_n214), .A2(new_n215), .B1(G29gat), .B2(G36gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(G43gat), .B(G50gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT15), .ZN(new_n218));
  OR2_X1    g017(.A1(G43gat), .A2(G50gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT15), .ZN(new_n220));
  NAND2_X1  g019(.A1(G43gat), .A2(G50gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n216), .A2(new_n218), .A3(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT93), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n216), .A2(new_n218), .A3(KEYINPUT93), .A4(new_n222), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n216), .A2(new_n218), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT94), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n225), .A2(KEYINPUT94), .A3(new_n226), .A4(new_n227), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G15gat), .B(G22gat), .ZN(new_n233));
  INV_X1    g032(.A(G1gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(KEYINPUT16), .A3(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n235), .B1(new_n234), .B2(new_n233), .ZN(new_n236));
  XOR2_X1   g035(.A(new_n236), .B(G8gat), .Z(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n232), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT17), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n228), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n230), .A2(new_n240), .A3(new_n231), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT95), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT95), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n230), .A2(new_n244), .A3(new_n240), .A4(new_n231), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n241), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n239), .B1(new_n246), .B2(new_n238), .ZN(new_n247));
  NAND2_X1  g046(.A1(G229gat), .A2(G233gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(KEYINPUT18), .A3(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(new_n248), .B(KEYINPUT13), .Z(new_n250));
  INV_X1    g049(.A(new_n232), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n251), .A2(new_n237), .ZN(new_n252));
  INV_X1    g051(.A(new_n239), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n252), .B1(KEYINPUT96), .B2(new_n253), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n252), .A2(KEYINPUT96), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n250), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n249), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT18), .B1(new_n247), .B2(new_n248), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n210), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n247), .A2(new_n248), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT18), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n262), .A2(new_n209), .A3(new_n249), .A4(new_n256), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  XOR2_X1   g063(.A(G183gat), .B(G211gat), .Z(new_n265));
  XNOR2_X1  g064(.A(G127gat), .B(G155gat), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  XOR2_X1   g066(.A(G57gat), .B(G64gat), .Z(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT97), .ZN(new_n269));
  XNOR2_X1  g068(.A(G57gat), .B(G64gat), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT97), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(G71gat), .A2(G78gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(G71gat), .A2(G78gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT9), .ZN(new_n275));
  AOI22_X1  g074(.A1(new_n269), .A2(new_n272), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n274), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(new_n273), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n278), .B1(new_n268), .B2(KEYINPUT9), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT98), .B1(new_n280), .B2(KEYINPUT21), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT98), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT21), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n282), .B(new_n283), .C1(new_n276), .C2(new_n279), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n281), .A2(G231gat), .A3(G233gat), .A4(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  AOI22_X1  g085(.A1(new_n281), .A2(new_n284), .B1(G231gat), .B2(G233gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n267), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n281), .A2(new_n284), .ZN(new_n289));
  NAND2_X1  g088(.A1(G231gat), .A2(G233gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(new_n285), .A3(new_n266), .ZN(new_n292));
  XOR2_X1   g091(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  AND3_X1   g093(.A1(new_n288), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n294), .B1(new_n288), .B2(new_n292), .ZN(new_n296));
  INV_X1    g095(.A(new_n276), .ZN(new_n297));
  INV_X1    g096(.A(new_n279), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(KEYINPUT99), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT99), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n300), .B1(new_n276), .B2(new_n279), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n237), .B1(new_n302), .B2(KEYINPUT21), .ZN(new_n303));
  NOR3_X1   g102(.A1(new_n295), .A2(new_n296), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n303), .ZN(new_n305));
  INV_X1    g104(.A(new_n292), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n266), .B1(new_n291), .B2(new_n285), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n293), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n288), .A2(new_n292), .A3(new_n294), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n305), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n265), .B1(new_n304), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n303), .B1(new_n295), .B2(new_n296), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n308), .A2(new_n305), .A3(new_n309), .ZN(new_n313));
  INV_X1    g112(.A(new_n265), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(G99gat), .A2(G106gat), .ZN(new_n317));
  INV_X1    g116(.A(G85gat), .ZN(new_n318));
  INV_X1    g117(.A(G92gat), .ZN(new_n319));
  AOI22_X1  g118(.A1(KEYINPUT8), .A2(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT101), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n320), .B(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G99gat), .B(G106gat), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT102), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n323), .B(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(G85gat), .A2(G92gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n326), .B(KEYINPUT7), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n322), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT103), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n322), .A2(new_n325), .A3(KEYINPUT103), .A4(new_n327), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n322), .A2(new_n327), .ZN(new_n332));
  INV_X1    g131(.A(new_n325), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n330), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n280), .ZN(new_n336));
  AND2_X1   g135(.A1(new_n280), .A2(new_n328), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n335), .A2(new_n336), .B1(new_n337), .B2(new_n334), .ZN(new_n338));
  NAND2_X1  g137(.A1(G230gat), .A2(G233gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G120gat), .B(G148gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(G176gat), .B(G204gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n339), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n299), .A2(new_n301), .A3(KEYINPUT10), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n346), .A2(new_n335), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT104), .B(KEYINPUT10), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n347), .B1(new_n338), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n344), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  XOR2_X1   g149(.A(new_n339), .B(KEYINPUT105), .Z(new_n351));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n334), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n352), .A2(new_n353), .A3(new_n348), .ZN(new_n354));
  OR2_X1    g153(.A1(new_n346), .A2(new_n335), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n351), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n343), .B1(new_n356), .B2(new_n340), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n350), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n246), .A2(new_n335), .ZN(new_n360));
  NAND2_X1  g159(.A1(G232gat), .A2(G233gat), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT41), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n363), .B1(new_n232), .B2(new_n335), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n360), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G190gat), .B(G218gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n367), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n360), .A2(new_n365), .A3(new_n369), .ZN(new_n370));
  XOR2_X1   g169(.A(G134gat), .B(G162gat), .Z(new_n371));
  NAND3_X1  g170(.A1(new_n368), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n371), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n369), .B1(new_n360), .B2(new_n365), .ZN(new_n374));
  AOI211_X1 g173(.A(new_n364), .B(new_n367), .C1(new_n246), .C2(new_n335), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n362), .A2(KEYINPUT41), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(KEYINPUT100), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n372), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n378), .B1(new_n372), .B2(new_n376), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n316), .B(new_n359), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT106), .ZN(new_n382));
  INV_X1    g181(.A(new_n378), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n371), .B1(new_n368), .B2(new_n370), .ZN(new_n384));
  NOR3_X1   g183(.A1(new_n374), .A2(new_n375), .A3(new_n373), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n372), .A2(new_n376), .A3(new_n378), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT106), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n388), .A2(new_n389), .A3(new_n316), .A4(new_n359), .ZN(new_n390));
  AND2_X1   g189(.A1(new_n382), .A2(new_n390), .ZN(new_n391));
  AND2_X1   g190(.A1(G155gat), .A2(G162gat), .ZN(new_n392));
  NOR2_X1   g191(.A1(G155gat), .A2(G162gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(G141gat), .B(G148gat), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n394), .B1(new_n395), .B2(KEYINPUT2), .ZN(new_n396));
  XNOR2_X1  g195(.A(G155gat), .B(G162gat), .ZN(new_n397));
  INV_X1    g196(.A(G141gat), .ZN(new_n398));
  INV_X1    g197(.A(G148gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(G155gat), .ZN(new_n401));
  INV_X1    g200(.A(G162gat), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT2), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(G141gat), .A2(G148gat), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n397), .A2(new_n400), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n396), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT22), .ZN(new_n407));
  XNOR2_X1  g206(.A(KEYINPUT76), .B(G218gat), .ZN(new_n408));
  INV_X1    g207(.A(G211gat), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(G197gat), .B(G204gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G211gat), .B(G218gat), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n414), .A2(KEYINPUT77), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(KEYINPUT77), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n417), .A2(new_n410), .A3(new_n411), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT29), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT3), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n406), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(G228gat), .A2(G233gat), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n396), .A2(new_n405), .A3(new_n422), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT81), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n396), .A2(new_n405), .A3(KEYINPUT81), .A4(new_n422), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n419), .B1(new_n429), .B2(new_n420), .ZN(new_n430));
  NOR3_X1   g229(.A1(new_n423), .A2(new_n424), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(G218gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT76), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT76), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(G218gat), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n409), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n411), .B(new_n413), .C1(new_n436), .C2(KEYINPUT22), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n413), .B1(new_n410), .B2(new_n411), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n420), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n406), .B1(new_n440), .B2(new_n422), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n424), .B1(new_n430), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT85), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT85), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n444), .B(new_n424), .C1(new_n430), .C2(new_n441), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n431), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(G22gat), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT86), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n446), .A2(new_n447), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OR3_X1    g249(.A1(new_n423), .A2(new_n424), .A3(new_n430), .ZN(new_n451));
  INV_X1    g250(.A(new_n445), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n436), .A2(KEYINPUT22), .ZN(new_n453));
  INV_X1    g252(.A(new_n411), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n414), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n437), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT3), .B1(new_n456), .B2(new_n420), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT29), .B1(new_n427), .B2(new_n428), .ZN(new_n458));
  OAI22_X1  g257(.A1(new_n457), .A2(new_n406), .B1(new_n458), .B2(new_n419), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n444), .B1(new_n459), .B2(new_n424), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n451), .B1(new_n452), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT86), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n462), .A3(G22gat), .ZN(new_n463));
  XOR2_X1   g262(.A(G78gat), .B(G106gat), .Z(new_n464));
  XNOR2_X1  g263(.A(new_n464), .B(KEYINPUT84), .ZN(new_n465));
  XOR2_X1   g264(.A(KEYINPUT31), .B(G50gat), .Z(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT87), .B1(new_n450), .B2(new_n468), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n447), .B(new_n451), .C1(new_n452), .C2(new_n460), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n462), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n461), .A2(G22gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT87), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n473), .A2(new_n474), .A3(new_n463), .A4(new_n467), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n472), .A2(new_n470), .ZN(new_n476));
  INV_X1    g275(.A(new_n467), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n469), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  XOR2_X1   g278(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n480));
  NOR2_X1   g279(.A1(G169gat), .A2(G176gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT23), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT23), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n483), .B1(G169gat), .B2(G176gat), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n482), .B1(new_n484), .B2(new_n481), .ZN(new_n485));
  AND3_X1   g284(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(G183gat), .A2(G190gat), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n480), .B1(new_n485), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT65), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT65), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n492), .B(new_n480), .C1(new_n485), .C2(new_n489), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n485), .A2(new_n489), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT25), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n491), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT27), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(G183gat), .ZN(new_n498));
  INV_X1    g297(.A(G183gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT27), .ZN(new_n500));
  INV_X1    g299(.A(G190gat), .ZN(new_n501));
  AND4_X1   g300(.A1(KEYINPUT28), .A2(new_n498), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT66), .B1(new_n499), .B2(KEYINPUT27), .ZN(new_n503));
  XNOR2_X1  g302(.A(KEYINPUT27), .B(G183gat), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n501), .B(new_n503), .C1(new_n504), .C2(KEYINPUT66), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT28), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n502), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT68), .ZN(new_n508));
  NAND2_X1  g307(.A1(G169gat), .A2(G176gat), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT26), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(G176gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n204), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT67), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n481), .A2(KEYINPUT67), .A3(new_n510), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n487), .ZN(new_n518));
  NOR3_X1   g317(.A1(new_n507), .A2(new_n508), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT66), .B1(new_n498), .B2(new_n500), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n501), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n506), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n502), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n515), .A2(new_n516), .B1(G183gat), .B2(G190gat), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT68), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n496), .B1(new_n519), .B2(new_n526), .ZN(new_n527));
  XOR2_X1   g326(.A(G113gat), .B(G120gat), .Z(new_n528));
  INV_X1    g327(.A(KEYINPUT1), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(G134gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(G127gat), .ZN(new_n532));
  INV_X1    g331(.A(G127gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(G134gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n532), .A2(new_n534), .A3(new_n529), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT69), .ZN(new_n538));
  INV_X1    g337(.A(G113gat), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n538), .B1(new_n539), .B2(G120gat), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT70), .ZN(new_n541));
  INV_X1    g340(.A(G120gat), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n541), .B1(new_n542), .B2(G113gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n542), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n539), .A2(KEYINPUT70), .A3(G120gat), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n540), .A2(new_n543), .A3(new_n544), .A4(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT71), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n537), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AND2_X1   g347(.A1(new_n543), .A2(new_n545), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n549), .A2(KEYINPUT71), .A3(new_n540), .A4(new_n544), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT72), .ZN(new_n551));
  AND3_X1   g350(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n551), .B1(new_n548), .B2(new_n550), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n536), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NOR3_X1   g353(.A1(new_n527), .A2(new_n554), .A3(KEYINPUT73), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n498), .A2(new_n500), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT66), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(G190gat), .B1(new_n498), .B2(KEYINPUT66), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT28), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n525), .B1(new_n560), .B2(new_n502), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n508), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n524), .A2(KEYINPUT68), .A3(new_n525), .ZN(new_n563));
  INV_X1    g362(.A(new_n480), .ZN(new_n564));
  NOR3_X1   g363(.A1(new_n483), .A2(G169gat), .A3(G176gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n509), .A2(KEYINPUT23), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n565), .B1(new_n513), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n488), .A2(new_n487), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT24), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n568), .B1(new_n569), .B2(new_n487), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n564), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g370(.A1(new_n571), .A2(new_n492), .B1(new_n494), .B2(KEYINPUT25), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n562), .A2(new_n563), .B1(new_n572), .B2(new_n491), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n548), .A2(new_n550), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT72), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(new_n576));
  AOI22_X1  g375(.A1(new_n575), .A2(new_n576), .B1(new_n530), .B2(new_n535), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT73), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n579), .B1(new_n573), .B2(new_n577), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n555), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G227gat), .A2(G233gat), .ZN(new_n582));
  OAI21_X1  g381(.A(KEYINPUT32), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT33), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n584), .B1(new_n581), .B2(new_n582), .ZN(new_n585));
  XNOR2_X1  g384(.A(G15gat), .B(G43gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT74), .ZN(new_n587));
  XOR2_X1   g386(.A(G71gat), .B(G99gat), .Z(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n583), .A2(new_n585), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n573), .A2(new_n579), .A3(new_n577), .ZN(new_n591));
  AOI21_X1  g390(.A(KEYINPUT73), .B1(new_n527), .B2(new_n554), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n527), .A2(new_n554), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n582), .B(new_n591), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT34), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT32), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n598));
  INV_X1    g397(.A(new_n582), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n589), .B(KEYINPUT75), .Z(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT33), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  AND3_X1   g402(.A1(new_n590), .A2(new_n596), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n596), .B1(new_n590), .B2(new_n603), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n479), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT91), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(KEYINPUT83), .B(KEYINPUT6), .ZN(new_n610));
  XNOR2_X1  g409(.A(G1gat), .B(G29gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT0), .ZN(new_n612));
  XNOR2_X1  g411(.A(G57gat), .B(G85gat), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n612), .B(new_n613), .Z(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n554), .B(new_n429), .C1(new_n422), .C2(new_n406), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n577), .A2(KEYINPUT4), .A3(new_n406), .ZN(new_n617));
  NAND2_X1  g416(.A1(G225gat), .A2(G233gat), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n536), .B(new_n406), .C1(new_n552), .C2(new_n553), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT4), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n616), .A2(new_n617), .A3(new_n618), .A4(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(KEYINPUT82), .B(KEYINPUT5), .Z(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n618), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n577), .A2(new_n406), .ZN(new_n626));
  INV_X1    g425(.A(new_n619), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n622), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n615), .B(new_n624), .C1(new_n629), .C2(new_n623), .ZN(new_n630));
  INV_X1    g429(.A(new_n624), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n623), .B1(new_n622), .B2(new_n628), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n614), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n610), .B1(new_n630), .B2(new_n633), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n630), .A2(new_n610), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AND2_X1   g435(.A1(G226gat), .A2(G233gat), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n573), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n496), .A2(new_n561), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(KEYINPUT78), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT78), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n496), .A2(new_n641), .A3(new_n561), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n637), .A2(KEYINPUT29), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n638), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(new_n419), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT79), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n562), .A2(new_n563), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n645), .B1(new_n649), .B2(new_n496), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n650), .B1(new_n643), .B2(new_n637), .ZN(new_n651));
  INV_X1    g450(.A(new_n419), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n648), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n642), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n641), .B1(new_n496), .B2(new_n561), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n637), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n650), .ZN(new_n657));
  AND4_X1   g456(.A1(new_n648), .A2(new_n656), .A3(new_n652), .A4(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n647), .B1(new_n653), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G8gat), .B(G36gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(G64gat), .B(G92gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n656), .A2(new_n657), .A3(new_n652), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT79), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n651), .A2(new_n648), .A3(new_n652), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n662), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n667), .A2(KEYINPUT30), .A3(new_n668), .A4(new_n647), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n663), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(KEYINPUT80), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n668), .B(new_n647), .C1(new_n653), .C2(new_n658), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT30), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT80), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n663), .A2(new_n669), .A3(new_n675), .ZN(new_n676));
  AND4_X1   g475(.A1(new_n636), .A2(new_n671), .A3(new_n674), .A4(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n479), .A2(new_n606), .A3(KEYINPUT91), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n609), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n674), .A2(new_n663), .A3(new_n669), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n636), .ZN(new_n682));
  AOI21_X1  g481(.A(KEYINPUT35), .B1(new_n682), .B2(KEYINPUT89), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT90), .B1(new_n604), .B2(new_n605), .ZN(new_n684));
  INV_X1    g483(.A(new_n596), .ZN(new_n685));
  AOI21_X1  g484(.A(KEYINPUT33), .B1(new_n598), .B2(new_n599), .ZN(new_n686));
  INV_X1    g485(.A(new_n589), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n600), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n603), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n685), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n590), .A2(new_n596), .A3(new_n603), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT90), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n684), .A2(new_n479), .A3(new_n693), .ZN(new_n694));
  NOR4_X1   g493(.A1(new_n680), .A2(new_n634), .A3(new_n635), .A4(KEYINPUT89), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI22_X1  g495(.A1(new_n679), .A2(KEYINPUT35), .B1(new_n683), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(KEYINPUT36), .B1(new_n604), .B2(new_n605), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT36), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n690), .A2(new_n691), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n616), .A2(new_n617), .A3(new_n621), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n625), .ZN(new_n703));
  OR3_X1    g502(.A1(new_n626), .A2(new_n625), .A3(new_n627), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(KEYINPUT39), .A3(new_n704), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n705), .B(new_n614), .C1(KEYINPUT39), .C2(new_n703), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT40), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n707), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n680), .A2(new_n708), .A3(new_n630), .A4(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT37), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n711), .B(new_n647), .C1(new_n653), .C2(new_n658), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(new_n662), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n711), .B1(new_n667), .B2(new_n647), .ZN(new_n714));
  OAI21_X1  g513(.A(KEYINPUT38), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n711), .B1(new_n651), .B2(new_n419), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n646), .A2(new_n652), .ZN(new_n717));
  AOI21_X1  g516(.A(KEYINPUT38), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n712), .A2(new_n718), .A3(new_n662), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT88), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n712), .A2(new_n718), .A3(KEYINPUT88), .A4(new_n662), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n715), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n672), .B1(new_n634), .B2(new_n635), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n710), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n479), .ZN(new_n726));
  INV_X1    g525(.A(new_n479), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n677), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n701), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n264), .B(new_n391), .C1(new_n697), .C2(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(new_n636), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(new_n234), .ZN(G1324gat));
  OR2_X1    g531(.A1(new_n730), .A2(new_n681), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT16), .B(G8gat), .Z(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(KEYINPUT42), .ZN(new_n735));
  OR3_X1    g534(.A1(new_n733), .A2(KEYINPUT108), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n734), .B(KEYINPUT107), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n737), .A2(KEYINPUT42), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT42), .ZN(new_n739));
  OAI22_X1  g538(.A1(new_n733), .A2(new_n738), .B1(new_n739), .B2(G8gat), .ZN(new_n740));
  OAI21_X1  g539(.A(KEYINPUT108), .B1(new_n733), .B2(new_n735), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n736), .A2(new_n740), .A3(new_n741), .ZN(G1325gat));
  NOR3_X1   g541(.A1(new_n604), .A2(new_n605), .A3(KEYINPUT36), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n699), .B1(new_n690), .B2(new_n691), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT109), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n698), .A2(new_n746), .A3(new_n700), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(G15gat), .B1(new_n730), .B2(new_n749), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n684), .A2(new_n693), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  OR2_X1    g551(.A1(new_n752), .A2(G15gat), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n750), .B1(new_n730), .B2(new_n753), .ZN(G1326gat));
  NOR2_X1   g553(.A1(new_n730), .A2(new_n479), .ZN(new_n755));
  XOR2_X1   g554(.A(KEYINPUT43), .B(G22gat), .Z(new_n756));
  XNOR2_X1  g555(.A(new_n755), .B(new_n756), .ZN(G1327gat));
  INV_X1    g556(.A(new_n316), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n359), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(new_n388), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n264), .B(new_n760), .C1(new_n697), .C2(new_n729), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n761), .A2(G29gat), .A3(new_n636), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n762), .B(KEYINPUT45), .Z(new_n763));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n679), .A2(KEYINPUT35), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n696), .A2(new_n683), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n726), .A2(new_n728), .ZN(new_n767));
  AOI22_X1  g566(.A1(new_n765), .A2(new_n766), .B1(new_n767), .B2(new_n749), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n764), .B1(new_n768), .B2(new_n388), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n379), .A2(new_n380), .ZN(new_n770));
  OAI211_X1 g569(.A(KEYINPUT44), .B(new_n770), .C1(new_n697), .C2(new_n729), .ZN(new_n771));
  INV_X1    g570(.A(new_n264), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n759), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n769), .A2(new_n771), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(G29gat), .B1(new_n774), .B2(new_n636), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n763), .A2(new_n775), .ZN(G1328gat));
  NOR3_X1   g575(.A1(new_n761), .A2(G36gat), .A3(new_n681), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT46), .ZN(new_n778));
  OAI21_X1  g577(.A(G36gat), .B1(new_n774), .B2(new_n681), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(G1329gat));
  OAI21_X1  g579(.A(G43gat), .B1(new_n774), .B2(new_n749), .ZN(new_n781));
  OR3_X1    g580(.A1(new_n761), .A2(G43gat), .A3(new_n752), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT47), .B1(new_n783), .B2(KEYINPUT110), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT110), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT47), .ZN(new_n786));
  AOI211_X1 g585(.A(new_n785), .B(new_n786), .C1(new_n781), .C2(new_n782), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n784), .A2(new_n787), .ZN(G1330gat));
  INV_X1    g587(.A(KEYINPUT48), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n761), .A2(G50gat), .A3(new_n479), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(KEYINPUT112), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n769), .A2(new_n727), .A3(new_n771), .A4(new_n773), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n790), .B1(new_n794), .B2(G50gat), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n796), .B(new_n789), .C1(new_n790), .C2(new_n791), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n793), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n795), .B1(new_n793), .B2(new_n797), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n798), .A2(new_n799), .ZN(G1331gat));
  NAND4_X1  g599(.A1(new_n388), .A2(new_n772), .A3(new_n316), .A4(new_n358), .ZN(new_n801));
  OR3_X1    g600(.A1(new_n768), .A2(KEYINPUT113), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(KEYINPUT113), .B1(new_n768), .B2(new_n801), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n636), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g606(.A(new_n681), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n804), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n810));
  XOR2_X1   g609(.A(new_n809), .B(new_n810), .Z(G1333gat));
  NAND3_X1  g610(.A1(new_n802), .A2(new_n748), .A3(new_n803), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(G71gat), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n752), .A2(G71gat), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n802), .A2(new_n803), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT50), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n816), .B(new_n817), .ZN(G1334gat));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n727), .A3(new_n803), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(KEYINPUT115), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n802), .A2(new_n821), .A3(new_n727), .A4(new_n803), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g622(.A(KEYINPUT114), .B(G78gat), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n823), .B(new_n824), .ZN(G1335gat));
  NOR3_X1   g624(.A1(new_n264), .A2(new_n316), .A3(new_n359), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n769), .A2(new_n771), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(G85gat), .B1(new_n827), .B2(new_n636), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n264), .A2(new_n316), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n748), .B1(new_n726), .B2(new_n728), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n770), .B(new_n829), .C1(new_n697), .C2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT51), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT116), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT116), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n831), .A2(new_n835), .A3(new_n832), .ZN(new_n836));
  INV_X1    g635(.A(new_n830), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n765), .A2(new_n766), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n839), .A2(KEYINPUT51), .A3(new_n770), .A4(new_n829), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n834), .A2(new_n836), .A3(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n805), .A2(new_n318), .A3(new_n358), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n828), .B1(new_n842), .B2(new_n843), .ZN(G1336gat));
  XNOR2_X1  g643(.A(KEYINPUT118), .B(KEYINPUT52), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n769), .A2(new_n680), .A3(new_n771), .A4(new_n826), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n845), .B1(new_n846), .B2(G92gat), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n681), .A2(G92gat), .A3(new_n359), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n836), .A2(new_n840), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n835), .B1(new_n831), .B2(new_n832), .ZN(new_n850));
  OAI211_X1 g649(.A(KEYINPUT117), .B(new_n848), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT117), .B1(new_n841), .B2(new_n848), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n847), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n846), .A2(G92gat), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n840), .A2(new_n833), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n856), .A2(new_n848), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT52), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n854), .A2(new_n858), .ZN(G1337gat));
  OAI21_X1  g658(.A(G99gat), .B1(new_n827), .B2(new_n749), .ZN(new_n860));
  OR3_X1    g659(.A1(new_n752), .A2(G99gat), .A3(new_n359), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n860), .B1(new_n842), .B2(new_n861), .ZN(G1338gat));
  NOR3_X1   g661(.A1(new_n479), .A2(G106gat), .A3(new_n359), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n841), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n769), .A2(new_n727), .A3(new_n771), .A4(new_n826), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(G106gat), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI22_X1  g667(.A1(new_n865), .A2(G106gat), .B1(new_n856), .B2(new_n863), .ZN(new_n869));
  OAI22_X1  g668(.A1(new_n864), .A2(new_n868), .B1(new_n867), .B2(new_n869), .ZN(G1339gat));
  NOR2_X1   g669(.A1(new_n381), .A2(new_n264), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT55), .ZN(new_n872));
  INV_X1    g671(.A(new_n343), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n873), .B1(new_n356), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n354), .A2(new_n355), .A3(new_n351), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n876), .B(KEYINPUT54), .C1(new_n349), .C2(new_n345), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT119), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n354), .A2(new_n355), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n874), .B1(new_n880), .B2(new_n339), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT119), .B1(new_n881), .B2(new_n876), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n872), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT120), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI211_X1 g684(.A(KEYINPUT120), .B(new_n872), .C1(new_n879), .C2(new_n882), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n207), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n254), .A2(new_n255), .A3(new_n250), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n247), .A2(new_n248), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n263), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n878), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n881), .A2(KEYINPUT119), .A3(new_n876), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n893), .A2(new_n894), .A3(KEYINPUT55), .A4(new_n875), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n895), .A2(new_n350), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n770), .A2(new_n887), .A3(new_n892), .A4(new_n896), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n263), .A2(new_n358), .A3(new_n891), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n895), .A2(new_n350), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n899), .B1(new_n259), .B2(new_n263), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n898), .B1(new_n900), .B2(new_n887), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n897), .B1(new_n901), .B2(new_n770), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n871), .B1(new_n902), .B2(new_n758), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n903), .A2(new_n636), .A3(new_n680), .ZN(new_n904));
  INV_X1    g703(.A(new_n694), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n906), .A2(new_n539), .A3(new_n772), .ZN(new_n907));
  INV_X1    g706(.A(new_n609), .ZN(new_n908));
  INV_X1    g707(.A(new_n678), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n904), .A2(new_n910), .A3(new_n264), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n907), .B1(new_n539), .B2(new_n911), .ZN(G1340gat));
  NOR3_X1   g711(.A1(new_n906), .A2(new_n542), .A3(new_n359), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n904), .A2(new_n910), .A3(new_n358), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n913), .B1(new_n542), .B2(new_n914), .ZN(G1341gat));
  OAI21_X1  g714(.A(G127gat), .B1(new_n906), .B2(new_n758), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n904), .A2(new_n533), .A3(new_n910), .A4(new_n316), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1342gat));
  NOR2_X1   g717(.A1(new_n903), .A2(new_n636), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n388), .A2(new_n680), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n919), .A2(new_n531), .A3(new_n910), .A4(new_n920), .ZN(new_n921));
  XOR2_X1   g720(.A(new_n921), .B(KEYINPUT56), .Z(new_n922));
  OAI21_X1  g721(.A(G134gat), .B1(new_n906), .B2(new_n388), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1343gat));
  AOI21_X1  g723(.A(new_n898), .B1(new_n900), .B2(new_n883), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n897), .B1(new_n925), .B2(new_n770), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n871), .B1(new_n926), .B2(new_n758), .ZN(new_n927));
  OAI21_X1  g726(.A(KEYINPUT57), .B1(new_n927), .B2(new_n479), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n748), .A2(new_n636), .A3(new_n680), .ZN(new_n929));
  INV_X1    g728(.A(new_n903), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n727), .ZN(new_n931));
  OAI211_X1 g730(.A(new_n928), .B(new_n929), .C1(new_n931), .C2(KEYINPUT57), .ZN(new_n932));
  OAI21_X1  g731(.A(G141gat), .B1(new_n932), .B2(new_n772), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n748), .A2(new_n479), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n904), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(new_n398), .A3(new_n264), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT58), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT121), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n938), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n937), .B(new_n940), .ZN(G1344gat));
  NAND3_X1  g740(.A1(new_n935), .A2(new_n399), .A3(new_n358), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT59), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n479), .A2(KEYINPUT57), .ZN(new_n944));
  AND4_X1   g743(.A1(new_n770), .A2(new_n887), .A3(new_n892), .A4(new_n896), .ZN(new_n945));
  INV_X1    g744(.A(new_n898), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n264), .A2(new_n896), .A3(new_n883), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n770), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g747(.A(KEYINPUT123), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT123), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n950), .B(new_n897), .C1(new_n925), .C2(new_n770), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n316), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n382), .A2(new_n772), .A3(new_n390), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT122), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n382), .A2(new_n390), .A3(KEYINPUT122), .A4(new_n772), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n944), .B1(new_n952), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g757(.A(KEYINPUT57), .B1(new_n903), .B2(new_n479), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n958), .A2(new_n959), .A3(new_n358), .A4(new_n929), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n399), .B1(new_n961), .B2(KEYINPUT124), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT124), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n943), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n932), .A2(new_n359), .ZN(new_n966));
  NOR3_X1   g765(.A1(new_n966), .A2(KEYINPUT59), .A3(new_n399), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n942), .B1(new_n965), .B2(new_n967), .ZN(G1345gat));
  OAI21_X1  g767(.A(G155gat), .B1(new_n932), .B2(new_n758), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n935), .A2(new_n401), .A3(new_n316), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(G1346gat));
  OAI21_X1  g770(.A(G162gat), .B1(new_n932), .B2(new_n388), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n919), .A2(new_n402), .A3(new_n920), .A4(new_n934), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n974), .B(KEYINPUT125), .ZN(G1347gat));
  NOR2_X1   g774(.A1(new_n805), .A2(new_n681), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n908), .A2(new_n977), .A3(new_n909), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n930), .A2(new_n978), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n980), .A2(new_n204), .A3(new_n264), .ZN(new_n981));
  NOR3_X1   g780(.A1(new_n903), .A2(new_n694), .A3(new_n977), .ZN(new_n982));
  INV_X1    g781(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g782(.A(G169gat), .B1(new_n983), .B2(new_n772), .ZN(new_n984));
  AND2_X1   g783(.A1(new_n984), .A2(KEYINPUT126), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n984), .A2(KEYINPUT126), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n981), .B1(new_n985), .B2(new_n986), .ZN(G1348gat));
  OAI21_X1  g786(.A(G176gat), .B1(new_n983), .B2(new_n359), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n980), .A2(new_n512), .A3(new_n358), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n988), .A2(new_n989), .ZN(G1349gat));
  NOR3_X1   g789(.A1(new_n979), .A2(new_n556), .A3(new_n758), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n499), .B1(new_n982), .B2(new_n316), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  XOR2_X1   g792(.A(new_n993), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g793(.A1(new_n980), .A2(new_n501), .A3(new_n770), .ZN(new_n995));
  OAI21_X1  g794(.A(G190gat), .B1(new_n983), .B2(new_n388), .ZN(new_n996));
  AND2_X1   g795(.A1(new_n996), .A2(KEYINPUT61), .ZN(new_n997));
  NOR2_X1   g796(.A1(new_n996), .A2(KEYINPUT61), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n995), .B1(new_n997), .B2(new_n998), .ZN(G1351gat));
  NOR2_X1   g798(.A1(new_n903), .A2(new_n479), .ZN(new_n1000));
  NOR2_X1   g799(.A1(new_n748), .A2(new_n977), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g801(.A(new_n206), .B1(new_n1002), .B2(new_n772), .ZN(new_n1003));
  NOR2_X1   g802(.A1(new_n772), .A2(new_n206), .ZN(new_n1004));
  NAND4_X1  g803(.A1(new_n958), .A2(new_n959), .A3(new_n1001), .A4(new_n1004), .ZN(new_n1005));
  AND2_X1   g804(.A1(new_n1003), .A2(new_n1005), .ZN(G1352gat));
  NAND4_X1  g805(.A1(new_n958), .A2(new_n959), .A3(new_n358), .A4(new_n1001), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1007), .A2(G204gat), .ZN(new_n1008));
  INV_X1    g807(.A(new_n1002), .ZN(new_n1009));
  NOR2_X1   g808(.A1(new_n359), .A2(G204gat), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g810(.A(KEYINPUT127), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g812(.A1(new_n1009), .A2(KEYINPUT127), .A3(new_n1010), .ZN(new_n1014));
  AND3_X1   g813(.A1(new_n1013), .A2(KEYINPUT62), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g814(.A(KEYINPUT62), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1016));
  OAI21_X1  g815(.A(new_n1008), .B1(new_n1015), .B2(new_n1016), .ZN(G1353gat));
  NAND3_X1  g816(.A1(new_n1009), .A2(new_n409), .A3(new_n316), .ZN(new_n1018));
  NAND4_X1  g817(.A1(new_n958), .A2(new_n959), .A3(new_n316), .A4(new_n1001), .ZN(new_n1019));
  AND3_X1   g818(.A1(new_n1019), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1020));
  AOI21_X1  g819(.A(KEYINPUT63), .B1(new_n1019), .B2(G211gat), .ZN(new_n1021));
  OAI21_X1  g820(.A(new_n1018), .B1(new_n1020), .B2(new_n1021), .ZN(G1354gat));
  OAI21_X1  g821(.A(new_n432), .B1(new_n1002), .B2(new_n388), .ZN(new_n1023));
  NOR2_X1   g822(.A1(new_n388), .A2(new_n408), .ZN(new_n1024));
  NAND4_X1  g823(.A1(new_n958), .A2(new_n959), .A3(new_n1001), .A4(new_n1024), .ZN(new_n1025));
  AND2_X1   g824(.A1(new_n1023), .A2(new_n1025), .ZN(G1355gat));
endmodule


