//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 0 1 0 1 0 0 1 0 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 0 1 0 1 1 1 1 0 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT79), .ZN(new_n188));
  INV_X1    g002(.A(G237), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  NAND4_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G143), .A4(G214), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT64), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT64), .A2(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  AND3_X1   g010(.A1(new_n189), .A2(new_n190), .A3(G214), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n188), .B(new_n191), .C1(new_n196), .C2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(KEYINPUT79), .A3(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT17), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n198), .A2(G131), .A3(new_n199), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT81), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n202), .A2(KEYINPUT81), .A3(new_n203), .A4(new_n204), .ZN(new_n208));
  INV_X1    g022(.A(G140), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G125), .ZN(new_n210));
  INV_X1    g024(.A(G125), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G140), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n210), .A2(new_n212), .A3(KEYINPUT16), .ZN(new_n213));
  OR3_X1    g027(.A1(new_n211), .A2(KEYINPUT16), .A3(G140), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(G146), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(G146), .B1(new_n213), .B2(new_n214), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n198), .A2(KEYINPUT17), .A3(G131), .A4(new_n199), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n207), .A2(new_n208), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n204), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT18), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n210), .A2(new_n212), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT80), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(G125), .B(G140), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT80), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n226), .A2(new_n228), .A3(G146), .ZN(new_n229));
  INV_X1    g043(.A(G146), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT18), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n200), .B1(new_n233), .B2(new_n201), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n223), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n221), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(G113), .B(G122), .ZN(new_n237));
  INV_X1    g051(.A(G104), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT83), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n187), .B1(new_n236), .B2(new_n241), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n223), .A2(new_n232), .A3(new_n234), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n208), .A2(new_n220), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n243), .B1(new_n244), .B2(new_n207), .ZN(new_n245));
  INV_X1    g059(.A(new_n241), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(G475), .B1(new_n242), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT20), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n202), .A2(new_n204), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT19), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n251), .B1(new_n226), .B2(new_n228), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n227), .A2(KEYINPUT19), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n230), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n250), .A2(new_n215), .A3(new_n254), .ZN(new_n255));
  AND3_X1   g069(.A1(new_n235), .A2(new_n255), .A3(new_n240), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n256), .B1(new_n236), .B2(new_n239), .ZN(new_n257));
  NOR2_X1   g071(.A1(G475), .A2(G902), .ZN(new_n258));
  XOR2_X1   g072(.A(new_n258), .B(KEYINPUT82), .Z(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n249), .B1(new_n257), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n240), .B1(new_n221), .B2(new_n235), .ZN(new_n262));
  NOR4_X1   g076(.A1(new_n262), .A2(new_n256), .A3(KEYINPUT20), .A4(new_n259), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n248), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT87), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT85), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n194), .A2(G128), .A3(new_n195), .ZN(new_n267));
  INV_X1    g081(.A(G134), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n267), .B(new_n268), .C1(G128), .C2(new_n193), .ZN(new_n269));
  INV_X1    g083(.A(G116), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n270), .A2(G122), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT84), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n272), .A2(new_n270), .A3(G122), .ZN(new_n273));
  INV_X1    g087(.A(G122), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT84), .B1(new_n274), .B2(G116), .ZN(new_n275));
  AOI211_X1 g089(.A(G107), .B(new_n271), .C1(new_n273), .C2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G107), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n273), .ZN(new_n278));
  INV_X1    g092(.A(new_n271), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n269), .B1(new_n276), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT13), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n194), .A2(new_n282), .A3(G128), .A4(new_n195), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G134), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n193), .A2(G128), .ZN(new_n285));
  AND2_X1   g099(.A1(KEYINPUT64), .A2(G143), .ZN(new_n286));
  NOR2_X1   g100(.A1(KEYINPUT64), .A2(G143), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n285), .B1(new_n288), .B2(G128), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n284), .B1(KEYINPUT13), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n266), .B1(new_n281), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n278), .A2(new_n279), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G107), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n278), .A2(new_n277), .A3(new_n279), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n267), .B(KEYINPUT13), .C1(G128), .C2(new_n193), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n296), .A2(G134), .A3(new_n283), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n295), .A2(new_n297), .A3(KEYINPUT85), .A4(new_n269), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT14), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n275), .A2(new_n273), .A3(new_n299), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n300), .A2(new_n279), .ZN(new_n301));
  AOI21_X1  g115(.A(KEYINPUT86), .B1(new_n278), .B2(KEYINPUT14), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT86), .ZN(new_n303));
  AOI211_X1 g117(.A(new_n303), .B(new_n299), .C1(new_n275), .C2(new_n273), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n301), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G107), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n267), .B1(G128), .B2(new_n193), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G134), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n276), .B1(new_n308), .B2(new_n269), .ZN(new_n309));
  AOI22_X1  g123(.A1(new_n291), .A2(new_n298), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT9), .B(G234), .ZN(new_n311));
  INV_X1    g125(.A(G217), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n311), .A2(new_n312), .A3(G953), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n265), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n306), .A2(new_n309), .ZN(new_n315));
  AOI22_X1  g129(.A1(new_n293), .A2(new_n294), .B1(new_n268), .B2(new_n289), .ZN(new_n316));
  AOI21_X1  g130(.A(KEYINPUT85), .B1(new_n316), .B2(new_n297), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n281), .A2(new_n290), .A3(new_n266), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n315), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n313), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n314), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n319), .A2(new_n265), .A3(new_n320), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(new_n187), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G478), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n325), .A2(KEYINPUT15), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n190), .A2(G952), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n328), .B1(G234), .B2(G237), .ZN(new_n329));
  NAND2_X1  g143(.A1(G234), .A2(G237), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(G902), .A3(G953), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(KEYINPUT88), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT21), .B(G898), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n329), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n326), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n322), .A2(new_n187), .A3(new_n323), .A4(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n327), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n264), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(G214), .B1(G237), .B2(G902), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n194), .A2(G146), .A3(new_n195), .ZN(new_n342));
  AND2_X1   g156(.A1(KEYINPUT0), .A2(G128), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n193), .A2(G146), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  AND3_X1   g159(.A1(new_n342), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(KEYINPUT0), .B(G128), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n230), .B1(new_n286), .B2(new_n287), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n230), .A2(G143), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n347), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(G125), .B1(new_n346), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT1), .ZN(new_n353));
  OAI21_X1  g167(.A(G128), .B1(new_n344), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(G146), .B1(new_n194), .B2(new_n195), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n354), .B1(new_n355), .B2(new_n349), .ZN(new_n356));
  INV_X1    g170(.A(G128), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n357), .A2(KEYINPUT1), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n342), .A2(new_n345), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(new_n211), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n352), .A2(KEYINPUT76), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT7), .ZN(new_n362));
  INV_X1    g176(.A(G224), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n363), .A2(G953), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT76), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n356), .A2(new_n366), .A3(new_n211), .A4(new_n359), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n361), .A2(new_n362), .A3(new_n365), .A4(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT3), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n369), .B1(new_n238), .B2(G107), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n277), .A2(KEYINPUT3), .A3(G104), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n277), .A2(G104), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G101), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT4), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n373), .B1(new_n370), .B2(new_n371), .ZN(new_n378));
  INV_X1    g192(.A(G101), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G113), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT2), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT2), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G113), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(G116), .B(G119), .ZN(new_n387));
  OR2_X1    g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n387), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n375), .A2(new_n377), .A3(G101), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n381), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n270), .A2(G119), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT5), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n382), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G119), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G116), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n270), .A2(G119), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n398), .A3(KEYINPUT5), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n395), .A2(new_n399), .B1(new_n387), .B2(new_n386), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT73), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n401), .B1(new_n277), .B2(G104), .ZN(new_n402));
  OAI21_X1  g216(.A(KEYINPUT72), .B1(new_n238), .B2(G107), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT72), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(new_n277), .A3(G104), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n238), .A2(KEYINPUT73), .A3(G107), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n402), .A2(new_n403), .A3(new_n405), .A4(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G101), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n378), .A2(new_n379), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n400), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT75), .ZN(new_n411));
  XOR2_X1   g225(.A(G110), .B(G122), .Z(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT75), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n400), .A2(new_n408), .A3(new_n414), .A4(new_n409), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n392), .A2(new_n411), .A3(new_n413), .A4(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT77), .B(KEYINPUT8), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n412), .B(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n410), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n400), .B1(new_n409), .B2(new_n408), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n368), .A2(new_n416), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n361), .A2(new_n367), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n364), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n361), .A2(new_n365), .A3(new_n367), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n365), .A2(new_n362), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(G902), .B1(new_n422), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(G210), .B1(G237), .B2(G902), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n392), .A2(new_n411), .A3(new_n415), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n412), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(KEYINPUT6), .A3(new_n416), .ZN(new_n432));
  INV_X1    g246(.A(new_n425), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n365), .B1(new_n361), .B2(new_n367), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT6), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n430), .A2(new_n436), .A3(new_n412), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n432), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n428), .A2(new_n429), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n429), .B1(new_n428), .B2(new_n438), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n341), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT78), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT78), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n443), .B(new_n341), .C1(new_n439), .C2(new_n440), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n340), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT32), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n189), .A2(new_n190), .A3(G210), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(KEYINPUT27), .ZN(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT26), .B(G101), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n448), .B(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(KEYINPUT65), .B1(new_n346), .B2(new_n351), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT11), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n452), .B1(new_n268), .B2(G137), .ZN(new_n453));
  INV_X1    g267(.A(G137), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n454), .A2(KEYINPUT11), .A3(G134), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n268), .A2(G137), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n453), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G131), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n453), .A2(new_n455), .A3(new_n201), .A4(new_n456), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT65), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n342), .A2(new_n343), .A3(new_n345), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n349), .B1(new_n196), .B2(new_n230), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n461), .B(new_n462), .C1(new_n463), .C2(new_n347), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n451), .A2(new_n460), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n390), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n268), .A2(G137), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n454), .A2(G134), .ZN(new_n468));
  OAI21_X1  g282(.A(G131), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n459), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n470), .B1(new_n356), .B2(new_n359), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n465), .A2(new_n466), .A3(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(KEYINPUT28), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n458), .A2(new_n459), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n462), .B1(new_n463), .B2(new_n347), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n390), .B1(new_n477), .B2(new_n471), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n450), .B1(new_n474), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n465), .A2(KEYINPUT30), .A3(new_n472), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT30), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n481), .B1(new_n477), .B2(new_n471), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(new_n482), .A3(new_n390), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT66), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n480), .A2(new_n482), .A3(KEYINPUT66), .A4(new_n390), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n473), .A2(new_n450), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT67), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT67), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n473), .A2(new_n490), .A3(new_n450), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT31), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n487), .A2(KEYINPUT31), .A3(new_n492), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n479), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G472), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n187), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n446), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n479), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n487), .A2(KEYINPUT31), .A3(new_n492), .ZN(new_n502));
  AOI21_X1  g316(.A(KEYINPUT31), .B1(new_n487), .B2(new_n492), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n504), .A2(KEYINPUT32), .A3(new_n498), .A4(new_n187), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n465), .A2(new_n472), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n390), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n474), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n450), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT29), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(G902), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n450), .B1(new_n487), .B2(new_n473), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n474), .A2(new_n478), .A3(new_n450), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n510), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n512), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(G472), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n500), .A2(new_n505), .A3(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(KEYINPUT70), .A2(KEYINPUT25), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n520), .B(KEYINPUT68), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT22), .B(G137), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n521), .B(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT23), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n524), .B1(new_n396), .B2(G128), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n357), .A2(KEYINPUT23), .A3(G119), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n525), .B(new_n526), .C1(G119), .C2(new_n357), .ZN(new_n527));
  XNOR2_X1  g341(.A(G119), .B(G128), .ZN(new_n528));
  XOR2_X1   g342(.A(KEYINPUT24), .B(G110), .Z(new_n529));
  AOI22_X1  g343(.A1(new_n527), .A2(G110), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n530), .B1(new_n216), .B2(new_n217), .ZN(new_n531));
  OAI22_X1  g345(.A1(new_n527), .A2(G110), .B1(new_n528), .B2(new_n529), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(new_n215), .A3(new_n231), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n534), .A2(KEYINPUT69), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT69), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n536), .B1(new_n531), .B2(new_n533), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n523), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n523), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n539), .B1(new_n534), .B2(KEYINPUT69), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n519), .B1(new_n541), .B2(G902), .ZN(new_n542));
  INV_X1    g356(.A(new_n519), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n538), .A2(new_n187), .A3(new_n540), .A4(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(KEYINPUT70), .A2(KEYINPUT25), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n542), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n312), .B1(G234), .B2(new_n187), .ZN(new_n547));
  INV_X1    g361(.A(new_n541), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n547), .A2(G902), .ZN(new_n549));
  AOI22_X1  g363(.A1(new_n546), .A2(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(G221), .B1(new_n311), .B2(G902), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(G469), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n553), .A2(new_n187), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT10), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n342), .A2(new_n345), .A3(new_n358), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n342), .A2(new_n345), .ZN(new_n557));
  OAI21_X1  g371(.A(G128), .B1(new_n355), .B2(new_n353), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n408), .A2(new_n409), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n555), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n451), .A2(new_n381), .A3(new_n464), .A4(new_n391), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n408), .A2(new_n409), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n555), .B1(new_n356), .B2(new_n359), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n561), .A2(new_n562), .A3(new_n475), .A4(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT74), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n357), .B1(new_n348), .B2(KEYINPUT1), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n344), .B1(new_n288), .B2(G146), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n359), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n563), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g386(.A1(new_n572), .A2(new_n555), .B1(new_n563), .B2(new_n564), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n573), .A2(KEYINPUT74), .A3(new_n475), .A4(new_n562), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n568), .A2(new_n574), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n560), .A2(new_n356), .A3(new_n359), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n558), .A2(new_n557), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n560), .B1(new_n359), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n460), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT12), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g395(.A(KEYINPUT12), .B(new_n460), .C1(new_n576), .C2(new_n578), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n575), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(G110), .B(G140), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n190), .A2(G227), .ZN(new_n586));
  XOR2_X1   g400(.A(new_n585), .B(new_n586), .Z(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(KEYINPUT71), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n587), .B1(new_n568), .B2(new_n574), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n573), .A2(new_n562), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n460), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n584), .A2(new_n588), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n554), .B1(new_n592), .B2(G469), .ZN(new_n593));
  INV_X1    g407(.A(new_n587), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n575), .A2(new_n594), .A3(new_n583), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n594), .B1(new_n575), .B2(new_n591), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n553), .B(new_n187), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n552), .B1(new_n593), .B2(new_n597), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n445), .A2(new_n518), .A3(new_n550), .A4(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(G101), .ZN(G3));
  NOR2_X1   g414(.A1(new_n498), .A2(KEYINPUT89), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n601), .B1(new_n497), .B2(G902), .ZN(new_n602));
  INV_X1    g416(.A(new_n601), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n504), .A2(new_n187), .A3(new_n603), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n598), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT33), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n322), .A2(new_n606), .A3(new_n323), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n310), .A2(new_n313), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n321), .A2(KEYINPUT33), .A3(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n325), .A2(G902), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n607), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT90), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n607), .A2(KEYINPUT90), .A3(new_n609), .A4(new_n610), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n324), .A2(new_n325), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n264), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n341), .ZN(new_n618));
  INV_X1    g432(.A(new_n440), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n428), .A2(new_n438), .A3(new_n429), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n336), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n605), .A2(new_n550), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT34), .B(G104), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G6));
  INV_X1    g440(.A(KEYINPUT92), .ZN(new_n627));
  INV_X1    g441(.A(G475), .ZN(new_n628));
  AOI21_X1  g442(.A(G902), .B1(new_n245), .B2(new_n246), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n236), .A2(new_n241), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n631), .B1(new_n327), .B2(new_n338), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT91), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n263), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n235), .A2(new_n255), .A3(new_n240), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n635), .B(new_n260), .C1(new_n245), .C2(new_n240), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(KEYINPUT20), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n257), .A2(new_n249), .A3(new_n260), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n637), .A2(new_n638), .A3(KEYINPUT91), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n632), .A2(new_n634), .A3(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n627), .B1(new_n622), .B2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n441), .A2(new_n335), .ZN(new_n642));
  AND2_X1   g456(.A1(new_n639), .A2(new_n634), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n642), .A2(new_n643), .A3(KEYINPUT92), .A4(new_n632), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n645), .A2(new_n550), .A3(new_n605), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT35), .B(G107), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G9));
  NAND2_X1  g462(.A1(new_n546), .A2(new_n547), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n539), .A2(KEYINPUT36), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(new_n534), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n549), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n605), .A2(new_n445), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT37), .B(G110), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT93), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n654), .B(new_n656), .ZN(G12));
  INV_X1    g471(.A(new_n554), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n589), .A2(new_n591), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n575), .A2(new_n583), .ZN(new_n660));
  INV_X1    g474(.A(new_n588), .ZN(new_n661));
  OAI211_X1 g475(.A(G469), .B(new_n659), .C1(new_n660), .C2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n597), .A2(new_n658), .A3(new_n662), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n663), .A2(new_n551), .A3(new_n621), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n518), .A2(new_n664), .A3(new_n653), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n329), .B(KEYINPUT94), .Z(new_n666));
  OAI21_X1  g480(.A(new_n666), .B1(G900), .B2(new_n332), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n632), .A2(new_n639), .A3(new_n634), .A4(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT95), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n665), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G128), .ZN(G30));
  NAND3_X1  g486(.A1(new_n619), .A2(KEYINPUT38), .A3(new_n620), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT38), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n674), .B1(new_n439), .B2(new_n440), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n327), .A2(new_n338), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n264), .A2(new_n677), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n676), .A2(new_n678), .A3(new_n618), .ZN(new_n679));
  INV_X1    g493(.A(new_n653), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n450), .B1(new_n507), .B2(new_n473), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n681), .B1(new_n487), .B2(new_n492), .ZN(new_n682));
  OAI21_X1  g496(.A(G472), .B1(new_n682), .B2(G902), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n500), .A2(new_n505), .A3(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n679), .A2(new_n680), .A3(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT96), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n667), .B(KEYINPUT39), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n598), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT40), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n679), .A2(new_n684), .A3(KEYINPUT96), .A4(new_n680), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n687), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n196), .ZN(G45));
  NAND2_X1  g508(.A1(new_n611), .A2(new_n612), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n695), .A2(new_n615), .A3(new_n614), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(new_n264), .A3(new_n667), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n698), .A2(new_n518), .A3(new_n653), .A4(new_n664), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G146), .ZN(G48));
  AND2_X1   g514(.A1(new_n518), .A2(new_n550), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n575), .A2(new_n591), .ZN(new_n702));
  AOI22_X1  g516(.A1(new_n702), .A2(new_n587), .B1(new_n589), .B2(new_n583), .ZN(new_n703));
  OAI21_X1  g517(.A(G469), .B1(new_n703), .B2(G902), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(KEYINPUT97), .A3(new_n597), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT97), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n706), .B(G469), .C1(new_n703), .C2(G902), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n552), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n701), .A2(new_n623), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT41), .B(G113), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G15));
  NAND3_X1  g525(.A1(new_n701), .A2(new_n645), .A3(new_n708), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G116), .ZN(G18));
  AOI211_X1 g527(.A(new_n552), .B(new_n441), .C1(new_n705), .C2(new_n707), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n714), .A2(new_n518), .A3(new_n340), .A4(new_n653), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G119), .ZN(G21));
  NOR2_X1   g530(.A1(new_n622), .A2(new_n678), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n708), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n474), .A2(new_n507), .ZN(new_n719));
  AOI22_X1  g533(.A1(new_n495), .A2(new_n496), .B1(new_n509), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g534(.A(KEYINPUT98), .B1(new_n720), .B2(new_n499), .ZN(new_n721));
  OAI21_X1  g535(.A(G472), .B1(new_n497), .B2(G902), .ZN(new_n722));
  OAI22_X1  g536(.A1(new_n502), .A2(new_n503), .B1(new_n450), .B2(new_n508), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT98), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n723), .A2(new_n724), .A3(new_n498), .A4(new_n187), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n721), .A2(new_n722), .A3(new_n725), .A4(new_n550), .ZN(new_n726));
  OAI21_X1  g540(.A(KEYINPUT99), .B1(new_n718), .B2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n726), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT99), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n728), .A2(new_n729), .A3(new_n708), .A4(new_n717), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  AND4_X1   g546(.A1(new_n653), .A2(new_n721), .A3(new_n722), .A4(new_n725), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(new_n714), .A3(new_n698), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G125), .ZN(G27));
  NOR3_X1   g549(.A1(new_n439), .A2(new_n440), .A3(new_n618), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n663), .A2(new_n551), .A3(new_n736), .ZN(new_n737));
  AND2_X1   g551(.A1(KEYINPUT100), .A2(KEYINPUT42), .ZN(new_n738));
  NOR2_X1   g552(.A1(KEYINPUT100), .A2(KEYINPUT42), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n701), .A2(new_n698), .A3(new_n737), .A4(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n698), .A2(new_n518), .A3(new_n550), .A4(new_n737), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n738), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n201), .ZN(G33));
  AND3_X1   g559(.A1(new_n518), .A2(new_n737), .A3(new_n550), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n670), .ZN(new_n747));
  XNOR2_X1  g561(.A(KEYINPUT101), .B(G134), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(G36));
  AOI21_X1  g563(.A(new_n631), .B1(new_n637), .B2(new_n638), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n696), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT104), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n751), .A2(new_n752), .A3(KEYINPUT43), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n680), .B1(new_n602), .B2(new_n604), .ZN(new_n754));
  XNOR2_X1  g568(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n696), .A2(new_n750), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n753), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT106), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n758), .B1(new_n757), .B2(new_n759), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n736), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n753), .A2(new_n754), .A3(KEYINPUT44), .A4(new_n756), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT105), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n764), .B(new_n765), .ZN(new_n766));
  OAI21_X1  g580(.A(KEYINPUT107), .B1(new_n763), .B2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(new_n736), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n757), .A2(new_n759), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(KEYINPUT106), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n768), .B1(new_n770), .B2(new_n760), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT107), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n764), .B(KEYINPUT105), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n553), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n592), .A2(KEYINPUT45), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n554), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(KEYINPUT102), .B1(new_n779), .B2(KEYINPUT46), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n575), .A2(new_n591), .A3(new_n594), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n661), .B1(new_n575), .B2(new_n583), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n776), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n778), .A2(G469), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT46), .B1(new_n784), .B2(new_n658), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT102), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n784), .A2(KEYINPUT46), .A3(new_n658), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n780), .A2(new_n787), .A3(new_n597), .A4(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(new_n551), .A3(new_n688), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT103), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n789), .A2(KEYINPUT103), .A3(new_n551), .A4(new_n688), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n767), .A2(new_n774), .A3(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G137), .ZN(G39));
  NOR4_X1   g610(.A1(new_n518), .A2(new_n697), .A3(new_n550), .A4(new_n768), .ZN(new_n797));
  INV_X1    g611(.A(new_n787), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n597), .B(new_n788), .C1(new_n785), .C2(new_n786), .ZN(new_n799));
  OAI211_X1 g613(.A(KEYINPUT47), .B(new_n551), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT47), .B1(new_n789), .B2(new_n551), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n797), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G140), .ZN(G42));
  NAND2_X1  g618(.A1(new_n708), .A2(new_n736), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n753), .A2(new_n756), .ZN(new_n806));
  OR3_X1    g620(.A1(new_n806), .A2(KEYINPUT114), .A3(new_n666), .ZN(new_n807));
  OAI21_X1  g621(.A(KEYINPUT114), .B1(new_n806), .B2(new_n666), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n805), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n701), .ZN(new_n810));
  XOR2_X1   g624(.A(KEYINPUT118), .B(KEYINPUT48), .Z(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n809), .A2(KEYINPUT118), .A3(KEYINPUT48), .A4(new_n701), .ZN(new_n813));
  XOR2_X1   g627(.A(new_n328), .B(KEYINPUT117), .Z(new_n814));
  INV_X1    g628(.A(new_n684), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n815), .A2(new_n550), .A3(new_n329), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n816), .A2(new_n805), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n814), .B1(new_n817), .B2(new_n617), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n726), .B1(new_n807), .B2(new_n808), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n818), .B1(new_n819), .B2(new_n714), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n812), .A2(new_n813), .A3(new_n820), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n817), .A2(new_n264), .A3(new_n696), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n822), .B1(new_n809), .B2(new_n733), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT50), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n341), .B1(new_n824), .B2(new_n825), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n708), .A2(new_n676), .A3(new_n827), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n819), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n826), .B1(new_n819), .B2(new_n828), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n823), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n801), .A2(new_n802), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n551), .B1(new_n705), .B2(new_n707), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n736), .B(new_n819), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT51), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n821), .B1(new_n831), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n831), .A2(KEYINPUT116), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n838), .B(new_n823), .C1(new_n829), .C2(new_n830), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n837), .A2(new_n839), .A3(new_n834), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT51), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n836), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT110), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n518), .A2(new_n653), .ZN(new_n844));
  INV_X1    g658(.A(new_n667), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n677), .A2(new_n631), .A3(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n598), .A2(new_n846), .A3(new_n643), .A4(new_n736), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n843), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  AND4_X1   g662(.A1(new_n598), .A2(new_n643), .A3(new_n846), .A4(new_n736), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(KEYINPUT110), .A3(new_n518), .A4(new_n653), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n721), .A2(new_n722), .A3(new_n725), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n851), .A2(new_n697), .A3(new_n680), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n848), .A2(new_n850), .B1(new_n852), .B2(new_n737), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n853), .A2(new_n743), .A3(new_n741), .A4(new_n747), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT109), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n750), .A2(new_n855), .A3(new_n677), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n327), .A2(new_n338), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT109), .B1(new_n857), .B2(new_n264), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n617), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n442), .A2(new_n444), .A3(new_n336), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n605), .A2(new_n859), .A3(new_n550), .A4(new_n860), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n861), .A2(new_n599), .A3(new_n654), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n701), .B(new_n708), .C1(new_n645), .C2(new_n623), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n862), .A2(new_n731), .A3(new_n715), .A4(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n854), .A2(new_n864), .ZN(new_n865));
  XOR2_X1   g679(.A(new_n667), .B(KEYINPUT111), .Z(new_n866));
  AND2_X1   g680(.A1(new_n598), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n678), .A2(new_n441), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n867), .A2(new_n680), .A3(new_n684), .A4(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n671), .A2(new_n699), .A3(new_n734), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT52), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n665), .B1(new_n670), .B2(new_n698), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT52), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n872), .A2(new_n873), .A3(new_n734), .A4(new_n869), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n865), .A2(new_n875), .A3(KEYINPUT53), .ZN(new_n876));
  XOR2_X1   g690(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n877));
  NAND3_X1  g691(.A1(new_n861), .A2(new_n599), .A3(new_n654), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n878), .B1(new_n730), .B2(new_n727), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n863), .A2(new_n715), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n741), .A2(new_n743), .A3(new_n747), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n879), .A2(new_n880), .A3(new_n881), .A4(new_n853), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n871), .A2(new_n874), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n877), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n876), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n885), .A2(KEYINPUT54), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n865), .A2(new_n875), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT112), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n888), .A2(new_n889), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n891), .B1(new_n888), .B2(new_n877), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n890), .B1(new_n892), .B2(KEYINPUT112), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT54), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n842), .B(new_n887), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  OR2_X1    g709(.A1(G952), .A2(G953), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n550), .A2(new_n551), .A3(new_n341), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT108), .ZN(new_n899));
  AOI211_X1 g713(.A(new_n751), .B(new_n899), .C1(new_n673), .C2(new_n675), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n705), .A2(new_n707), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT49), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n900), .A2(new_n815), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n897), .A2(new_n903), .ZN(G75));
  INV_X1    g718(.A(new_n885), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n905), .A2(new_n187), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(G210), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT56), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n432), .A2(new_n437), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(new_n435), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT55), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n907), .A2(new_n908), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n911), .B1(new_n907), .B2(new_n908), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n190), .A2(G952), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(G51));
  XNOR2_X1  g729(.A(new_n554), .B(KEYINPUT57), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n905), .A2(new_n894), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n916), .B1(new_n917), .B2(new_n886), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n918), .B1(new_n596), .B2(new_n595), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n906), .A2(new_n778), .A3(new_n777), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n914), .B1(new_n919), .B2(new_n920), .ZN(G54));
  NAND3_X1  g735(.A1(new_n906), .A2(KEYINPUT58), .A3(G475), .ZN(new_n922));
  INV_X1    g736(.A(new_n257), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n922), .A2(new_n923), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n924), .A2(new_n925), .A3(new_n914), .ZN(G60));
  NAND2_X1  g740(.A1(new_n607), .A2(new_n609), .ZN(new_n927));
  NAND2_X1  g741(.A1(G478), .A2(G902), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT59), .Z(new_n929));
  NOR2_X1   g743(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n930), .B1(new_n917), .B2(new_n886), .ZN(new_n931));
  INV_X1    g745(.A(new_n914), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n887), .B1(new_n893), .B2(new_n894), .ZN(new_n934));
  INV_X1    g748(.A(new_n929), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n933), .B1(new_n936), .B2(new_n927), .ZN(G63));
  INV_X1    g751(.A(KEYINPUT119), .ZN(new_n938));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT60), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  AND4_X1   g755(.A1(new_n938), .A2(new_n885), .A3(new_n651), .A4(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n940), .B1(new_n876), .B2(new_n884), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n938), .B1(new_n943), .B2(new_n651), .ZN(new_n944));
  OAI21_X1  g758(.A(KEYINPUT120), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n885), .A2(new_n651), .A3(new_n941), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(KEYINPUT119), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT120), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n943), .A2(new_n938), .A3(new_n651), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n943), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n914), .B1(new_n951), .B2(new_n541), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n945), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT61), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n942), .A2(new_n944), .ZN(new_n956));
  OAI211_X1 g770(.A(KEYINPUT61), .B(new_n932), .C1(new_n943), .C2(new_n548), .ZN(new_n957));
  OAI21_X1  g771(.A(KEYINPUT121), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n957), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT121), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n959), .B(new_n960), .C1(new_n942), .C2(new_n944), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n955), .A2(new_n962), .ZN(G66));
  OAI21_X1  g777(.A(G953), .B1(new_n334), .B2(new_n363), .ZN(new_n964));
  INV_X1    g778(.A(new_n864), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n964), .B1(new_n965), .B2(G953), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n909), .B1(G898), .B2(new_n190), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(G69));
  AOI21_X1  g782(.A(new_n190), .B1(G227), .B2(G900), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT62), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n693), .A2(new_n970), .A3(new_n734), .A4(new_n872), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n746), .A2(new_n688), .A3(new_n859), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(KEYINPUT123), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT123), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n746), .A2(new_n974), .A3(new_n688), .A4(new_n859), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n803), .A2(new_n971), .A3(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n693), .A2(new_n734), .A3(new_n872), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(KEYINPUT62), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT122), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n978), .A2(KEYINPUT122), .A3(KEYINPUT62), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n977), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n795), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n190), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT124), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n480), .A2(new_n482), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n252), .A2(new_n253), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n987), .B(new_n988), .Z(new_n989));
  NAND3_X1  g803(.A1(new_n985), .A2(new_n986), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(G953), .B1(new_n983), .B2(new_n795), .ZN(new_n991));
  INV_X1    g805(.A(new_n989), .ZN(new_n992));
  OAI21_X1  g806(.A(KEYINPUT124), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n190), .A2(G900), .ZN(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n872), .A2(new_n734), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n803), .A2(new_n881), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n701), .A2(new_n868), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n999), .B1(new_n792), .B2(new_n793), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n795), .A2(new_n1001), .ZN(new_n1002));
  OAI211_X1 g816(.A(KEYINPUT125), .B(new_n996), .C1(new_n1002), .C2(G953), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT125), .ZN(new_n1004));
  AOI21_X1  g818(.A(G953), .B1(new_n795), .B2(new_n1001), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1004), .B1(new_n1005), .B2(new_n995), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n1003), .A2(new_n1006), .A3(new_n992), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n969), .B1(new_n994), .B2(new_n1007), .ZN(new_n1008));
  AND4_X1   g822(.A1(new_n1007), .A2(new_n993), .A3(new_n990), .A4(new_n969), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1008), .A2(new_n1009), .ZN(G72));
  NAND2_X1  g824(.A1(new_n487), .A2(new_n473), .ZN(new_n1011));
  NAND2_X1  g825(.A1(G472), .A2(G902), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT63), .Z(new_n1013));
  OAI21_X1  g827(.A(new_n1013), .B1(new_n984), .B2(new_n864), .ZN(new_n1014));
  AND2_X1   g828(.A1(new_n1014), .A2(KEYINPUT126), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n1014), .A2(KEYINPUT126), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n450), .B(new_n1011), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n1011), .A2(new_n450), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT127), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1002), .A2(new_n965), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1019), .B1(new_n1020), .B2(new_n1013), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1013), .ZN(new_n1022));
  AOI211_X1 g836(.A(KEYINPUT127), .B(new_n1022), .C1(new_n1002), .C2(new_n965), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1018), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g838(.A(new_n893), .ZN(new_n1025));
  INV_X1    g839(.A(new_n513), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1022), .B1(new_n1026), .B2(new_n493), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n914), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  AND3_X1   g842(.A1(new_n1017), .A2(new_n1024), .A3(new_n1028), .ZN(G57));
endmodule


