//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 0 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(new_n202));
  XOR2_X1   g0002(.A(new_n202), .B(KEYINPUT64), .Z(G355));
  NAND2_X1  g0003(.A1(G1), .A2(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G13), .ZN(new_n205));
  OAI211_X1 g0005(.A(new_n205), .B(G250), .C1(G257), .C2(G264), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT0), .Z(new_n207));
  INV_X1    g0007(.A(G58), .ZN(new_n208));
  INV_X1    g0008(.A(G232), .ZN(new_n209));
  INV_X1    g0009(.A(G77), .ZN(new_n210));
  INV_X1    g0010(.A(G244), .ZN(new_n211));
  OAI22_X1  g0011(.A1(new_n208), .A2(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G50), .ZN(new_n213));
  INV_X1    g0013(.A(G226), .ZN(new_n214));
  INV_X1    g0014(.A(G116), .ZN(new_n215));
  INV_X1    g0015(.A(G270), .ZN(new_n216));
  OAI22_X1  g0016(.A1(new_n213), .A2(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G87), .A2(G250), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G97), .A2(G257), .ZN(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT65), .B(G238), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(G68), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G107), .ZN(new_n224));
  INV_X1    g0024(.A(G264), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n204), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT66), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(G68), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n208), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n234), .A2(G50), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  AOI211_X1 g0036(.A(new_n207), .B(new_n229), .C1(new_n232), .C2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G264), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(new_n216), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT67), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G232), .ZN(new_n243));
  XOR2_X1   g0043(.A(G238), .B(G244), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT68), .ZN(new_n250));
  XOR2_X1   g0050(.A(G68), .B(G77), .Z(new_n251));
  XOR2_X1   g0051(.A(G50), .B(G58), .Z(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  INV_X1    g0054(.A(KEYINPUT14), .ZN(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT69), .B(G41), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n256), .B(G274), .C1(new_n257), .C2(G45), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT70), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n258), .B(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n230), .B1(G33), .B2(G41), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n256), .B1(G41), .B2(G45), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G238), .ZN(new_n266));
  XNOR2_X1  g0066(.A(new_n261), .B(KEYINPUT72), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT3), .B(G33), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(G232), .A3(G1698), .ZN(new_n269));
  INV_X1    g0069(.A(G1698), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n269), .B1(new_n271), .B2(new_n214), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  INV_X1    g0073(.A(G97), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n267), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n260), .A2(new_n266), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT13), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT13), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n260), .A2(new_n276), .A3(new_n279), .A4(new_n266), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n255), .B1(new_n281), .B2(G169), .ZN(new_n282));
  INV_X1    g0082(.A(G169), .ZN(new_n283));
  AOI211_X1 g0083(.A(KEYINPUT14), .B(new_n283), .C1(new_n278), .C2(new_n280), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G179), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n230), .B1(new_n204), .B2(new_n273), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT73), .ZN(new_n291));
  XNOR2_X1  g0091(.A(new_n290), .B(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n233), .A2(G20), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n231), .A2(G33), .ZN(new_n294));
  NOR2_X1   g0094(.A1(G20), .A2(G33), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  OAI221_X1 g0096(.A(new_n293), .B1(new_n294), .B2(new_n210), .C1(new_n296), .C2(new_n213), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n298), .B(KEYINPUT11), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n290), .B(KEYINPUT73), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n256), .A2(G20), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n299), .B1(new_n233), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G13), .ZN(new_n304));
  NOR3_X1   g0104(.A1(new_n304), .A2(new_n231), .A3(G1), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n305), .A2(KEYINPUT79), .A3(new_n233), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT12), .ZN(new_n307));
  AOI21_X1  g0107(.A(KEYINPUT79), .B1(new_n305), .B2(new_n233), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n307), .B(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n303), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n289), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n281), .A2(G200), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n278), .A2(G190), .A3(new_n280), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n313), .A2(new_n310), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n268), .A2(G1698), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n317), .B(KEYINPUT71), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n318), .A2(G223), .ZN(new_n319));
  INV_X1    g0119(.A(G222), .ZN(new_n320));
  OAI22_X1  g0120(.A1(new_n271), .A2(new_n320), .B1(new_n210), .B2(new_n268), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n267), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  OR2_X1    g0122(.A1(new_n258), .A2(new_n259), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n258), .A2(new_n259), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n323), .A2(new_n324), .B1(G226), .B2(new_n265), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n322), .A2(G190), .A3(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(G20), .B1(new_n234), .B2(G50), .ZN(new_n327));
  INV_X1    g0127(.A(G150), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT8), .B(G58), .ZN(new_n329));
  OAI221_X1 g0129(.A(new_n327), .B1(new_n328), .B2(new_n296), .C1(new_n329), .C2(new_n294), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n292), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n300), .A2(G50), .A3(new_n301), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n305), .A2(new_n213), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n334), .B(KEYINPUT9), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n326), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G200), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n337), .B1(new_n322), .B2(new_n325), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT78), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n339), .A2(new_n340), .A3(KEYINPUT10), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(KEYINPUT10), .ZN(new_n342));
  OR2_X1    g0142(.A1(new_n340), .A2(KEYINPUT10), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n342), .B(new_n343), .C1(new_n336), .C2(new_n338), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n322), .A2(new_n325), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n283), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n346), .B(new_n334), .C1(G179), .C2(new_n345), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n341), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n316), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(G58), .A2(G68), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT80), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT80), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n352), .A2(G58), .A3(G68), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n351), .A2(new_n353), .A3(new_n234), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G20), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n295), .A2(G159), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT81), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n295), .A2(KEYINPUT81), .A3(G159), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT82), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT7), .ZN(new_n363));
  NOR3_X1   g0163(.A1(new_n268), .A2(new_n363), .A3(G20), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n273), .A2(KEYINPUT3), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT3), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(G33), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(KEYINPUT7), .B1(new_n368), .B2(new_n231), .ZN(new_n369));
  OAI21_X1  g0169(.A(G68), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT82), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n355), .A2(new_n360), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n362), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT16), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n362), .A2(KEYINPUT16), .A3(new_n370), .A4(new_n372), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n375), .A2(new_n292), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n329), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n302), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(new_n378), .B2(new_n305), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n365), .A2(new_n367), .A3(G226), .A4(G1698), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT83), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n268), .A2(KEYINPUT83), .A3(G226), .A4(G1698), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n365), .A2(new_n367), .A3(G223), .A4(new_n270), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G33), .A2(G87), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(KEYINPUT84), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n388), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT84), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n390), .A2(new_n391), .A3(new_n383), .A4(new_n384), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n389), .A2(new_n267), .A3(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(G190), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n394), .A2(KEYINPUT85), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(KEYINPUT85), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n323), .A2(new_n324), .B1(G232), .B2(new_n265), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n393), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(G200), .B1(new_n393), .B2(new_n398), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n377), .B(new_n380), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT17), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n393), .A2(new_n398), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n337), .ZN(new_n405));
  INV_X1    g0205(.A(new_n397), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n405), .B1(new_n406), .B2(new_n404), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n407), .A2(KEYINPUT17), .A3(new_n380), .A4(new_n377), .ZN(new_n408));
  AND3_X1   g0208(.A1(new_n393), .A2(new_n286), .A3(new_n398), .ZN(new_n409));
  AOI21_X1  g0209(.A(G169), .B1(new_n393), .B2(new_n398), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n377), .A2(new_n380), .ZN(new_n412));
  AND3_X1   g0212(.A1(new_n411), .A2(new_n412), .A3(KEYINPUT18), .ZN(new_n413));
  AOI21_X1  g0213(.A(KEYINPUT18), .B1(new_n411), .B2(new_n412), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n403), .B(new_n408), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n378), .A2(new_n295), .B1(G20), .B2(G77), .ZN(new_n417));
  XNOR2_X1  g0217(.A(KEYINPUT15), .B(G87), .ZN(new_n418));
  XNOR2_X1  g0218(.A(new_n418), .B(KEYINPUT74), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n417), .B1(new_n419), .B2(new_n294), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n420), .A2(new_n292), .B1(new_n210), .B2(new_n305), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT75), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n302), .B2(new_n210), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n300), .A2(KEYINPUT75), .A3(G77), .A4(new_n301), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n421), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT76), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n421), .A2(KEYINPUT76), .A3(new_n423), .A4(new_n424), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n267), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n268), .A2(new_n224), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(new_n318), .B2(new_n221), .ZN(new_n432));
  NOR3_X1   g0232(.A1(new_n368), .A2(new_n209), .A3(G1698), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n430), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n260), .B1(new_n211), .B2(new_n264), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n283), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n436), .ZN(new_n438));
  AOI211_X1 g0238(.A(new_n431), .B(new_n433), .C1(new_n318), .C2(new_n221), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n438), .B(new_n286), .C1(new_n439), .C2(new_n430), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n429), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT77), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n438), .B(G190), .C1(new_n439), .C2(new_n430), .ZN(new_n443));
  OAI21_X1  g0243(.A(G200), .B1(new_n435), .B2(new_n436), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n443), .A2(new_n444), .A3(new_n427), .A4(new_n428), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n441), .A2(new_n442), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n442), .B1(new_n441), .B2(new_n445), .ZN(new_n447));
  OR2_X1    g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n349), .A2(KEYINPUT86), .A3(new_n416), .A4(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT86), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n341), .A2(new_n344), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n451), .A2(new_n312), .A3(new_n315), .A4(new_n347), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n416), .B1(new_n446), .B2(new_n447), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n450), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n268), .A2(new_n231), .A3(G87), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT22), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT22), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n268), .A2(new_n459), .A3(new_n231), .A4(G87), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n231), .A2(G33), .A3(G116), .ZN(new_n462));
  XOR2_X1   g0262(.A(new_n462), .B(KEYINPUT93), .Z(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n231), .A2(G107), .ZN(new_n465));
  XNOR2_X1  g0265(.A(new_n465), .B(KEYINPUT23), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n461), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT24), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n463), .B1(new_n458), .B2(new_n460), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT24), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n469), .A2(new_n470), .A3(new_n466), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n292), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n273), .A2(G1), .ZN(new_n474));
  OR2_X1    g0274(.A1(new_n474), .A2(KEYINPUT88), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n305), .B1(KEYINPUT88), .B2(new_n474), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n300), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n477), .A2(new_n224), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n304), .A2(G1), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n465), .ZN(new_n480));
  XNOR2_X1  g0280(.A(new_n480), .B(KEYINPUT25), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n473), .A2(KEYINPUT94), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT94), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n300), .B1(new_n468), .B2(new_n471), .ZN(new_n485));
  INV_X1    g0285(.A(new_n482), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n268), .B1(G250), .B2(G1698), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n270), .A2(G257), .ZN(new_n489));
  INV_X1    g0289(.A(G294), .ZN(new_n490));
  OAI22_X1  g0290(.A1(new_n488), .A2(new_n489), .B1(new_n273), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n267), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT5), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n257), .A2(new_n493), .ZN(new_n494));
  OR2_X1    g0294(.A1(new_n493), .A2(G41), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n494), .A2(new_n256), .A3(G45), .A4(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n496), .A2(G264), .A3(new_n262), .ZN(new_n497));
  OR2_X1    g0297(.A1(new_n495), .A2(KEYINPUT89), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n256), .A2(G45), .A3(G274), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n495), .A2(KEYINPUT89), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n498), .A2(new_n494), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n492), .A2(new_n497), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G169), .ZN(new_n503));
  OR2_X1    g0303(.A1(new_n502), .A2(new_n286), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n483), .A2(new_n487), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n502), .A2(G200), .ZN(new_n506));
  OR2_X1    g0306(.A1(new_n502), .A2(new_n394), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n473), .A2(new_n482), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n305), .A2(new_n274), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(G107), .B1(new_n364), .B2(new_n369), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT87), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n224), .A2(KEYINPUT6), .A3(G97), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n274), .A2(new_n224), .ZN(new_n517));
  NOR2_X1   g0317(.A1(G97), .A2(G107), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n516), .B1(new_n519), .B2(KEYINPUT6), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n520), .A2(G20), .B1(G77), .B2(new_n295), .ZN(new_n521));
  OAI211_X1 g0321(.A(KEYINPUT87), .B(G107), .C1(new_n364), .C2(new_n369), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n515), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n512), .B1(new_n523), .B2(new_n292), .ZN(new_n524));
  INV_X1    g0324(.A(new_n477), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G97), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n268), .A2(G244), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT4), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n528), .A2(new_n529), .B1(G33), .B2(G283), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n268), .A2(KEYINPUT4), .A3(G244), .A4(new_n270), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n529), .B1(new_n268), .B2(G250), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n530), .B(new_n531), .C1(new_n270), .C2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n267), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n496), .A2(G257), .A3(new_n262), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n534), .A2(new_n535), .A3(new_n501), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n283), .ZN(new_n537));
  INV_X1    g0337(.A(new_n501), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(new_n533), .B2(new_n267), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n539), .A2(new_n286), .A3(new_n535), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n527), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n536), .A2(G200), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n539), .A2(G190), .A3(new_n535), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n542), .A2(new_n524), .A3(new_n526), .A4(new_n543), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT21), .ZN(new_n546));
  AOI21_X1  g0346(.A(G20), .B1(G33), .B2(G283), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(G33), .B2(new_n274), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n548), .B(new_n290), .C1(new_n231), .C2(G116), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT20), .ZN(new_n550));
  XNOR2_X1  g0350(.A(new_n549), .B(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n305), .A2(new_n215), .ZN(new_n552));
  XOR2_X1   g0352(.A(new_n552), .B(KEYINPUT91), .Z(new_n553));
  NAND4_X1  g0353(.A1(new_n300), .A2(G116), .A3(new_n475), .A4(new_n476), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n551), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(G303), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n368), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n270), .A2(G257), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n268), .B(new_n559), .C1(new_n225), .C2(new_n270), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n267), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n496), .A2(G270), .A3(new_n262), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n561), .A2(new_n562), .A3(new_n501), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G169), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n546), .B1(new_n556), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n563), .A2(new_n286), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n555), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n555), .A2(KEYINPUT21), .A3(G169), .A4(new_n563), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n565), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT92), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n563), .A2(G200), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n556), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n570), .B1(new_n556), .B2(new_n571), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OR2_X1    g0374(.A1(new_n563), .A2(new_n397), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n569), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n211), .A2(G1698), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(G238), .B2(G1698), .ZN(new_n578));
  OAI22_X1  g0378(.A1(new_n578), .A2(new_n368), .B1(new_n273), .B2(new_n215), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n499), .B1(new_n267), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n256), .A2(G45), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n262), .A2(G250), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(G200), .ZN(new_n584));
  OR3_X1    g0384(.A1(new_n583), .A2(KEYINPUT90), .A3(new_n394), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n525), .A2(G87), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT19), .ZN(new_n587));
  INV_X1    g0387(.A(G87), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n587), .B1(new_n518), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(G20), .B2(new_n275), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n268), .A2(new_n231), .A3(G68), .ZN(new_n591));
  NOR3_X1   g0391(.A1(new_n273), .A2(new_n274), .A3(G20), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n590), .B(new_n591), .C1(KEYINPUT19), .C2(new_n592), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n593), .A2(new_n292), .B1(new_n419), .B2(new_n305), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n586), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(KEYINPUT90), .B1(new_n583), .B2(new_n394), .ZN(new_n596));
  AND4_X1   g0396(.A1(new_n584), .A2(new_n585), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n583), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n286), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n583), .A2(new_n283), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n594), .B1(new_n419), .B2(new_n477), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n597), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n510), .A2(new_n545), .A3(new_n576), .A4(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n456), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g0406(.A(new_n606), .B(KEYINPUT95), .Z(G372));
  INV_X1    g0407(.A(new_n347), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n413), .A2(new_n414), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n315), .ZN(new_n611));
  OR2_X1    g0411(.A1(new_n611), .A2(new_n441), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n312), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT96), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n612), .A2(new_n312), .A3(KEYINPUT96), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n408), .A2(new_n403), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n610), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n608), .B1(new_n619), .B2(new_n451), .ZN(new_n620));
  INV_X1    g0420(.A(new_n541), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n598), .A2(G190), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n595), .A2(new_n622), .A3(new_n584), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n623), .A2(new_n602), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT26), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n621), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n541), .A2(new_n544), .A3(new_n508), .A4(new_n623), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n473), .A2(new_n482), .B1(new_n504), .B2(new_n503), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n569), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n626), .B(new_n602), .C1(new_n627), .C2(new_n629), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n597), .A2(new_n541), .A3(new_n603), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n631), .A2(new_n625), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n620), .B1(new_n456), .B2(new_n634), .ZN(G369));
  NAND2_X1  g0435(.A1(new_n479), .A2(new_n231), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n636), .A2(KEYINPUT27), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(KEYINPUT27), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(new_n638), .A3(G213), .ZN(new_n639));
  INV_X1    g0439(.A(G343), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n576), .B1(new_n556), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n569), .A2(new_n555), .A3(new_n641), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(KEYINPUT97), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT97), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n643), .A2(new_n647), .A3(new_n644), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n483), .A2(new_n487), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n510), .B1(new_n651), .B2(new_n642), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n504), .A2(new_n503), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n652), .B1(new_n654), .B2(new_n642), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n649), .A2(G330), .A3(new_n655), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(KEYINPUT98), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(KEYINPUT98), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n569), .A2(new_n642), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n510), .A2(new_n661), .B1(new_n628), .B2(new_n642), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n659), .A2(new_n662), .ZN(G399));
  INV_X1    g0463(.A(new_n205), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(new_n257), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n518), .A2(new_n588), .A3(new_n215), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n665), .A2(new_n256), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n667), .B1(new_n236), .B2(new_n665), .ZN(new_n668));
  XNOR2_X1  g0468(.A(KEYINPUT99), .B(KEYINPUT28), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n668), .B(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n642), .B1(new_n630), .B2(new_n632), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT103), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OAI211_X1 g0473(.A(KEYINPUT103), .B(new_n642), .C1(new_n630), .C2(new_n632), .ZN(new_n674));
  XNOR2_X1  g0474(.A(KEYINPUT104), .B(KEYINPUT29), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n623), .A2(new_n602), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n677), .A2(new_n541), .A3(new_n625), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT105), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n603), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n621), .A2(new_n624), .A3(KEYINPUT26), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n681), .B(KEYINPUT105), .C1(new_n631), .C2(KEYINPUT26), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT106), .ZN(new_n683));
  INV_X1    g0483(.A(new_n569), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n654), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(KEYINPUT106), .B1(new_n505), .B2(new_n569), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n680), .B(new_n682), .C1(new_n687), .C2(new_n627), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n688), .A2(KEYINPUT29), .A3(new_n642), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n536), .A2(new_n502), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT102), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n536), .A2(KEYINPUT102), .A3(new_n502), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n692), .A2(new_n286), .A3(new_n563), .A4(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(new_n598), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n580), .A2(new_n492), .A3(new_n497), .A4(new_n582), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(KEYINPUT100), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n566), .ZN(new_n698));
  OAI211_X1 g0498(.A(new_n539), .B(new_n535), .C1(new_n696), .C2(KEYINPUT100), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT101), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(KEYINPUT30), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT30), .ZN(new_n702));
  OAI211_X1 g0502(.A(KEYINPUT101), .B(new_n702), .C1(new_n698), .C2(new_n699), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n641), .B1(new_n695), .B2(new_n704), .ZN(new_n705));
  OAI211_X1 g0505(.A(KEYINPUT31), .B(new_n705), .C1(new_n605), .C2(new_n641), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n705), .A2(KEYINPUT31), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI22_X1  g0508(.A1(new_n676), .A2(new_n689), .B1(new_n708), .B2(G330), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n670), .B1(new_n709), .B2(G1), .ZN(G364));
  INV_X1    g0510(.A(new_n665), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n304), .A2(G20), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G45), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n711), .A2(G1), .A3(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n649), .ZN(new_n715));
  NOR2_X1   g0515(.A1(G13), .A2(G33), .ZN(new_n716));
  XOR2_X1   g0516(.A(new_n716), .B(KEYINPUT107), .Z(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(G20), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n714), .B1(new_n715), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n230), .B1(G20), .B2(new_n283), .ZN(new_n721));
  NOR2_X1   g0521(.A1(G179), .A2(G200), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT108), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(new_n394), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n231), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT109), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(new_n274), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n231), .A2(G179), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(G190), .A3(G200), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(new_n588), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n231), .A2(new_n286), .A3(G200), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n394), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AOI211_X1 g0534(.A(new_n368), .B(new_n731), .C1(G77), .C2(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n729), .A2(new_n394), .A3(G200), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n735), .B1(new_n224), .B2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT32), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n723), .A2(new_n231), .A3(G190), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(G159), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n738), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n739), .A2(KEYINPUT32), .A3(G159), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n737), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n406), .A2(new_n732), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n231), .A2(new_n286), .A3(new_n337), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n394), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n746), .A2(G58), .B1(new_n749), .B2(G68), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n728), .A2(new_n744), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n406), .A2(new_n747), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n751), .B1(G50), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g0554(.A(KEYINPUT110), .B(G326), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n753), .A2(new_n755), .B1(new_n739), .B2(G329), .ZN(new_n756));
  INV_X1    g0556(.A(G283), .ZN(new_n757));
  OAI221_X1 g0557(.A(new_n756), .B1(new_n757), .B2(new_n736), .C1(new_n557), .C2(new_n730), .ZN(new_n758));
  INV_X1    g0558(.A(G311), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n733), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n725), .A2(new_n490), .ZN(new_n761));
  INV_X1    g0561(.A(G317), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n748), .B1(KEYINPUT33), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(KEYINPUT33), .B2(new_n762), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n746), .A2(G322), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n764), .A2(new_n765), .A3(new_n368), .ZN(new_n766));
  NOR4_X1   g0566(.A1(new_n758), .A2(new_n760), .A3(new_n761), .A4(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n721), .B1(new_n754), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n253), .A2(G45), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n664), .A2(new_n268), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n769), .B(new_n770), .C1(G45), .C2(new_n235), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n664), .A2(new_n368), .ZN(new_n772));
  NAND2_X1  g0572(.A1(G355), .A2(new_n772), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n771), .B(new_n773), .C1(G116), .C2(new_n205), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n719), .A2(new_n721), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n720), .A2(new_n768), .A3(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n714), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n778), .B1(new_n649), .B2(G330), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(G330), .B2(new_n649), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n777), .A2(new_n780), .ZN(G396));
  INV_X1    g0581(.A(new_n721), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n746), .A2(G143), .B1(G159), .B2(new_n734), .ZN(new_n783));
  INV_X1    g0583(.A(G137), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n783), .B1(new_n784), .B2(new_n752), .C1(new_n328), .C2(new_n748), .ZN(new_n785));
  XOR2_X1   g0585(.A(new_n785), .B(KEYINPUT34), .Z(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n368), .ZN(new_n787));
  INV_X1    g0587(.A(new_n725), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G58), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n739), .A2(G132), .ZN(new_n790));
  INV_X1    g0590(.A(new_n730), .ZN(new_n791));
  INV_X1    g0591(.A(new_n736), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n791), .A2(G50), .B1(new_n792), .B2(G68), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n787), .A2(new_n789), .A3(new_n790), .A4(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n728), .B1(new_n490), .B2(new_n745), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n795), .B1(G303), .B2(new_n753), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n734), .A2(G116), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n368), .B1(new_n730), .B2(new_n224), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n798), .B(KEYINPUT112), .Z(new_n799));
  OAI22_X1  g0599(.A1(new_n740), .A2(new_n759), .B1(new_n588), .B2(new_n736), .ZN(new_n800));
  OR2_X1    g0600(.A1(new_n749), .A2(KEYINPUT111), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n749), .A2(KEYINPUT111), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n800), .B1(G283), .B2(new_n803), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n796), .A2(new_n797), .A3(new_n799), .A4(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n782), .B1(new_n794), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n429), .A2(new_n437), .A3(new_n440), .A4(new_n642), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n429), .A2(new_n641), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n445), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n808), .B1(new_n441), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n718), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n721), .A2(new_n716), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(G77), .ZN(new_n815));
  NOR4_X1   g0615(.A1(new_n806), .A2(new_n812), .A3(new_n714), .A4(new_n815), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n811), .B(new_n642), .C1(new_n630), .C2(new_n632), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n673), .A2(new_n674), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n810), .A2(new_n441), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n807), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n818), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n708), .A2(G330), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n822), .B(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n816), .B1(new_n824), .B2(new_n714), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G384));
  INV_X1    g0626(.A(KEYINPUT115), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT37), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n411), .A2(new_n412), .ZN(new_n829));
  INV_X1    g0629(.A(new_n639), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n412), .A2(new_n830), .ZN(new_n831));
  AND4_X1   g0631(.A1(new_n828), .A2(new_n829), .A3(new_n401), .A4(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n412), .B1(new_n411), .B2(new_n830), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n828), .B1(new_n833), .B2(new_n401), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n827), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n831), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n415), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n404), .A2(new_n283), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n393), .A2(new_n286), .A3(new_n398), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n840), .A2(new_n639), .B1(new_n380), .B2(new_n377), .ZN(new_n841));
  INV_X1    g0641(.A(new_n401), .ZN(new_n842));
  OAI21_X1  g0642(.A(KEYINPUT37), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n833), .A2(new_n828), .A3(new_n401), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n843), .A2(KEYINPUT115), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n835), .A2(new_n837), .A3(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT38), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT116), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n843), .A2(new_n844), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT114), .ZN(new_n852));
  AND3_X1   g0652(.A1(new_n415), .A2(new_n852), .A3(new_n836), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n852), .B1(new_n415), .B2(new_n836), .ZN(new_n854));
  OAI211_X1 g0654(.A(KEYINPUT38), .B(new_n851), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n846), .A2(KEYINPUT116), .A3(new_n847), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n850), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT39), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n312), .A2(new_n641), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n851), .B1(new_n853), .B2(new_n854), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n847), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n862), .A2(KEYINPUT39), .A3(new_n855), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n859), .A2(new_n860), .A3(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n311), .B(new_n641), .C1(new_n289), .C2(new_n611), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n311), .A2(new_n641), .ZN(new_n866));
  NOR3_X1   g0666(.A1(new_n282), .A2(new_n284), .A3(new_n287), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n315), .B(new_n866), .C1(new_n867), .C2(new_n310), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n817), .B2(new_n807), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n862), .A2(new_n855), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n871), .A2(new_n872), .B1(new_n609), .B2(new_n639), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n864), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n455), .A2(new_n676), .A3(new_n689), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n620), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n874), .B(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n708), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n456), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n821), .B1(new_n865), .B2(new_n868), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n706), .A2(new_n707), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n837), .A2(KEYINPUT114), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n415), .A2(new_n852), .A3(new_n836), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT38), .B1(new_n885), .B2(new_n851), .ZN(new_n886));
  INV_X1    g0686(.A(new_n855), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n882), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT40), .ZN(new_n889));
  AND4_X1   g0689(.A1(KEYINPUT40), .A2(new_n706), .A3(new_n707), .A4(new_n881), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n888), .A2(new_n889), .B1(new_n857), .B2(new_n890), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n880), .B(new_n891), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n892), .A2(G330), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n877), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n877), .A2(new_n893), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n894), .B(new_n895), .C1(new_n256), .C2(new_n712), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n215), .B1(new_n520), .B2(KEYINPUT35), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n897), .B(new_n232), .C1(KEYINPUT35), .C2(new_n520), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n898), .B(KEYINPUT36), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n236), .A2(G77), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n351), .A2(new_n353), .ZN(new_n901));
  OAI22_X1  g0701(.A1(new_n900), .A2(new_n901), .B1(G50), .B2(new_n233), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n902), .A2(G1), .A3(new_n304), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n903), .B(KEYINPUT113), .Z(new_n904));
  NAND3_X1  g0704(.A1(new_n896), .A2(new_n899), .A3(new_n904), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT117), .ZN(G367));
  AOI22_X1  g0706(.A1(new_n803), .A2(G159), .B1(G50), .B2(new_n734), .ZN(new_n907));
  OAI221_X1 g0707(.A(new_n907), .B1(new_n210), .B2(new_n736), .C1(new_n784), .C2(new_n740), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n726), .A2(new_n233), .ZN(new_n909));
  OAI22_X1  g0709(.A1(new_n745), .A2(new_n328), .B1(new_n208), .B2(new_n730), .ZN(new_n910));
  NOR3_X1   g0710(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(G143), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n911), .B(new_n268), .C1(new_n912), .C2(new_n752), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n791), .A2(KEYINPUT46), .A3(G116), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n368), .B(new_n914), .C1(new_n725), .C2(new_n224), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n733), .A2(new_n757), .B1(new_n736), .B2(new_n274), .ZN(new_n916));
  AOI21_X1  g0716(.A(KEYINPUT46), .B1(new_n791), .B2(G116), .ZN(new_n917));
  NOR3_X1   g0717(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AOI22_X1  g0718(.A1(G303), .A2(new_n746), .B1(new_n753), .B2(G311), .ZN(new_n919));
  INV_X1    g0719(.A(new_n803), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n918), .B(new_n919), .C1(new_n490), .C2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n740), .A2(new_n762), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n913), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT47), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n721), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n595), .A2(new_n642), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n624), .A2(new_n926), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n926), .A2(new_n602), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n927), .A2(new_n719), .A3(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n770), .ZN(new_n930));
  OAI221_X1 g0730(.A(new_n775), .B1(new_n205), .B2(new_n419), .C1(new_n240), .C2(new_n930), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n925), .A2(new_n778), .A3(new_n929), .A4(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n510), .A2(new_n545), .A3(new_n661), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n933), .B(KEYINPUT42), .Z(new_n934));
  NAND2_X1  g0734(.A1(new_n927), .A2(new_n928), .ZN(new_n935));
  XOR2_X1   g0735(.A(KEYINPUT118), .B(KEYINPUT43), .Z(new_n936));
  NOR2_X1   g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n527), .A2(new_n641), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n545), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n541), .B1(new_n939), .B2(new_n654), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n642), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n934), .A2(new_n937), .A3(new_n941), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT119), .Z(new_n943));
  NAND2_X1  g0743(.A1(new_n934), .A2(new_n941), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n937), .B1(KEYINPUT43), .B2(new_n935), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(KEYINPUT120), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT120), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n943), .A2(new_n949), .A3(new_n946), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n659), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n621), .A2(new_n641), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n939), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n951), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n948), .A2(new_n952), .A3(new_n954), .A4(new_n950), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n713), .A2(G1), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n662), .A2(new_n954), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT45), .Z(new_n961));
  NOR2_X1   g0761(.A1(new_n662), .A2(new_n954), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT44), .ZN(new_n963));
  AND4_X1   g0763(.A1(new_n657), .A2(new_n658), .A3(new_n961), .A4(new_n963), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n657), .A2(new_n658), .B1(new_n961), .B2(new_n963), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n649), .A2(G330), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n510), .A2(new_n661), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n655), .B2(new_n661), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n967), .B(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n709), .B1(new_n966), .B2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n665), .B(KEYINPUT41), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n959), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n932), .B1(new_n958), .B2(new_n973), .ZN(G387));
  INV_X1    g0774(.A(new_n970), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n975), .A2(new_n709), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n709), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n976), .A2(new_n665), .A3(new_n977), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n803), .A2(G311), .B1(G322), .B2(new_n753), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n979), .B1(new_n557), .B2(new_n733), .C1(new_n762), .C2(new_n745), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT48), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n981), .B1(new_n757), .B2(new_n725), .C1(new_n490), .C2(new_n730), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT49), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n368), .B1(new_n736), .B2(new_n215), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(new_n739), .B2(new_n755), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n726), .A2(new_n419), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n745), .A2(new_n213), .B1(new_n274), .B2(new_n736), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n791), .A2(G77), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n989), .B1(new_n741), .B2(new_n752), .C1(new_n740), .C2(new_n328), .ZN(new_n990));
  NOR4_X1   g0790(.A1(new_n987), .A2(new_n368), .A3(new_n988), .A4(new_n990), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n991), .B1(new_n233), .B2(new_n733), .C1(new_n329), .C2(new_n748), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n782), .B1(new_n986), .B2(new_n992), .ZN(new_n993));
  NOR3_X1   g0793(.A1(new_n655), .A2(G20), .A3(new_n718), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n930), .B1(new_n245), .B2(G45), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(new_n666), .B2(new_n772), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n378), .A2(new_n213), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT50), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n233), .A2(new_n210), .ZN(new_n999));
  NOR4_X1   g0799(.A1(new_n998), .A2(G45), .A3(new_n999), .A4(new_n666), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n996), .A2(new_n1000), .B1(G107), .B2(new_n205), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n1001), .A2(new_n775), .ZN(new_n1002));
  NOR4_X1   g0802(.A1(new_n993), .A2(new_n714), .A3(new_n994), .A4(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(new_n975), .B2(new_n959), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n978), .A2(new_n1004), .ZN(G393));
  NOR2_X1   g0805(.A1(new_n733), .A2(new_n329), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n726), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(G77), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G159), .A2(new_n746), .B1(new_n753), .B2(G150), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1009), .A2(KEYINPUT51), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n740), .A2(new_n912), .B1(new_n588), .B2(new_n736), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n368), .B1(new_n803), .B2(G50), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n791), .A2(G68), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1008), .A2(new_n1012), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n1006), .B(new_n1015), .C1(KEYINPUT51), .C2(new_n1009), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n759), .A2(new_n745), .B1(new_n752), .B2(new_n762), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT52), .Z(new_n1018));
  AOI22_X1  g0818(.A1(new_n803), .A2(G303), .B1(G107), .B2(new_n792), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n730), .A2(new_n757), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n268), .B(new_n1020), .C1(new_n739), .C2(G322), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1019), .B(new_n1021), .C1(new_n215), .C2(new_n725), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1018), .B(new_n1022), .C1(G294), .C2(new_n734), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n721), .B1(new_n1016), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n939), .A2(new_n719), .A3(new_n953), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n249), .A2(new_n770), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n775), .B(new_n1026), .C1(new_n274), .C2(new_n205), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1024), .A2(new_n778), .A3(new_n1025), .A4(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n959), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1028), .B1(new_n966), .B2(new_n1029), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n966), .A2(new_n977), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n711), .B1(new_n966), .B2(new_n977), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1030), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(G390));
  NAND3_X1  g0834(.A1(new_n708), .A2(G330), .A3(new_n881), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n871), .A2(new_n860), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n859), .B2(new_n863), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n688), .A2(new_n642), .A3(new_n820), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n807), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n860), .B1(new_n1040), .B2(new_n869), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n1041), .A2(new_n857), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1036), .B1(new_n1038), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1041), .A2(new_n857), .ZN(new_n1044));
  AND3_X1   g0844(.A1(new_n862), .A2(KEYINPUT39), .A3(new_n855), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n858), .B2(new_n857), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1044), .B(new_n1035), .C1(new_n1046), .C2(new_n1037), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1043), .A2(new_n1047), .A3(new_n959), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1046), .A2(new_n718), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n813), .A2(new_n329), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n1007), .A2(G77), .B1(G68), .B2(new_n792), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n734), .A2(G97), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n268), .B1(new_n803), .B2(G107), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n215), .A2(new_n745), .B1(new_n752), .B2(new_n757), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n731), .B(new_n1054), .C1(G294), .C2(new_n739), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .A4(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(G125), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n920), .A2(new_n784), .B1(new_n1057), .B2(new_n740), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n1007), .B2(G159), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n746), .A2(G132), .ZN(new_n1060));
  XOR2_X1   g0860(.A(KEYINPUT54), .B(G143), .Z(new_n1061));
  AOI22_X1  g0861(.A1(new_n753), .A2(G128), .B1(new_n734), .B2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n730), .A2(new_n328), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT53), .ZN(new_n1064));
  AND3_X1   g0864(.A1(new_n1062), .A2(new_n268), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1059), .A2(new_n1060), .A3(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n736), .A2(new_n213), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1056), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n721), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1049), .A2(new_n778), .A3(new_n1050), .A4(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n455), .A2(G330), .A3(new_n708), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n620), .A2(new_n875), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n817), .A2(new_n807), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n706), .A2(new_n707), .A3(G330), .A4(new_n811), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n870), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1073), .B1(new_n1036), .B2(new_n1076), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1035), .A2(new_n1075), .A3(new_n807), .A4(new_n1039), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1072), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1043), .A2(new_n1047), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n665), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1079), .B1(new_n1043), .B2(new_n1047), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1048), .B(new_n1070), .C1(new_n1081), .C2(new_n1082), .ZN(G378));
  AOI211_X1 g0883(.A(new_n268), .B(new_n257), .C1(new_n746), .C2(G107), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n419), .B2(new_n733), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n1085), .B(new_n909), .C1(G283), .C2(new_n739), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n208), .B2(new_n736), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n989), .B1(new_n748), .B2(new_n274), .C1(new_n752), .C2(new_n215), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT58), .Z(new_n1090));
  OAI221_X1 g0890(.A(new_n213), .B1(G33), .B2(G41), .C1(new_n268), .C2(new_n257), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1007), .A2(G150), .B1(G137), .B2(new_n734), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n746), .A2(G128), .B1(new_n749), .B2(G132), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1092), .B(new_n1093), .C1(new_n1057), .C2(new_n752), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(new_n791), .B2(new_n1061), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT59), .Z(new_n1096));
  AOI211_X1 g0896(.A(G33), .B(G41), .C1(new_n739), .C2(G124), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n741), .B2(new_n736), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1090), .B(new_n1091), .C1(new_n1096), .C2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n714), .B1(new_n1099), .B2(new_n721), .ZN(new_n1100));
  XOR2_X1   g0900(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1101));
  XNOR2_X1  g0901(.A(new_n348), .B(new_n1101), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n334), .A2(new_n830), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1102), .B(new_n1103), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n1100), .B1(G50), .B2(new_n814), .C1(new_n718), .C2(new_n1104), .ZN(new_n1105));
  XOR2_X1   g0905(.A(new_n1105), .B(KEYINPUT121), .Z(new_n1106));
  NAND2_X1  g0906(.A1(new_n864), .A2(new_n873), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n888), .A2(new_n889), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n857), .A2(new_n890), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1104), .ZN(new_n1110));
  AND4_X1   g0910(.A1(G330), .A2(new_n1108), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1110), .B1(new_n891), .B2(G330), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1107), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1108), .A2(G330), .A3(new_n1109), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n1104), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n891), .A2(G330), .A3(new_n1110), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n874), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1106), .B1(new_n1118), .B2(new_n1029), .ZN(new_n1119));
  AND3_X1   g0919(.A1(new_n1113), .A2(new_n1117), .A3(KEYINPUT57), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n1072), .B(KEYINPUT122), .Z(new_n1121));
  NAND2_X1  g0921(.A1(new_n1080), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n711), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT57), .ZN(new_n1124));
  AND2_X1   g0924(.A1(new_n1080), .A2(new_n1121), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1124), .B1(new_n1125), .B2(new_n1118), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1119), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(G375));
  AND2_X1   g0928(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1129), .A2(new_n1029), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n813), .A2(new_n233), .ZN(new_n1131));
  NOR3_X1   g0931(.A1(new_n869), .A2(G13), .A3(G33), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n726), .A2(new_n419), .B1(new_n920), .B2(new_n215), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n740), .A2(new_n557), .B1(new_n210), .B2(new_n736), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n757), .A2(new_n745), .B1(new_n752), .B2(new_n490), .ZN(new_n1135));
  NOR4_X1   g0935(.A1(new_n1133), .A2(new_n268), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n1136), .B1(new_n274), .B2(new_n730), .C1(new_n224), .C2(new_n733), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n745), .A2(new_n784), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n739), .A2(G128), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT123), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n368), .B1(new_n792), .B2(G58), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n1139), .B1(new_n1140), .B2(new_n1141), .C1(new_n328), .C2(new_n733), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1138), .B(new_n1142), .C1(new_n803), .C2(new_n1061), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1141), .A2(new_n1140), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n791), .A2(G159), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n1007), .A2(G50), .B1(G132), .B2(new_n753), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .A4(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n782), .B1(new_n1137), .B2(new_n1147), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n1132), .A2(new_n714), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1130), .B1(new_n1131), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1129), .A2(new_n1072), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1079), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1151), .A2(new_n972), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1150), .A2(new_n1153), .ZN(G381));
  OAI211_X1 g0954(.A(new_n932), .B(new_n1033), .C1(new_n958), .C2(new_n973), .ZN(new_n1155));
  OR2_X1    g0955(.A1(G393), .A2(G396), .ZN(new_n1156));
  NOR4_X1   g0956(.A1(new_n1155), .A2(G384), .A3(G381), .A4(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(G378), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1157), .A2(new_n1158), .A3(new_n1127), .ZN(G407));
  NAND2_X1  g0959(.A1(new_n640), .A2(G213), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n1160), .B(KEYINPUT124), .Z(new_n1161));
  NOR2_X1   g0961(.A1(new_n1157), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1127), .A2(new_n1158), .ZN(new_n1163));
  OAI21_X1  g0963(.A(G213), .B1(new_n1162), .B2(new_n1163), .ZN(G409));
  NAND2_X1  g0964(.A1(G393), .A2(G396), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1156), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(KEYINPUT126), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT126), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1156), .A2(new_n1168), .A3(new_n1165), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(G387), .A2(G390), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n1155), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1167), .A2(new_n1169), .B1(new_n1171), .B2(new_n1155), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT60), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n665), .B(new_n1152), .C1(new_n1151), .C2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(KEYINPUT60), .B1(new_n1129), .B2(new_n1072), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1150), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n825), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1150), .B(G384), .C1(new_n1177), .C2(new_n1178), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1161), .A2(G2897), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1182), .A2(G2897), .A3(new_n1161), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(new_n1111), .A2(new_n1112), .A3(new_n1107), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n1115), .A2(new_n1116), .B1(new_n864), .B2(new_n873), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  AND2_X1   g0989(.A1(new_n1122), .A2(new_n972), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1189), .B1(new_n1190), .B2(new_n959), .ZN(new_n1191));
  AOI21_X1  g0991(.A(G378), .B1(new_n1191), .B2(new_n1105), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1105), .B(KEYINPUT121), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n1189), .B2(new_n959), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1113), .A2(new_n1117), .A3(KEYINPUT57), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n665), .B1(new_n1125), .B2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT57), .B1(new_n1189), .B2(new_n1122), .ZN(new_n1197));
  OAI211_X1 g0997(.A(G378), .B(new_n1194), .C1(new_n1196), .C2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(KEYINPUT125), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT125), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1200), .A2(new_n1201), .A3(G378), .A4(new_n1194), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1192), .B1(new_n1199), .B2(new_n1202), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1185), .B(new_n1186), .C1(new_n1203), .C2(new_n1161), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n1203), .A2(new_n1161), .A3(new_n1182), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT62), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1204), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1192), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1201), .B1(new_n1127), .B2(G378), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1198), .A2(KEYINPUT125), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1208), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1161), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1211), .A2(new_n1206), .A3(new_n1212), .A4(new_n1183), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT61), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1175), .B1(new_n1207), .B2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1211), .A2(new_n1212), .A3(new_n1183), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT63), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1217), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1214), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n1205), .B2(KEYINPUT63), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1221), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1216), .A2(new_n1224), .ZN(G405));
  NAND2_X1  g1025(.A1(new_n1199), .A2(new_n1202), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(G375), .A2(new_n1158), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT127), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1228), .A2(new_n1229), .A3(new_n1182), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1183), .A2(KEYINPUT127), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1182), .A2(new_n1229), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1226), .A2(new_n1231), .A3(new_n1232), .A4(new_n1227), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1230), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1175), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1234), .B(new_n1235), .ZN(G402));
endmodule


