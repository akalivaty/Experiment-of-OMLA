//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 1 1 1 0 1 0 1 0 0 1 0 0 0 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985;
  XOR2_X1   g000(.A(G155gat), .B(G162gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G141gat), .B(G148gat), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(KEYINPUT2), .B2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT78), .B(G162gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G155gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT2), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n202), .A2(new_n203), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT79), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT79), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n208), .A2(new_n212), .A3(new_n209), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n205), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G211gat), .B(G218gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n215), .B(KEYINPUT74), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n217));
  OR2_X1    g016(.A1(G197gat), .A2(G204gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(G197gat), .A2(G204gat), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n216), .B(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT29), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n214), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT82), .ZN(new_n226));
  INV_X1    g025(.A(G228gat), .ZN(new_n227));
  INV_X1    g026(.A(G233gat), .ZN(new_n228));
  OAI22_X1  g027(.A1(new_n225), .A2(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G22gat), .ZN(new_n230));
  INV_X1    g029(.A(G22gat), .ZN(new_n231));
  OAI221_X1 g030(.A(new_n231), .B1(new_n227), .B2(new_n228), .C1(new_n225), .C2(new_n226), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT31), .B(G50gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n234), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n230), .A2(new_n232), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n214), .A2(new_n224), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n221), .B1(new_n239), .B2(new_n222), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n240), .A2(new_n225), .ZN(new_n241));
  XNOR2_X1  g040(.A(G78gat), .B(G106gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n238), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n235), .A2(new_n243), .A3(new_n237), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(KEYINPUT80), .B(KEYINPUT4), .Z(new_n248));
  INV_X1    g047(.A(G120gat), .ZN(new_n249));
  AND2_X1   g048(.A1(new_n249), .A2(G113gat), .ZN(new_n250));
  OR2_X1    g049(.A1(new_n250), .A2(KEYINPUT70), .ZN(new_n251));
  OAI21_X1  g050(.A(KEYINPUT71), .B1(new_n249), .B2(G113gat), .ZN(new_n252));
  OR3_X1    g051(.A1(new_n249), .A2(KEYINPUT71), .A3(G113gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n250), .A2(KEYINPUT70), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n251), .A2(new_n252), .A3(new_n253), .A4(new_n254), .ZN(new_n255));
  XOR2_X1   g054(.A(G127gat), .B(G134gat), .Z(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(KEYINPUT1), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n249), .A2(G113gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n250), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n256), .B1(new_n260), .B2(KEYINPUT1), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(new_n214), .ZN(new_n264));
  MUX2_X1   g063(.A(new_n248), .B(KEYINPUT4), .S(new_n264), .Z(new_n265));
  INV_X1    g064(.A(KEYINPUT5), .ZN(new_n266));
  NAND2_X1  g065(.A1(G225gat), .A2(G233gat), .ZN(new_n267));
  INV_X1    g066(.A(new_n213), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n212), .B1(new_n208), .B2(new_n209), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n204), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n271), .A2(new_n239), .A3(new_n262), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n265), .A2(new_n266), .A3(new_n267), .A4(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n264), .A2(new_n248), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n263), .A2(new_n214), .A3(KEYINPUT4), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n272), .A2(new_n274), .A3(new_n267), .A4(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n270), .A2(new_n262), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n264), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n267), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n266), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AND3_X1   g079(.A1(new_n276), .A2(KEYINPUT81), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT81), .B1(new_n276), .B2(new_n280), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n273), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G1gat), .B(G29gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(KEYINPUT0), .ZN(new_n285));
  XNOR2_X1  g084(.A(G57gat), .B(G85gat), .ZN(new_n286));
  XOR2_X1   g085(.A(new_n285), .B(new_n286), .Z(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n283), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n273), .B(new_n287), .C1(new_n281), .C2(new_n282), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n283), .A2(KEYINPUT6), .A3(new_n288), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G8gat), .B(G36gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(G64gat), .B(G92gat), .ZN(new_n297));
  XOR2_X1   g096(.A(new_n296), .B(new_n297), .Z(new_n298));
  NAND2_X1  g097(.A1(G226gat), .A2(G233gat), .ZN(new_n299));
  XOR2_X1   g098(.A(new_n299), .B(KEYINPUT75), .Z(new_n300));
  INV_X1    g099(.A(KEYINPUT69), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT27), .B(G183gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n302), .B(KEYINPUT68), .ZN(new_n303));
  INV_X1    g102(.A(G190gat), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n304), .A2(KEYINPUT28), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n302), .A2(new_n304), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n307));
  AOI22_X1  g106(.A1(new_n303), .A2(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(G183gat), .A2(G190gat), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NOR2_X1   g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n310), .B1(KEYINPUT26), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT26), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n312), .B1(new_n311), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n301), .B1(new_n308), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NOR3_X1   g117(.A1(new_n308), .A2(new_n301), .A3(new_n316), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT25), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT24), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n310), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G183gat), .B(G190gat), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n322), .B1(new_n323), .B2(new_n321), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n311), .A2(KEYINPUT23), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT23), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n326), .B1(G169gat), .B2(G176gat), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n325), .A2(new_n313), .A3(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n320), .B1(new_n324), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n324), .A2(KEYINPUT64), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT64), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n322), .B(new_n332), .C1(new_n323), .C2(new_n321), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n328), .A2(new_n320), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n331), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT65), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT65), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n331), .A2(new_n337), .A3(new_n333), .A4(new_n334), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n330), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT66), .ZN(new_n340));
  OAI22_X1  g139(.A1(new_n318), .A2(new_n319), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AOI211_X1 g140(.A(KEYINPUT66), .B(new_n330), .C1(new_n336), .C2(new_n338), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n300), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n303), .A2(new_n305), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n306), .A2(new_n307), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n316), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n339), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n299), .B1(new_n347), .B2(KEYINPUT29), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n343), .A2(new_n221), .A3(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n347), .A2(new_n299), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n222), .B1(new_n341), .B2(new_n342), .ZN(new_n351));
  INV_X1    g150(.A(new_n300), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n298), .B(new_n349), .C1(new_n353), .C2(new_n221), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT30), .ZN(new_n355));
  INV_X1    g154(.A(new_n221), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n336), .A2(new_n338), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(new_n329), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n346), .A2(KEYINPUT69), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n358), .A2(KEYINPUT66), .B1(new_n317), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n342), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n300), .B1(new_n362), .B2(new_n222), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n356), .B1(new_n363), .B2(new_n350), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT30), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n364), .A2(new_n365), .A3(new_n298), .A4(new_n349), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n355), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n349), .B1(new_n353), .B2(new_n221), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT77), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n298), .B(KEYINPUT76), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n369), .B1(new_n368), .B2(new_n370), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n367), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n247), .B1(new_n295), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT73), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT36), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(KEYINPUT73), .A2(KEYINPUT36), .ZN(new_n379));
  XNOR2_X1  g178(.A(G15gat), .B(G43gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(G71gat), .B(G99gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n380), .B(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(G227gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n383), .A2(new_n228), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n263), .B1(new_n360), .B2(new_n361), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n341), .A2(new_n262), .A3(new_n342), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n382), .B1(new_n387), .B2(KEYINPUT32), .ZN(new_n388));
  INV_X1    g187(.A(new_n384), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n262), .B1(new_n341), .B2(new_n342), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n360), .A2(new_n263), .A3(new_n361), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT72), .B1(new_n392), .B2(KEYINPUT33), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT72), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT33), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n387), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n388), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n390), .A2(new_n391), .A3(new_n389), .ZN(new_n398));
  XOR2_X1   g197(.A(new_n398), .B(KEYINPUT34), .Z(new_n399));
  OAI211_X1 g198(.A(new_n387), .B(KEYINPUT32), .C1(new_n395), .C2(new_n382), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n397), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n399), .B1(new_n397), .B2(new_n400), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n378), .B(new_n379), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n397), .A2(new_n400), .ZN(new_n404));
  INV_X1    g203(.A(new_n399), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n397), .A2(new_n399), .A3(new_n400), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n406), .A2(new_n376), .A3(new_n377), .A4(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n375), .A2(new_n403), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT83), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT83), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n375), .A2(new_n403), .A3(new_n408), .A4(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n298), .B1(new_n368), .B2(KEYINPUT37), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT86), .ZN(new_n414));
  OAI22_X1  g213(.A1(new_n413), .A2(new_n414), .B1(KEYINPUT37), .B2(new_n368), .ZN(new_n415));
  AND2_X1   g214(.A1(new_n413), .A2(new_n414), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT38), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n343), .A2(new_n356), .A3(new_n348), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n418), .B(KEYINPUT37), .C1(new_n353), .C2(new_n356), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT38), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n370), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n419), .B(new_n421), .C1(new_n368), .C2(KEYINPUT37), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT85), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n417), .A2(new_n295), .A3(new_n424), .A4(new_n354), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n267), .B1(new_n265), .B2(new_n272), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n278), .A2(new_n279), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n428), .B(KEYINPUT84), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n427), .A2(new_n429), .A3(KEYINPUT39), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT39), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n288), .B1(new_n426), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT40), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n430), .A2(KEYINPUT40), .A3(new_n432), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n435), .A2(new_n289), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n247), .B1(new_n437), .B2(new_n374), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n425), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n410), .A2(new_n412), .A3(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(KEYINPUT87), .B(KEYINPUT35), .ZN(new_n441));
  NOR3_X1   g240(.A1(new_n401), .A2(new_n402), .A3(new_n247), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n295), .A2(new_n374), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n245), .A2(new_n246), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n406), .A2(new_n407), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n373), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n371), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n294), .A2(new_n448), .A3(new_n367), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT35), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n450), .A2(KEYINPUT87), .ZN(new_n451));
  NOR3_X1   g250(.A1(new_n446), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n444), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n440), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT89), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI211_X1 g257(.A(KEYINPUT89), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g259(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n461));
  INV_X1    g260(.A(G36gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT90), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n458), .A2(new_n459), .B1(new_n462), .B2(new_n461), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT90), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(KEYINPUT91), .B(G36gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(G29gat), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n465), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(G43gat), .B(G50gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT15), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n463), .A2(new_n456), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n475), .B(KEYINPUT92), .ZN(new_n476));
  OR2_X1    g275(.A1(new_n472), .A2(KEYINPUT15), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n477), .A2(new_n473), .A3(new_n470), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n471), .A2(new_n474), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT17), .ZN(new_n480));
  INV_X1    g279(.A(new_n468), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n470), .B1(new_n466), .B2(new_n467), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n474), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n478), .A2(new_n476), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT17), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(G15gat), .B(G22gat), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n488), .A2(G1gat), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT93), .ZN(new_n490));
  OAI21_X1  g289(.A(G8gat), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT16), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n488), .B1(new_n492), .B2(G1gat), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n493), .B1(G1gat), .B2(new_n488), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n491), .B(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n480), .A2(new_n487), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(G229gat), .A2(G233gat), .ZN(new_n497));
  INV_X1    g296(.A(new_n495), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n485), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n496), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT18), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n496), .A2(KEYINPUT18), .A3(new_n497), .A4(new_n499), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n479), .A2(new_n495), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(KEYINPUT94), .B(KEYINPUT13), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(new_n497), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G113gat), .B(G141gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(G169gat), .B(G197gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n512), .B(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT12), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n502), .A2(new_n503), .A3(new_n509), .A4(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT95), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n500), .A2(new_n501), .B1(new_n505), .B2(new_n508), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT95), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n518), .A2(new_n519), .A3(new_n503), .A4(new_n515), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n518), .A2(new_n503), .ZN(new_n522));
  INV_X1    g321(.A(new_n515), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(G230gat), .A2(G233gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT102), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT7), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n529), .A2(G85gat), .A3(G92gat), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G99gat), .A2(G106gat), .ZN(new_n532));
  INV_X1    g331(.A(G85gat), .ZN(new_n533));
  INV_X1    g332(.A(G92gat), .ZN(new_n534));
  AOI22_X1  g333(.A1(KEYINPUT8), .A2(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n533), .A2(new_n534), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n531), .B(new_n535), .C1(new_n536), .C2(new_n529), .ZN(new_n537));
  XNOR2_X1  g336(.A(G99gat), .B(G106gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G71gat), .A2(G78gat), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT9), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(KEYINPUT97), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  AND2_X1   g343(.A1(G71gat), .A2(G78gat), .ZN(new_n545));
  NOR2_X1   g344(.A1(G71gat), .A2(G78gat), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT97), .B1(new_n541), .B2(new_n542), .ZN(new_n548));
  NOR3_X1   g347(.A1(new_n544), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(G57gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT98), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT98), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(G57gat), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n551), .A2(new_n553), .A3(G64gat), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT99), .ZN(new_n555));
  INV_X1    g354(.A(G64gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(G57gat), .ZN(new_n557));
  AND3_X1   g356(.A1(new_n554), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n555), .B1(new_n554), .B2(new_n557), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n549), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT97), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n561), .B1(new_n545), .B2(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n550), .A2(G64gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n557), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n562), .A2(new_n543), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n546), .A2(KEYINPUT96), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n546), .A2(KEYINPUT96), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n565), .A2(new_n541), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  AND3_X1   g367(.A1(new_n560), .A2(KEYINPUT100), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(KEYINPUT100), .B1(new_n560), .B2(new_n568), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n540), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n560), .A2(new_n568), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n539), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT10), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n539), .A2(KEYINPUT10), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT100), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n562), .B(new_n543), .C1(new_n545), .C2(new_n546), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n554), .A2(new_n557), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT99), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n554), .A2(new_n555), .A3(new_n557), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n577), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n567), .A2(new_n541), .A3(new_n566), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n544), .A2(new_n548), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n582), .B1(new_n583), .B2(new_n564), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n576), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n560), .A2(KEYINPUT100), .A3(new_n568), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n575), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n526), .B1(new_n574), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n526), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n571), .A2(new_n589), .A3(new_n573), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G120gat), .B(G148gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(G176gat), .B(G204gat), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n592), .B(new_n593), .Z(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n588), .A2(new_n590), .A3(new_n594), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n585), .A2(new_n586), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT21), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(new_n495), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT101), .B(KEYINPUT19), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G231gat), .A2(G233gat), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n605), .B1(new_n599), .B2(KEYINPUT21), .ZN(new_n606));
  XNOR2_X1  g405(.A(G127gat), .B(G155gat), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n607), .B(KEYINPUT20), .Z(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT21), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n585), .A2(new_n610), .A3(new_n586), .A4(new_n604), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n606), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(G183gat), .B(G211gat), .Z(new_n614));
  AOI21_X1  g413(.A(new_n609), .B1(new_n606), .B2(new_n611), .ZN(new_n615));
  NOR3_X1   g414(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n614), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n606), .A2(new_n611), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(new_n608), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n617), .B1(new_n619), .B2(new_n612), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n603), .B1(new_n616), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n480), .A2(new_n487), .A3(new_n540), .ZN(new_n622));
  AND2_X1   g421(.A1(G232gat), .A2(G233gat), .ZN(new_n623));
  AOI22_X1  g422(.A1(new_n485), .A2(new_n539), .B1(KEYINPUT41), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(G190gat), .B(G218gat), .Z(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n626), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n622), .A2(new_n628), .A3(new_n624), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n623), .A2(KEYINPUT41), .ZN(new_n631));
  XNOR2_X1  g430(.A(G134gat), .B(G162gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n627), .A2(new_n633), .A3(new_n629), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n603), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n614), .B1(new_n613), .B2(new_n615), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n619), .A2(new_n617), .A3(new_n612), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n598), .A2(new_n621), .A3(new_n637), .A4(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT103), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n621), .A2(new_n641), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT103), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n644), .A2(new_n645), .A3(new_n637), .A4(new_n598), .ZN(new_n646));
  AND4_X1   g445(.A1(new_n455), .A2(new_n525), .A3(new_n643), .A4(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n295), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g448(.A(KEYINPUT16), .B(G8gat), .Z(new_n650));
  AND3_X1   g449(.A1(new_n647), .A2(new_n374), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(G8gat), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n652), .B1(new_n647), .B2(new_n374), .ZN(new_n653));
  OAI21_X1  g452(.A(KEYINPUT42), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n654), .B1(KEYINPUT42), .B2(new_n651), .ZN(G1325gat));
  AND2_X1   g454(.A1(new_n403), .A2(new_n408), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  AND3_X1   g456(.A1(new_n647), .A2(G15gat), .A3(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n401), .A2(new_n402), .ZN(new_n659));
  AOI21_X1  g458(.A(G15gat), .B1(new_n647), .B2(new_n659), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n660), .A2(KEYINPUT104), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(KEYINPUT104), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n658), .B1(new_n661), .B2(new_n662), .ZN(G1326gat));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n247), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT43), .B(G22gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(G1327gat));
  AOI21_X1  g465(.A(new_n637), .B1(new_n440), .B2(new_n454), .ZN(new_n667));
  INV_X1    g466(.A(G29gat), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n521), .A2(new_n524), .ZN(new_n669));
  INV_X1    g468(.A(new_n598), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n669), .A2(new_n644), .A3(new_n670), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n667), .A2(new_n668), .A3(new_n295), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT45), .ZN(new_n673));
  INV_X1    g472(.A(new_n671), .ZN(new_n674));
  AOI22_X1  g473(.A1(new_n409), .A2(KEYINPUT83), .B1(new_n425), .B2(new_n438), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n453), .B1(new_n675), .B2(new_n412), .ZN(new_n676));
  OAI21_X1  g475(.A(KEYINPUT44), .B1(new_n676), .B2(new_n637), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n425), .A2(new_n438), .ZN(new_n678));
  OAI22_X1  g477(.A1(new_n678), .A2(new_n409), .B1(new_n444), .B2(new_n452), .ZN(new_n679));
  INV_X1    g478(.A(new_n637), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n674), .B1(new_n677), .B2(new_n682), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n683), .A2(new_n295), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n673), .B1(new_n684), .B2(new_n668), .ZN(G1328gat));
  INV_X1    g484(.A(new_n469), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n686), .B1(new_n683), .B2(new_n374), .ZN(new_n687));
  INV_X1    g486(.A(new_n374), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n688), .A2(new_n469), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n455), .A2(new_n680), .A3(new_n671), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(KEYINPUT106), .B(KEYINPUT46), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(KEYINPUT107), .B1(new_n687), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n682), .B1(new_n667), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n695), .A2(new_n374), .A3(new_n671), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n469), .ZN(new_n697));
  INV_X1    g496(.A(new_n691), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n690), .B(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT107), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n697), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n693), .A2(new_n701), .ZN(G1329gat));
  NAND4_X1  g501(.A1(new_n695), .A2(G43gat), .A3(new_n657), .A4(new_n671), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n667), .A2(new_n671), .ZN(new_n704));
  INV_X1    g503(.A(new_n659), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n703), .B1(G43gat), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(KEYINPUT47), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT47), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n703), .B(new_n709), .C1(G43gat), .C2(new_n706), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(G1330gat));
  NAND4_X1  g510(.A1(new_n695), .A2(G50gat), .A3(new_n247), .A4(new_n671), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n704), .A2(new_n445), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n712), .B1(G50gat), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(KEYINPUT48), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT48), .ZN(new_n716));
  OAI211_X1 g515(.A(new_n712), .B(new_n716), .C1(G50gat), .C2(new_n713), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(G1331gat));
  INV_X1    g517(.A(new_n644), .ZN(new_n719));
  NOR4_X1   g518(.A1(new_n719), .A2(new_n525), .A3(new_n680), .A4(new_n598), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n679), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n295), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n551), .A2(new_n553), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1332gat));
  AOI21_X1  g523(.A(new_n688), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(KEYINPUT108), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT108), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n721), .A2(new_n728), .A3(new_n725), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  OR2_X1    g529(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(G1333gat));
  INV_X1    g531(.A(G71gat), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n721), .A2(new_n733), .A3(new_n659), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n721), .A2(new_n657), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n734), .B1(new_n735), .B2(new_n733), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT50), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1334gat));
  NAND2_X1  g537(.A1(new_n721), .A2(new_n247), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT109), .B(G78gat), .Z(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1335gat));
  NOR2_X1   g540(.A1(new_n525), .A2(new_n644), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n670), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n743), .B1(new_n677), .B2(new_n682), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n744), .A2(new_n295), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n679), .A2(new_n680), .A3(new_n742), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT51), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT51), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n679), .A2(new_n748), .A3(new_n680), .A4(new_n742), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n747), .A2(new_n670), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n295), .A2(new_n533), .ZN(new_n751));
  OAI22_X1  g550(.A1(new_n745), .A2(new_n533), .B1(new_n750), .B2(new_n751), .ZN(G1336gat));
  AOI21_X1  g551(.A(new_n534), .B1(new_n744), .B2(new_n374), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n688), .A2(G92gat), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n747), .A2(new_n670), .A3(new_n749), .A4(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(KEYINPUT52), .B1(new_n753), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT52), .ZN(new_n758));
  AOI211_X1 g557(.A(new_n688), .B(new_n743), .C1(new_n677), .C2(new_n682), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n758), .B(new_n755), .C1(new_n759), .C2(new_n534), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n757), .A2(new_n760), .ZN(G1337gat));
  OR3_X1    g560(.A1(new_n750), .A2(G99gat), .A3(new_n705), .ZN(new_n762));
  INV_X1    g561(.A(new_n743), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n695), .A2(new_n657), .A3(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT110), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(G99gat), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n764), .A2(new_n765), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n762), .B1(new_n767), .B2(new_n768), .ZN(G1338gat));
  INV_X1    g568(.A(G106gat), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n744), .B2(new_n247), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n445), .A2(G106gat), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n747), .A2(new_n670), .A3(new_n749), .A4(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(KEYINPUT53), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT53), .ZN(new_n776));
  AOI211_X1 g575(.A(new_n445), .B(new_n743), .C1(new_n677), .C2(new_n682), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n776), .B(new_n773), .C1(new_n777), .C2(new_n770), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n775), .A2(new_n778), .ZN(G1339gat));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT10), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n539), .B1(new_n585), .B2(new_n586), .ZN(new_n782));
  INV_X1    g581(.A(new_n573), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n599), .A2(KEYINPUT10), .A3(new_n539), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n780), .B1(new_n786), .B2(new_n526), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n571), .A2(new_n573), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n587), .B1(new_n788), .B2(new_n781), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT111), .B1(new_n789), .B2(new_n589), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n791));
  NOR4_X1   g590(.A1(new_n574), .A2(new_n791), .A3(new_n587), .A4(new_n526), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n787), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  AOI211_X1 g592(.A(KEYINPUT54), .B(new_n589), .C1(new_n784), .C2(new_n785), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT112), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n794), .A2(new_n795), .A3(new_n594), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n786), .A2(new_n780), .A3(new_n526), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT112), .B1(new_n797), .B2(new_n595), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n793), .B(KEYINPUT55), .C1(new_n796), .C2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n597), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n799), .A2(KEYINPUT113), .A3(new_n597), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n796), .A2(new_n798), .ZN(new_n805));
  INV_X1    g604(.A(new_n793), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n802), .A2(new_n525), .A3(new_n803), .A4(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(KEYINPUT114), .B1(new_n505), .B2(new_n508), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n499), .A2(new_n504), .A3(new_n810), .A4(new_n507), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n497), .B1(new_n496), .B2(new_n499), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n514), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT115), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n816), .B(new_n514), .C1(new_n812), .C2(new_n813), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n670), .A2(new_n818), .A3(new_n521), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n680), .B1(new_n808), .B2(new_n819), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n818), .A2(new_n521), .A3(new_n680), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n802), .A2(new_n821), .A3(new_n803), .A4(new_n807), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n719), .B1(new_n820), .B2(new_n823), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n642), .A2(new_n525), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n446), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n374), .A2(new_n294), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n525), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n670), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n249), .A2(KEYINPUT116), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n249), .A2(KEYINPUT116), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n834), .B1(new_n831), .B2(new_n832), .ZN(G1341gat));
  NAND2_X1  g634(.A1(new_n828), .A2(new_n644), .ZN(new_n836));
  INV_X1    g635(.A(G127gat), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n836), .A2(KEYINPUT117), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n828), .A2(G127gat), .A3(new_n644), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n839), .A2(KEYINPUT117), .ZN(new_n840));
  AOI211_X1 g639(.A(new_n838), .B(new_n840), .C1(new_n837), .C2(new_n836), .ZN(G1342gat));
  INV_X1    g640(.A(G134gat), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n374), .A2(new_n294), .A3(new_n637), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n826), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(KEYINPUT56), .ZN(new_n845));
  XOR2_X1   g644(.A(new_n845), .B(KEYINPUT118), .Z(new_n846));
  NAND2_X1  g645(.A1(new_n826), .A2(new_n843), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(G134gat), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n846), .B(new_n848), .C1(KEYINPUT56), .C2(new_n844), .ZN(G1343gat));
  INV_X1    g648(.A(KEYINPUT120), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n656), .A2(new_n827), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n824), .A2(new_n825), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT57), .B1(new_n852), .B2(new_n247), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n445), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n597), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n795), .B1(new_n794), .B2(new_n594), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n797), .A2(KEYINPUT112), .A3(new_n595), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n789), .A2(KEYINPUT111), .A3(new_n589), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n784), .A2(new_n589), .A3(new_n785), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n791), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  AOI22_X1  g662(.A1(new_n858), .A2(new_n859), .B1(new_n863), .B2(new_n787), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n857), .B1(new_n864), .B2(KEYINPUT55), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n804), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n793), .B(new_n866), .C1(new_n796), .C2(new_n798), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n525), .B(new_n865), .C1(new_n867), .C2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n680), .B1(new_n870), .B2(new_n819), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n719), .B1(new_n871), .B2(new_n823), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n856), .B1(new_n872), .B2(new_n825), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n525), .B(new_n851), .C1(new_n853), .C2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n850), .B1(new_n874), .B2(G141gat), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n445), .B1(new_n824), .B2(new_n825), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n669), .A2(G141gat), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n876), .A2(new_n851), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n878), .B1(new_n874), .B2(G141gat), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n875), .A2(new_n879), .A3(KEYINPUT58), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT58), .ZN(new_n881));
  AOI221_X4 g680(.A(new_n878), .B1(new_n850), .B2(new_n881), .C1(new_n874), .C2(G141gat), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n880), .A2(new_n882), .ZN(G1344gat));
  INV_X1    g682(.A(G148gat), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(KEYINPUT59), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n851), .B1(new_n853), .B2(new_n873), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n885), .B1(new_n886), .B2(new_n598), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n851), .A2(new_n670), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n646), .A2(new_n643), .A3(new_n669), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(KEYINPUT121), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n646), .A2(new_n643), .A3(new_n891), .A4(new_n669), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n819), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n669), .A2(new_n800), .ZN(new_n895));
  OAI21_X1  g694(.A(KEYINPUT119), .B1(new_n805), .B2(new_n806), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n896), .A2(new_n804), .A3(new_n868), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n894), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n822), .B1(new_n898), .B2(new_n680), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n893), .B1(new_n899), .B2(new_n719), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n854), .B1(new_n900), .B2(new_n445), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n852), .A2(new_n855), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n888), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(KEYINPUT59), .B1(new_n903), .B2(new_n884), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n887), .A2(new_n904), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n876), .A2(new_n851), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(new_n884), .A3(new_n670), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n905), .A2(new_n907), .ZN(G1345gat));
  OAI21_X1  g707(.A(G155gat), .B1(new_n886), .B2(new_n719), .ZN(new_n909));
  INV_X1    g708(.A(G155gat), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n906), .A2(new_n910), .A3(new_n644), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n911), .ZN(G1346gat));
  OAI21_X1  g711(.A(new_n206), .B1(new_n886), .B2(new_n637), .ZN(new_n913));
  INV_X1    g712(.A(new_n843), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n657), .A2(new_n206), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n876), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT122), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n913), .A2(new_n917), .ZN(G1347gat));
  NOR2_X1   g717(.A1(new_n688), .A2(new_n295), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(KEYINPUT124), .A3(new_n659), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT124), .ZN(new_n921));
  INV_X1    g720(.A(new_n919), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n921), .B1(new_n922), .B2(new_n705), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n852), .A2(new_n445), .A3(new_n920), .A4(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(G169gat), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n924), .A2(new_n925), .A3(new_n669), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n852), .A2(KEYINPUT123), .A3(new_n294), .ZN(new_n927));
  AOI21_X1  g726(.A(KEYINPUT123), .B1(new_n852), .B2(new_n294), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n446), .A2(new_n688), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n929), .A2(new_n525), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n926), .B1(new_n931), .B2(new_n925), .ZN(G1348gat));
  INV_X1    g731(.A(G176gat), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n924), .A2(new_n933), .A3(new_n598), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT125), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n670), .B(new_n930), .C1(new_n927), .C2(new_n928), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n935), .B1(new_n937), .B2(G176gat), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n936), .A2(KEYINPUT125), .A3(new_n933), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n934), .B1(new_n938), .B2(new_n939), .ZN(G1349gat));
  AND2_X1   g739(.A1(new_n644), .A2(new_n303), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n930), .B(new_n941), .C1(new_n927), .C2(new_n928), .ZN(new_n942));
  OAI21_X1  g741(.A(G183gat), .B1(new_n924), .B2(new_n719), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT60), .ZN(G1350gat));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n680), .A2(new_n304), .ZN(new_n947));
  OAI21_X1  g746(.A(G190gat), .B1(new_n924), .B2(new_n637), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n948), .A2(KEYINPUT61), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n948), .A2(KEYINPUT61), .ZN(new_n950));
  OAI22_X1  g749(.A1(new_n946), .A2(new_n947), .B1(new_n949), .B2(new_n950), .ZN(G1351gat));
  NOR3_X1   g750(.A1(new_n657), .A2(new_n688), .A3(new_n445), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n929), .A2(new_n525), .A3(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(G197gat), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n657), .A2(new_n922), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n956), .B1(new_n901), .B2(new_n902), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n669), .A2(new_n954), .ZN(new_n958));
  AOI22_X1  g757(.A1(new_n953), .A2(new_n954), .B1(new_n957), .B2(new_n958), .ZN(G1352gat));
  INV_X1    g758(.A(new_n957), .ZN(new_n960));
  OAI21_X1  g759(.A(G204gat), .B1(new_n960), .B2(new_n598), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n598), .A2(G204gat), .ZN(new_n962));
  OAI211_X1 g761(.A(new_n952), .B(new_n962), .C1(new_n927), .C2(new_n928), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n963), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n964));
  AOI21_X1  g763(.A(KEYINPUT126), .B1(new_n963), .B2(KEYINPUT62), .ZN(new_n965));
  OAI221_X1 g764(.A(new_n961), .B1(KEYINPUT62), .B2(new_n963), .C1(new_n964), .C2(new_n965), .ZN(G1353gat));
  INV_X1    g765(.A(KEYINPUT63), .ZN(new_n967));
  INV_X1    g766(.A(new_n893), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n872), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g768(.A(KEYINPUT57), .B1(new_n969), .B2(new_n247), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n856), .B1(new_n824), .B2(new_n825), .ZN(new_n971));
  OAI211_X1 g770(.A(new_n644), .B(new_n955), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  OAI21_X1  g771(.A(G211gat), .B1(new_n972), .B2(KEYINPUT127), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT127), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n974), .B1(new_n957), .B2(new_n644), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n967), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n972), .A2(KEYINPUT127), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n957), .A2(new_n974), .A3(new_n644), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n977), .A2(new_n978), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n929), .A2(new_n952), .ZN(new_n981));
  OR3_X1    g780(.A1(new_n981), .A2(G211gat), .A3(new_n719), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n980), .A2(new_n982), .ZN(G1354gat));
  OAI21_X1  g782(.A(G218gat), .B1(new_n960), .B2(new_n637), .ZN(new_n984));
  OR2_X1    g783(.A1(new_n637), .A2(G218gat), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n984), .B1(new_n981), .B2(new_n985), .ZN(G1355gat));
endmodule


