

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U558 ( .A(KEYINPUT23), .B(KEYINPUT65), .ZN(n522) );
  INV_X1 U559 ( .A(KEYINPUT26), .ZN(n684) );
  XNOR2_X1 U560 ( .A(KEYINPUT96), .B(KEYINPUT27), .ZN(n678) );
  XNOR2_X1 U561 ( .A(n679), .B(n678), .ZN(n681) );
  XNOR2_X1 U562 ( .A(n712), .B(KEYINPUT97), .ZN(n713) );
  XNOR2_X1 U563 ( .A(n714), .B(n713), .ZN(n715) );
  NOR2_X1 U564 ( .A1(n718), .A2(n717), .ZN(n720) );
  NOR2_X1 U565 ( .A1(G1966), .A2(n766), .ZN(n734) );
  NAND2_X1 U566 ( .A1(n677), .A2(n772), .ZN(n723) );
  AND2_X1 U567 ( .A1(n527), .A2(G2104), .ZN(n873) );
  NOR2_X1 U568 ( .A1(G2104), .A2(n527), .ZN(n876) );
  NOR2_X1 U569 ( .A1(G651), .A2(n631), .ZN(n638) );
  XNOR2_X1 U570 ( .A(n523), .B(n522), .ZN(n526) );
  NOR2_X1 U571 ( .A1(n531), .A2(n530), .ZN(G160) );
  INV_X1 U572 ( .A(G2105), .ZN(n527) );
  NAND2_X1 U573 ( .A1(G101), .A2(n873), .ZN(n523) );
  NOR2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  XOR2_X2 U575 ( .A(KEYINPUT17), .B(n524), .Z(n872) );
  NAND2_X1 U576 ( .A1(G137), .A2(n872), .ZN(n525) );
  NAND2_X1 U577 ( .A1(n526), .A2(n525), .ZN(n531) );
  NAND2_X1 U578 ( .A1(G125), .A2(n876), .ZN(n529) );
  AND2_X1 U579 ( .A1(G2104), .A2(G2105), .ZN(n877) );
  NAND2_X1 U580 ( .A1(G113), .A2(n877), .ZN(n528) );
  NAND2_X1 U581 ( .A1(n529), .A2(n528), .ZN(n530) );
  NAND2_X1 U582 ( .A1(G114), .A2(n877), .ZN(n533) );
  NAND2_X1 U583 ( .A1(G102), .A2(n873), .ZN(n532) );
  AND2_X1 U584 ( .A1(n533), .A2(n532), .ZN(n535) );
  NAND2_X1 U585 ( .A1(G126), .A2(n876), .ZN(n534) );
  AND2_X1 U586 ( .A1(n535), .A2(n534), .ZN(n537) );
  NAND2_X1 U587 ( .A1(n872), .A2(G138), .ZN(n536) );
  AND2_X1 U588 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U589 ( .A(n538), .B(KEYINPUT85), .Z(G164) );
  NOR2_X1 U590 ( .A1(G651), .A2(G543), .ZN(n637) );
  NAND2_X1 U591 ( .A1(n637), .A2(G85), .ZN(n542) );
  XOR2_X1 U592 ( .A(G651), .B(KEYINPUT66), .Z(n543) );
  NOR2_X1 U593 ( .A1(G543), .A2(n543), .ZN(n539) );
  XNOR2_X1 U594 ( .A(n539), .B(KEYINPUT1), .ZN(n540) );
  XNOR2_X1 U595 ( .A(KEYINPUT67), .B(n540), .ZN(n646) );
  NAND2_X1 U596 ( .A1(G60), .A2(n646), .ZN(n541) );
  NAND2_X1 U597 ( .A1(n542), .A2(n541), .ZN(n547) );
  XOR2_X1 U598 ( .A(KEYINPUT0), .B(G543), .Z(n631) );
  NAND2_X1 U599 ( .A1(n638), .A2(G47), .ZN(n545) );
  NOR2_X1 U600 ( .A1(n631), .A2(n543), .ZN(n641) );
  NAND2_X1 U601 ( .A1(G72), .A2(n641), .ZN(n544) );
  NAND2_X1 U602 ( .A1(n545), .A2(n544), .ZN(n546) );
  OR2_X1 U603 ( .A1(n547), .A2(n546), .ZN(G290) );
  NAND2_X1 U604 ( .A1(n638), .A2(G52), .ZN(n549) );
  NAND2_X1 U605 ( .A1(G64), .A2(n646), .ZN(n548) );
  NAND2_X1 U606 ( .A1(n549), .A2(n548), .ZN(n555) );
  NAND2_X1 U607 ( .A1(G90), .A2(n637), .ZN(n551) );
  NAND2_X1 U608 ( .A1(G77), .A2(n641), .ZN(n550) );
  NAND2_X1 U609 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U610 ( .A(KEYINPUT9), .B(n552), .Z(n553) );
  XNOR2_X1 U611 ( .A(KEYINPUT68), .B(n553), .ZN(n554) );
  NOR2_X1 U612 ( .A1(n555), .A2(n554), .ZN(G171) );
  AND2_X1 U613 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U614 ( .A1(n876), .A2(G123), .ZN(n556) );
  XNOR2_X1 U615 ( .A(n556), .B(KEYINPUT18), .ZN(n558) );
  NAND2_X1 U616 ( .A1(G111), .A2(n877), .ZN(n557) );
  NAND2_X1 U617 ( .A1(n558), .A2(n557), .ZN(n562) );
  NAND2_X1 U618 ( .A1(G135), .A2(n872), .ZN(n560) );
  NAND2_X1 U619 ( .A1(G99), .A2(n873), .ZN(n559) );
  NAND2_X1 U620 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U621 ( .A1(n562), .A2(n561), .ZN(n925) );
  XNOR2_X1 U622 ( .A(n925), .B(G2096), .ZN(n563) );
  XNOR2_X1 U623 ( .A(n563), .B(KEYINPUT75), .ZN(n564) );
  OR2_X1 U624 ( .A1(G2100), .A2(n564), .ZN(G156) );
  INV_X1 U625 ( .A(G132), .ZN(G219) );
  INV_X1 U626 ( .A(G57), .ZN(G237) );
  NAND2_X1 U627 ( .A1(n638), .A2(G53), .ZN(n566) );
  NAND2_X1 U628 ( .A1(G65), .A2(n646), .ZN(n565) );
  NAND2_X1 U629 ( .A1(n566), .A2(n565), .ZN(n570) );
  NAND2_X1 U630 ( .A1(G91), .A2(n637), .ZN(n568) );
  NAND2_X1 U631 ( .A1(G78), .A2(n641), .ZN(n567) );
  NAND2_X1 U632 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X1 U633 ( .A1(n570), .A2(n569), .ZN(n696) );
  INV_X1 U634 ( .A(n696), .ZN(G299) );
  NAND2_X1 U635 ( .A1(n638), .A2(G51), .ZN(n571) );
  XNOR2_X1 U636 ( .A(KEYINPUT73), .B(n571), .ZN(n574) );
  NAND2_X1 U637 ( .A1(G63), .A2(n646), .ZN(n572) );
  XOR2_X1 U638 ( .A(KEYINPUT72), .B(n572), .Z(n573) );
  NOR2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(KEYINPUT6), .ZN(n581) );
  NAND2_X1 U641 ( .A1(n637), .A2(G89), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n576), .B(KEYINPUT4), .ZN(n578) );
  NAND2_X1 U643 ( .A1(G76), .A2(n641), .ZN(n577) );
  NAND2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(KEYINPUT5), .B(n579), .ZN(n580) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U648 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U649 ( .A1(G7), .A2(G661), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n583), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U651 ( .A(G223), .ZN(n827) );
  NAND2_X1 U652 ( .A1(n827), .A2(G567), .ZN(n584) );
  XOR2_X1 U653 ( .A(KEYINPUT11), .B(n584), .Z(G234) );
  NAND2_X1 U654 ( .A1(n646), .A2(G56), .ZN(n585) );
  XOR2_X1 U655 ( .A(KEYINPUT14), .B(n585), .Z(n591) );
  NAND2_X1 U656 ( .A1(n637), .A2(G81), .ZN(n586) );
  XNOR2_X1 U657 ( .A(n586), .B(KEYINPUT12), .ZN(n588) );
  NAND2_X1 U658 ( .A1(G68), .A2(n641), .ZN(n587) );
  NAND2_X1 U659 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U660 ( .A(KEYINPUT13), .B(n589), .Z(n590) );
  NOR2_X1 U661 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U662 ( .A1(n638), .A2(G43), .ZN(n592) );
  NAND2_X1 U663 ( .A1(n593), .A2(n592), .ZN(n987) );
  INV_X1 U664 ( .A(G860), .ZN(n607) );
  OR2_X1 U665 ( .A1(n987), .A2(n607), .ZN(G153) );
  XOR2_X1 U666 ( .A(G171), .B(KEYINPUT70), .Z(G301) );
  NAND2_X1 U667 ( .A1(G868), .A2(G301), .ZN(n594) );
  XOR2_X1 U668 ( .A(KEYINPUT71), .B(n594), .Z(n603) );
  NAND2_X1 U669 ( .A1(n637), .A2(G92), .ZN(n596) );
  NAND2_X1 U670 ( .A1(G66), .A2(n646), .ZN(n595) );
  NAND2_X1 U671 ( .A1(n596), .A2(n595), .ZN(n600) );
  NAND2_X1 U672 ( .A1(n638), .A2(G54), .ZN(n598) );
  NAND2_X1 U673 ( .A1(G79), .A2(n641), .ZN(n597) );
  NAND2_X1 U674 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U675 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U676 ( .A(KEYINPUT15), .B(n601), .Z(n971) );
  OR2_X1 U677 ( .A1(n971), .A2(G868), .ZN(n602) );
  NAND2_X1 U678 ( .A1(n603), .A2(n602), .ZN(G284) );
  INV_X1 U679 ( .A(G868), .ZN(n657) );
  NOR2_X1 U680 ( .A1(G286), .A2(n657), .ZN(n604) );
  XNOR2_X1 U681 ( .A(n604), .B(KEYINPUT74), .ZN(n606) );
  NOR2_X1 U682 ( .A1(G299), .A2(G868), .ZN(n605) );
  NOR2_X1 U683 ( .A1(n606), .A2(n605), .ZN(G297) );
  NAND2_X1 U684 ( .A1(n607), .A2(G559), .ZN(n608) );
  NAND2_X1 U685 ( .A1(n608), .A2(n971), .ZN(n609) );
  XNOR2_X1 U686 ( .A(n609), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U687 ( .A1(G868), .A2(n987), .ZN(n612) );
  NAND2_X1 U688 ( .A1(G868), .A2(n971), .ZN(n610) );
  NOR2_X1 U689 ( .A1(G559), .A2(n610), .ZN(n611) );
  NOR2_X1 U690 ( .A1(n612), .A2(n611), .ZN(G282) );
  NAND2_X1 U691 ( .A1(n971), .A2(G559), .ZN(n655) );
  XNOR2_X1 U692 ( .A(n987), .B(n655), .ZN(n613) );
  NOR2_X1 U693 ( .A1(n613), .A2(G860), .ZN(n622) );
  NAND2_X1 U694 ( .A1(G93), .A2(n637), .ZN(n615) );
  NAND2_X1 U695 ( .A1(G55), .A2(n638), .ZN(n614) );
  NAND2_X1 U696 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U697 ( .A1(G80), .A2(n641), .ZN(n616) );
  XNOR2_X1 U698 ( .A(KEYINPUT77), .B(n616), .ZN(n617) );
  NOR2_X1 U699 ( .A1(n618), .A2(n617), .ZN(n620) );
  NAND2_X1 U700 ( .A1(G67), .A2(n646), .ZN(n619) );
  NAND2_X1 U701 ( .A1(n620), .A2(n619), .ZN(n658) );
  XOR2_X1 U702 ( .A(n658), .B(KEYINPUT76), .Z(n621) );
  XNOR2_X1 U703 ( .A(n622), .B(n621), .ZN(G145) );
  NAND2_X1 U704 ( .A1(G62), .A2(n646), .ZN(n624) );
  NAND2_X1 U705 ( .A1(G75), .A2(n641), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U707 ( .A1(n637), .A2(G88), .ZN(n625) );
  XOR2_X1 U708 ( .A(KEYINPUT80), .B(n625), .Z(n626) );
  NOR2_X1 U709 ( .A1(n627), .A2(n626), .ZN(n629) );
  NAND2_X1 U710 ( .A1(n638), .A2(G50), .ZN(n628) );
  NAND2_X1 U711 ( .A1(n629), .A2(n628), .ZN(G303) );
  INV_X1 U712 ( .A(G303), .ZN(G166) );
  NAND2_X1 U713 ( .A1(G74), .A2(G651), .ZN(n630) );
  XNOR2_X1 U714 ( .A(n630), .B(KEYINPUT78), .ZN(n636) );
  NAND2_X1 U715 ( .A1(G49), .A2(n638), .ZN(n633) );
  NAND2_X1 U716 ( .A1(G87), .A2(n631), .ZN(n632) );
  NAND2_X1 U717 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U718 ( .A1(n646), .A2(n634), .ZN(n635) );
  NAND2_X1 U719 ( .A1(n636), .A2(n635), .ZN(G288) );
  NAND2_X1 U720 ( .A1(G86), .A2(n637), .ZN(n640) );
  NAND2_X1 U721 ( .A1(G48), .A2(n638), .ZN(n639) );
  NAND2_X1 U722 ( .A1(n640), .A2(n639), .ZN(n645) );
  NAND2_X1 U723 ( .A1(n641), .A2(G73), .ZN(n642) );
  XNOR2_X1 U724 ( .A(n642), .B(KEYINPUT79), .ZN(n643) );
  XNOR2_X1 U725 ( .A(n643), .B(KEYINPUT2), .ZN(n644) );
  NOR2_X1 U726 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U727 ( .A1(G61), .A2(n646), .ZN(n647) );
  NAND2_X1 U728 ( .A1(n648), .A2(n647), .ZN(G305) );
  XNOR2_X1 U729 ( .A(KEYINPUT19), .B(G290), .ZN(n649) );
  XNOR2_X1 U730 ( .A(n649), .B(G288), .ZN(n650) );
  XNOR2_X1 U731 ( .A(G166), .B(n650), .ZN(n652) );
  XNOR2_X1 U732 ( .A(n987), .B(n696), .ZN(n651) );
  XNOR2_X1 U733 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U734 ( .A(n653), .B(G305), .ZN(n654) );
  XNOR2_X1 U735 ( .A(n654), .B(n658), .ZN(n897) );
  XOR2_X1 U736 ( .A(n897), .B(n655), .Z(n656) );
  NOR2_X1 U737 ( .A1(n657), .A2(n656), .ZN(n660) );
  NOR2_X1 U738 ( .A1(G868), .A2(n658), .ZN(n659) );
  NOR2_X1 U739 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U740 ( .A(KEYINPUT81), .B(n661), .Z(G295) );
  NAND2_X1 U741 ( .A1(G2078), .A2(G2084), .ZN(n662) );
  XOR2_X1 U742 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U743 ( .A1(n663), .A2(G2090), .ZN(n664) );
  XNOR2_X1 U744 ( .A(n664), .B(KEYINPUT21), .ZN(n665) );
  XNOR2_X1 U745 ( .A(KEYINPUT82), .B(n665), .ZN(n666) );
  NAND2_X1 U746 ( .A1(n666), .A2(G2072), .ZN(n667) );
  XOR2_X1 U747 ( .A(KEYINPUT83), .B(n667), .Z(G158) );
  XNOR2_X1 U748 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U749 ( .A(KEYINPUT69), .B(G82), .ZN(G220) );
  NAND2_X1 U750 ( .A1(G120), .A2(G69), .ZN(n668) );
  NOR2_X1 U751 ( .A1(G237), .A2(n668), .ZN(n669) );
  XNOR2_X1 U752 ( .A(KEYINPUT84), .B(n669), .ZN(n670) );
  NAND2_X1 U753 ( .A1(n670), .A2(G108), .ZN(n915) );
  NAND2_X1 U754 ( .A1(n915), .A2(G567), .ZN(n675) );
  NOR2_X1 U755 ( .A1(G219), .A2(G220), .ZN(n671) );
  XOR2_X1 U756 ( .A(KEYINPUT22), .B(n671), .Z(n672) );
  NOR2_X1 U757 ( .A1(G218), .A2(n672), .ZN(n673) );
  NAND2_X1 U758 ( .A1(G96), .A2(n673), .ZN(n916) );
  NAND2_X1 U759 ( .A1(n916), .A2(G2106), .ZN(n674) );
  NAND2_X1 U760 ( .A1(n675), .A2(n674), .ZN(n831) );
  NAND2_X1 U761 ( .A1(G483), .A2(G661), .ZN(n676) );
  NOR2_X1 U762 ( .A1(n831), .A2(n676), .ZN(n830) );
  NAND2_X1 U763 ( .A1(n830), .A2(G36), .ZN(G176) );
  NAND2_X1 U764 ( .A1(G160), .A2(G40), .ZN(n771) );
  INV_X1 U765 ( .A(n771), .ZN(n677) );
  NOR2_X2 U766 ( .A1(G164), .A2(G1384), .ZN(n772) );
  INV_X1 U767 ( .A(n723), .ZN(n704) );
  NAND2_X1 U768 ( .A1(G2072), .A2(n704), .ZN(n679) );
  INV_X1 U769 ( .A(G1956), .ZN(n998) );
  NOR2_X1 U770 ( .A1(n704), .A2(n998), .ZN(n680) );
  NOR2_X1 U771 ( .A1(n681), .A2(n680), .ZN(n697) );
  NOR2_X1 U772 ( .A1(n697), .A2(n696), .ZN(n683) );
  INV_X1 U773 ( .A(KEYINPUT28), .ZN(n682) );
  XNOR2_X1 U774 ( .A(n683), .B(n682), .ZN(n701) );
  INV_X1 U775 ( .A(G1996), .ZN(n945) );
  NOR2_X1 U776 ( .A1(n723), .A2(n945), .ZN(n685) );
  XNOR2_X1 U777 ( .A(n685), .B(n684), .ZN(n687) );
  NAND2_X1 U778 ( .A1(n723), .A2(G1341), .ZN(n686) );
  NAND2_X1 U779 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U780 ( .A1(n987), .A2(n688), .ZN(n693) );
  NAND2_X1 U781 ( .A1(n971), .A2(n693), .ZN(n692) );
  NAND2_X1 U782 ( .A1(G1348), .A2(n723), .ZN(n690) );
  NAND2_X1 U783 ( .A1(n704), .A2(G2067), .ZN(n689) );
  NAND2_X1 U784 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U785 ( .A1(n692), .A2(n691), .ZN(n695) );
  OR2_X1 U786 ( .A1(n971), .A2(n693), .ZN(n694) );
  NAND2_X1 U787 ( .A1(n695), .A2(n694), .ZN(n699) );
  NAND2_X1 U788 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U789 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U790 ( .A1(n701), .A2(n700), .ZN(n703) );
  INV_X1 U791 ( .A(KEYINPUT29), .ZN(n702) );
  XNOR2_X1 U792 ( .A(n703), .B(n702), .ZN(n710) );
  NOR2_X1 U793 ( .A1(n704), .A2(G1961), .ZN(n705) );
  XOR2_X1 U794 ( .A(KEYINPUT94), .B(n705), .Z(n708) );
  XOR2_X1 U795 ( .A(G2078), .B(KEYINPUT25), .Z(n955) );
  NOR2_X1 U796 ( .A1(n955), .A2(n723), .ZN(n706) );
  XNOR2_X1 U797 ( .A(KEYINPUT95), .B(n706), .ZN(n707) );
  NAND2_X1 U798 ( .A1(n708), .A2(n707), .ZN(n716) );
  NAND2_X1 U799 ( .A1(n716), .A2(G171), .ZN(n709) );
  NAND2_X1 U800 ( .A1(n710), .A2(n709), .ZN(n722) );
  NAND2_X1 U801 ( .A1(G8), .A2(n723), .ZN(n766) );
  NOR2_X1 U802 ( .A1(G2084), .A2(n723), .ZN(n733) );
  NOR2_X1 U803 ( .A1(n734), .A2(n733), .ZN(n711) );
  NAND2_X1 U804 ( .A1(G8), .A2(n711), .ZN(n714) );
  INV_X1 U805 ( .A(KEYINPUT30), .ZN(n712) );
  NOR2_X1 U806 ( .A1(G168), .A2(n715), .ZN(n718) );
  NOR2_X1 U807 ( .A1(G171), .A2(n716), .ZN(n717) );
  INV_X1 U808 ( .A(KEYINPUT31), .ZN(n719) );
  XNOR2_X1 U809 ( .A(n720), .B(n719), .ZN(n721) );
  NAND2_X1 U810 ( .A1(n722), .A2(n721), .ZN(n737) );
  NAND2_X1 U811 ( .A1(n737), .A2(G286), .ZN(n730) );
  INV_X1 U812 ( .A(G8), .ZN(n728) );
  NOR2_X1 U813 ( .A1(G1971), .A2(n766), .ZN(n725) );
  NOR2_X1 U814 ( .A1(G2090), .A2(n723), .ZN(n724) );
  NOR2_X1 U815 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U816 ( .A1(n726), .A2(G303), .ZN(n727) );
  OR2_X1 U817 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U818 ( .A1(n730), .A2(n729), .ZN(n732) );
  INV_X1 U819 ( .A(KEYINPUT32), .ZN(n731) );
  XNOR2_X1 U820 ( .A(n732), .B(n731), .ZN(n756) );
  AND2_X1 U821 ( .A1(G8), .A2(n733), .ZN(n735) );
  NOR2_X1 U822 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U823 ( .A1(n737), .A2(n736), .ZN(n757) );
  NAND2_X1 U824 ( .A1(G1976), .A2(G288), .ZN(n977) );
  AND2_X1 U825 ( .A1(n757), .A2(n977), .ZN(n738) );
  NAND2_X1 U826 ( .A1(n756), .A2(n738), .ZN(n744) );
  INV_X1 U827 ( .A(n977), .ZN(n741) );
  NOR2_X1 U828 ( .A1(G1976), .A2(G288), .ZN(n975) );
  NOR2_X1 U829 ( .A1(G1971), .A2(G303), .ZN(n739) );
  NOR2_X1 U830 ( .A1(n975), .A2(n739), .ZN(n740) );
  OR2_X1 U831 ( .A1(n741), .A2(n740), .ZN(n742) );
  OR2_X1 U832 ( .A1(n766), .A2(n742), .ZN(n743) );
  NAND2_X1 U833 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U834 ( .A(n745), .B(KEYINPUT64), .ZN(n746) );
  NOR2_X1 U835 ( .A1(KEYINPUT33), .A2(n746), .ZN(n751) );
  NAND2_X1 U836 ( .A1(KEYINPUT33), .A2(n975), .ZN(n747) );
  XNOR2_X1 U837 ( .A(KEYINPUT98), .B(n747), .ZN(n748) );
  NOR2_X1 U838 ( .A1(n766), .A2(n748), .ZN(n749) );
  XOR2_X1 U839 ( .A(KEYINPUT99), .B(n749), .Z(n750) );
  NOR2_X1 U840 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U841 ( .A(KEYINPUT100), .B(n752), .ZN(n754) );
  XNOR2_X1 U842 ( .A(G1981), .B(KEYINPUT101), .ZN(n753) );
  XNOR2_X1 U843 ( .A(n753), .B(G305), .ZN(n988) );
  NAND2_X1 U844 ( .A1(n754), .A2(n988), .ZN(n755) );
  XNOR2_X1 U845 ( .A(n755), .B(KEYINPUT102), .ZN(n770) );
  NAND2_X1 U846 ( .A1(n757), .A2(n756), .ZN(n760) );
  NOR2_X1 U847 ( .A1(G2090), .A2(G303), .ZN(n758) );
  NAND2_X1 U848 ( .A1(G8), .A2(n758), .ZN(n759) );
  NAND2_X1 U849 ( .A1(n760), .A2(n759), .ZN(n761) );
  AND2_X1 U850 ( .A1(n761), .A2(n766), .ZN(n768) );
  XNOR2_X1 U851 ( .A(KEYINPUT24), .B(KEYINPUT93), .ZN(n762) );
  XNOR2_X1 U852 ( .A(n762), .B(KEYINPUT92), .ZN(n764) );
  NOR2_X1 U853 ( .A1(G1981), .A2(G305), .ZN(n763) );
  XNOR2_X1 U854 ( .A(n764), .B(n763), .ZN(n765) );
  NOR2_X1 U855 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U856 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U857 ( .A1(n770), .A2(n769), .ZN(n808) );
  NOR2_X1 U858 ( .A1(n772), .A2(n771), .ZN(n822) );
  XNOR2_X1 U859 ( .A(KEYINPUT86), .B(KEYINPUT34), .ZN(n776) );
  NAND2_X1 U860 ( .A1(G140), .A2(n872), .ZN(n774) );
  NAND2_X1 U861 ( .A1(G104), .A2(n873), .ZN(n773) );
  NAND2_X1 U862 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U863 ( .A(n776), .B(n775), .ZN(n782) );
  NAND2_X1 U864 ( .A1(n876), .A2(G128), .ZN(n777) );
  XOR2_X1 U865 ( .A(KEYINPUT87), .B(n777), .Z(n779) );
  NAND2_X1 U866 ( .A1(n877), .A2(G116), .ZN(n778) );
  NAND2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U868 ( .A(KEYINPUT35), .B(n780), .Z(n781) );
  NOR2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n783) );
  XOR2_X1 U870 ( .A(KEYINPUT36), .B(n783), .Z(n894) );
  XOR2_X1 U871 ( .A(KEYINPUT37), .B(G2067), .Z(n819) );
  AND2_X1 U872 ( .A1(n894), .A2(n819), .ZN(n922) );
  NAND2_X1 U873 ( .A1(n822), .A2(n922), .ZN(n816) );
  INV_X1 U874 ( .A(n816), .ZN(n803) );
  XOR2_X1 U875 ( .A(KEYINPUT38), .B(KEYINPUT88), .Z(n785) );
  NAND2_X1 U876 ( .A1(G105), .A2(n873), .ZN(n784) );
  XNOR2_X1 U877 ( .A(n785), .B(n784), .ZN(n789) );
  NAND2_X1 U878 ( .A1(G129), .A2(n876), .ZN(n787) );
  NAND2_X1 U879 ( .A1(G141), .A2(n872), .ZN(n786) );
  NAND2_X1 U880 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U881 ( .A1(n789), .A2(n788), .ZN(n791) );
  NAND2_X1 U882 ( .A1(n877), .A2(G117), .ZN(n790) );
  NAND2_X1 U883 ( .A1(n791), .A2(n790), .ZN(n862) );
  NAND2_X1 U884 ( .A1(G1996), .A2(n862), .ZN(n792) );
  XNOR2_X1 U885 ( .A(n792), .B(KEYINPUT89), .ZN(n800) );
  INV_X1 U886 ( .A(G1991), .ZN(n809) );
  NAND2_X1 U887 ( .A1(G131), .A2(n872), .ZN(n794) );
  NAND2_X1 U888 ( .A1(G95), .A2(n873), .ZN(n793) );
  NAND2_X1 U889 ( .A1(n794), .A2(n793), .ZN(n798) );
  NAND2_X1 U890 ( .A1(G119), .A2(n876), .ZN(n796) );
  NAND2_X1 U891 ( .A1(G107), .A2(n877), .ZN(n795) );
  NAND2_X1 U892 ( .A1(n796), .A2(n795), .ZN(n797) );
  NOR2_X1 U893 ( .A1(n798), .A2(n797), .ZN(n891) );
  NOR2_X1 U894 ( .A1(n809), .A2(n891), .ZN(n799) );
  NOR2_X1 U895 ( .A1(n800), .A2(n799), .ZN(n927) );
  INV_X1 U896 ( .A(n822), .ZN(n801) );
  NOR2_X1 U897 ( .A1(n927), .A2(n801), .ZN(n812) );
  XNOR2_X1 U898 ( .A(KEYINPUT90), .B(n812), .ZN(n802) );
  NOR2_X1 U899 ( .A1(n803), .A2(n802), .ZN(n804) );
  XOR2_X1 U900 ( .A(n804), .B(KEYINPUT91), .Z(n806) );
  XNOR2_X1 U901 ( .A(G1986), .B(G290), .ZN(n982) );
  NAND2_X1 U902 ( .A1(n982), .A2(n822), .ZN(n805) );
  AND2_X1 U903 ( .A1(n806), .A2(n805), .ZN(n807) );
  NAND2_X1 U904 ( .A1(n808), .A2(n807), .ZN(n825) );
  NOR2_X1 U905 ( .A1(G1996), .A2(n862), .ZN(n919) );
  AND2_X1 U906 ( .A1(n809), .A2(n891), .ZN(n929) );
  NOR2_X1 U907 ( .A1(G1986), .A2(G290), .ZN(n810) );
  NOR2_X1 U908 ( .A1(n929), .A2(n810), .ZN(n811) );
  NOR2_X1 U909 ( .A1(n812), .A2(n811), .ZN(n813) );
  NOR2_X1 U910 ( .A1(n919), .A2(n813), .ZN(n815) );
  XOR2_X1 U911 ( .A(KEYINPUT39), .B(KEYINPUT103), .Z(n814) );
  XNOR2_X1 U912 ( .A(n815), .B(n814), .ZN(n817) );
  NAND2_X1 U913 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U914 ( .A(n818), .B(KEYINPUT104), .ZN(n821) );
  NOR2_X1 U915 ( .A1(n894), .A2(n819), .ZN(n820) );
  XNOR2_X1 U916 ( .A(KEYINPUT105), .B(n820), .ZN(n936) );
  NAND2_X1 U917 ( .A1(n821), .A2(n936), .ZN(n823) );
  NAND2_X1 U918 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U919 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U920 ( .A(n826), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n827), .ZN(G217) );
  AND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n828) );
  NAND2_X1 U923 ( .A1(G661), .A2(n828), .ZN(G259) );
  NAND2_X1 U924 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U925 ( .A1(n830), .A2(n829), .ZN(G188) );
  INV_X1 U926 ( .A(n831), .ZN(G319) );
  XOR2_X1 U927 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n833) );
  XNOR2_X1 U928 ( .A(KEYINPUT106), .B(G2096), .ZN(n832) );
  XNOR2_X1 U929 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U930 ( .A(n834), .B(G2678), .Z(n836) );
  XNOR2_X1 U931 ( .A(G2067), .B(G2078), .ZN(n835) );
  XNOR2_X1 U932 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U933 ( .A(G2100), .B(G2090), .Z(n838) );
  XNOR2_X1 U934 ( .A(G2072), .B(G2084), .ZN(n837) );
  XNOR2_X1 U935 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U936 ( .A(n840), .B(n839), .Z(n842) );
  XNOR2_X1 U937 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n841) );
  XNOR2_X1 U938 ( .A(n842), .B(n841), .ZN(G227) );
  XOR2_X1 U939 ( .A(G1976), .B(G1956), .Z(n844) );
  XNOR2_X1 U940 ( .A(G1986), .B(G1961), .ZN(n843) );
  XNOR2_X1 U941 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U942 ( .A(G1981), .B(G1966), .Z(n846) );
  XNOR2_X1 U943 ( .A(G1996), .B(G1991), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U945 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U946 ( .A(KEYINPUT109), .B(G2474), .ZN(n849) );
  XNOR2_X1 U947 ( .A(n850), .B(n849), .ZN(n852) );
  XOR2_X1 U948 ( .A(G1971), .B(KEYINPUT41), .Z(n851) );
  XNOR2_X1 U949 ( .A(n852), .B(n851), .ZN(G229) );
  NAND2_X1 U950 ( .A1(G124), .A2(n876), .ZN(n853) );
  XNOR2_X1 U951 ( .A(n853), .B(KEYINPUT110), .ZN(n854) );
  XNOR2_X1 U952 ( .A(n854), .B(KEYINPUT44), .ZN(n856) );
  NAND2_X1 U953 ( .A1(G112), .A2(n877), .ZN(n855) );
  NAND2_X1 U954 ( .A1(n856), .A2(n855), .ZN(n860) );
  NAND2_X1 U955 ( .A1(G136), .A2(n872), .ZN(n858) );
  NAND2_X1 U956 ( .A1(G100), .A2(n873), .ZN(n857) );
  NAND2_X1 U957 ( .A1(n858), .A2(n857), .ZN(n859) );
  NOR2_X1 U958 ( .A1(n860), .A2(n859), .ZN(G162) );
  XOR2_X1 U959 ( .A(G162), .B(n925), .Z(n861) );
  XNOR2_X1 U960 ( .A(n862), .B(n861), .ZN(n871) );
  NAND2_X1 U961 ( .A1(G130), .A2(n876), .ZN(n864) );
  NAND2_X1 U962 ( .A1(G118), .A2(n877), .ZN(n863) );
  NAND2_X1 U963 ( .A1(n864), .A2(n863), .ZN(n869) );
  NAND2_X1 U964 ( .A1(G142), .A2(n872), .ZN(n866) );
  NAND2_X1 U965 ( .A1(G106), .A2(n873), .ZN(n865) );
  NAND2_X1 U966 ( .A1(n866), .A2(n865), .ZN(n867) );
  XOR2_X1 U967 ( .A(KEYINPUT45), .B(n867), .Z(n868) );
  NOR2_X1 U968 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U969 ( .A(n871), .B(n870), .Z(n886) );
  NAND2_X1 U970 ( .A1(G139), .A2(n872), .ZN(n875) );
  NAND2_X1 U971 ( .A1(G103), .A2(n873), .ZN(n874) );
  NAND2_X1 U972 ( .A1(n875), .A2(n874), .ZN(n884) );
  XNOR2_X1 U973 ( .A(KEYINPUT47), .B(KEYINPUT112), .ZN(n882) );
  NAND2_X1 U974 ( .A1(n876), .A2(G127), .ZN(n880) );
  NAND2_X1 U975 ( .A1(n877), .A2(G115), .ZN(n878) );
  XOR2_X1 U976 ( .A(KEYINPUT111), .B(n878), .Z(n879) );
  NAND2_X1 U977 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U978 ( .A(n882), .B(n881), .Z(n883) );
  NOR2_X1 U979 ( .A1(n884), .A2(n883), .ZN(n932) );
  XNOR2_X1 U980 ( .A(G160), .B(n932), .ZN(n885) );
  XNOR2_X1 U981 ( .A(n886), .B(n885), .ZN(n890) );
  XOR2_X1 U982 ( .A(KEYINPUT46), .B(KEYINPUT113), .Z(n888) );
  XNOR2_X1 U983 ( .A(KEYINPUT114), .B(KEYINPUT48), .ZN(n887) );
  XNOR2_X1 U984 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U985 ( .A(n890), .B(n889), .Z(n893) );
  XNOR2_X1 U986 ( .A(G164), .B(n891), .ZN(n892) );
  XNOR2_X1 U987 ( .A(n893), .B(n892), .ZN(n895) );
  XOR2_X1 U988 ( .A(n895), .B(n894), .Z(n896) );
  NOR2_X1 U989 ( .A1(G37), .A2(n896), .ZN(G395) );
  XNOR2_X1 U990 ( .A(n971), .B(G286), .ZN(n898) );
  XNOR2_X1 U991 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U992 ( .A(n899), .B(G171), .ZN(n900) );
  NOR2_X1 U993 ( .A1(G37), .A2(n900), .ZN(G397) );
  XOR2_X1 U994 ( .A(G2451), .B(G2430), .Z(n902) );
  XNOR2_X1 U995 ( .A(G2438), .B(G2443), .ZN(n901) );
  XNOR2_X1 U996 ( .A(n902), .B(n901), .ZN(n908) );
  XOR2_X1 U997 ( .A(G2435), .B(G2454), .Z(n904) );
  XNOR2_X1 U998 ( .A(G1348), .B(G1341), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n904), .B(n903), .ZN(n906) );
  XOR2_X1 U1000 ( .A(G2446), .B(G2427), .Z(n905) );
  XNOR2_X1 U1001 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1002 ( .A(n908), .B(n907), .Z(n909) );
  NAND2_X1 U1003 ( .A1(G14), .A2(n909), .ZN(n917) );
  NAND2_X1 U1004 ( .A1(G319), .A2(n917), .ZN(n912) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n910) );
  XNOR2_X1 U1006 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1007 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1009 ( .A1(n914), .A2(n913), .ZN(G225) );
  XNOR2_X1 U1010 ( .A(KEYINPUT115), .B(G225), .ZN(G308) );
  INV_X1 U1012 ( .A(G120), .ZN(G236) );
  INV_X1 U1013 ( .A(G108), .ZN(G238) );
  INV_X1 U1014 ( .A(G96), .ZN(G221) );
  INV_X1 U1015 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1016 ( .A1(n916), .A2(n915), .ZN(G325) );
  INV_X1 U1017 ( .A(G325), .ZN(G261) );
  INV_X1 U1018 ( .A(n917), .ZN(G401) );
  XOR2_X1 U1019 ( .A(G2090), .B(G162), .Z(n918) );
  NOR2_X1 U1020 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1021 ( .A(n920), .B(KEYINPUT51), .ZN(n921) );
  NOR2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n931) );
  XOR2_X1 U1023 ( .A(G2084), .B(G160), .Z(n923) );
  XNOR2_X1 U1024 ( .A(KEYINPUT116), .B(n923), .ZN(n924) );
  NOR2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n928) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n939) );
  XOR2_X1 U1029 ( .A(G2072), .B(n932), .Z(n934) );
  XOR2_X1 U1030 ( .A(G164), .B(G2078), .Z(n933) );
  NOR2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1032 ( .A(n935), .B(KEYINPUT50), .ZN(n937) );
  NAND2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1035 ( .A(KEYINPUT52), .B(n940), .Z(n941) );
  NOR2_X1 U1036 ( .A1(KEYINPUT55), .A2(n941), .ZN(n942) );
  XNOR2_X1 U1037 ( .A(KEYINPUT117), .B(n942), .ZN(n943) );
  NAND2_X1 U1038 ( .A1(n943), .A2(G29), .ZN(n1026) );
  XOR2_X1 U1039 ( .A(KEYINPUT53), .B(KEYINPUT123), .Z(n960) );
  XNOR2_X1 U1040 ( .A(KEYINPUT119), .B(G1991), .ZN(n944) );
  XNOR2_X1 U1041 ( .A(n944), .B(G25), .ZN(n951) );
  XNOR2_X1 U1042 ( .A(G32), .B(n945), .ZN(n946) );
  NAND2_X1 U1043 ( .A1(n946), .A2(G28), .ZN(n949) );
  XOR2_X1 U1044 ( .A(KEYINPUT121), .B(G2072), .Z(n947) );
  XNOR2_X1 U1045 ( .A(G33), .B(n947), .ZN(n948) );
  NOR2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(KEYINPUT120), .B(G2067), .ZN(n952) );
  XNOR2_X1 U1049 ( .A(G26), .B(n952), .ZN(n953) );
  NOR2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n958) );
  XOR2_X1 U1051 ( .A(n955), .B(G27), .Z(n956) );
  XNOR2_X1 U1052 ( .A(KEYINPUT122), .B(n956), .ZN(n957) );
  NAND2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(n960), .B(n959), .ZN(n963) );
  XOR2_X1 U1055 ( .A(G2084), .B(G34), .Z(n961) );
  XNOR2_X1 U1056 ( .A(KEYINPUT54), .B(n961), .ZN(n962) );
  NAND2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(KEYINPUT118), .B(G2090), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(G35), .B(n964), .ZN(n965) );
  NOR2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1061 ( .A(KEYINPUT55), .B(n967), .Z(n968) );
  NOR2_X1 U1062 ( .A1(G29), .A2(n968), .ZN(n969) );
  XOR2_X1 U1063 ( .A(KEYINPUT124), .B(n969), .Z(n970) );
  NAND2_X1 U1064 ( .A1(G11), .A2(n970), .ZN(n1024) );
  XNOR2_X1 U1065 ( .A(G16), .B(KEYINPUT56), .ZN(n997) );
  XNOR2_X1 U1066 ( .A(G1348), .B(n971), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(G171), .B(G1961), .ZN(n972) );
  NAND2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n986) );
  XNOR2_X1 U1069 ( .A(G1971), .B(G166), .ZN(n974) );
  XNOR2_X1 U1070 ( .A(n974), .B(KEYINPUT126), .ZN(n981) );
  INV_X1 U1071 ( .A(n975), .ZN(n976) );
  NAND2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(G1956), .B(G299), .ZN(n978) );
  NOR2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1077 ( .A(KEYINPUT127), .B(n984), .ZN(n985) );
  NOR2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n995) );
  XNOR2_X1 U1079 ( .A(n987), .B(G1341), .ZN(n993) );
  XNOR2_X1 U1080 ( .A(G1966), .B(G168), .ZN(n989) );
  NAND2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1082 ( .A(n990), .B(KEYINPUT57), .ZN(n991) );
  XNOR2_X1 U1083 ( .A(KEYINPUT125), .B(n991), .ZN(n992) );
  NOR2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n1022) );
  INV_X1 U1087 ( .A(G16), .ZN(n1020) );
  XNOR2_X1 U1088 ( .A(G20), .B(n998), .ZN(n1002) );
  XNOR2_X1 U1089 ( .A(G1341), .B(G19), .ZN(n1000) );
  XNOR2_X1 U1090 ( .A(G6), .B(G1981), .ZN(n999) );
  NOR2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XOR2_X1 U1093 ( .A(KEYINPUT59), .B(G1348), .Z(n1003) );
  XNOR2_X1 U1094 ( .A(G4), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1096 ( .A(KEYINPUT60), .B(n1006), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(G1966), .B(G21), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(G5), .B(G1961), .ZN(n1007) );
  NOR2_X1 U1099 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1017) );
  XNOR2_X1 U1101 ( .A(G1971), .B(G22), .ZN(n1012) );
  XNOR2_X1 U1102 ( .A(G23), .B(G1976), .ZN(n1011) );
  NOR2_X1 U1103 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XOR2_X1 U1104 ( .A(G1986), .B(G24), .Z(n1013) );
  NAND2_X1 U1105 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1106 ( .A(KEYINPUT58), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1108 ( .A(KEYINPUT61), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1109 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1113 ( .A(KEYINPUT62), .B(n1027), .Z(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

