

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592;

  XOR2_X1 U324 ( .A(n453), .B(n452), .Z(n571) );
  XNOR2_X2 U325 ( .A(n368), .B(n367), .ZN(n404) );
  XNOR2_X1 U326 ( .A(n438), .B(n296), .ZN(n390) );
  XNOR2_X1 U327 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U328 ( .A(n476), .B(KEYINPUT120), .ZN(n477) );
  NOR2_X1 U329 ( .A1(n572), .A2(n483), .ZN(n569) );
  NAND2_X1 U330 ( .A1(n571), .A2(n404), .ZN(n292) );
  XNOR2_X1 U331 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n293) );
  XOR2_X1 U332 ( .A(KEYINPUT81), .B(G211GAT), .Z(n294) );
  AND2_X1 U333 ( .A1(n431), .A2(n430), .ZN(n295) );
  AND2_X1 U334 ( .A1(G226GAT), .A2(G233GAT), .ZN(n296) );
  INV_X1 U335 ( .A(n555), .ZN(n430) );
  XNOR2_X1 U336 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U337 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U338 ( .A(n400), .B(n332), .ZN(n333) );
  XNOR2_X1 U339 ( .A(n399), .B(n398), .ZN(n403) );
  XNOR2_X1 U340 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U341 ( .A(n487), .B(n293), .ZN(n488) );
  XNOR2_X1 U342 ( .A(n459), .B(G43GAT), .ZN(n460) );
  XNOR2_X1 U343 ( .A(n489), .B(n488), .ZN(G1349GAT) );
  XNOR2_X1 U344 ( .A(n461), .B(n460), .ZN(G1330GAT) );
  XOR2_X1 U345 ( .A(KEYINPUT38), .B(KEYINPUT100), .Z(n457) );
  XNOR2_X1 U346 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n297) );
  XNOR2_X1 U347 ( .A(n297), .B(G29GAT), .ZN(n298) );
  XOR2_X1 U348 ( .A(n298), .B(KEYINPUT7), .Z(n300) );
  XNOR2_X1 U349 ( .A(G43GAT), .B(G50GAT), .ZN(n299) );
  XNOR2_X1 U350 ( .A(n300), .B(n299), .ZN(n451) );
  XOR2_X1 U351 ( .A(KEYINPUT71), .B(G197GAT), .Z(n302) );
  XNOR2_X1 U352 ( .A(G169GAT), .B(G113GAT), .ZN(n301) );
  XNOR2_X1 U353 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U354 ( .A(G8GAT), .B(KEYINPUT66), .Z(n304) );
  XNOR2_X1 U355 ( .A(KEYINPUT69), .B(KEYINPUT68), .ZN(n303) );
  XNOR2_X1 U356 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U357 ( .A(n306), .B(n305), .Z(n316) );
  XOR2_X1 U358 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n308) );
  XNOR2_X1 U359 ( .A(KEYINPUT29), .B(KEYINPUT70), .ZN(n307) );
  XNOR2_X1 U360 ( .A(n308), .B(n307), .ZN(n314) );
  XOR2_X1 U361 ( .A(G141GAT), .B(G22GAT), .Z(n371) );
  XOR2_X1 U362 ( .A(KEYINPUT72), .B(KEYINPUT73), .Z(n310) );
  XNOR2_X1 U363 ( .A(G15GAT), .B(G1GAT), .ZN(n309) );
  XNOR2_X1 U364 ( .A(n310), .B(n309), .ZN(n347) );
  XOR2_X1 U365 ( .A(n371), .B(n347), .Z(n312) );
  NAND2_X1 U366 ( .A1(G229GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U367 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U368 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U369 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n451), .B(n317), .ZN(n578) );
  XNOR2_X1 U371 ( .A(KEYINPUT74), .B(n578), .ZN(n535) );
  XOR2_X1 U372 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n319) );
  XNOR2_X1 U373 ( .A(KEYINPUT76), .B(KEYINPUT31), .ZN(n318) );
  XOR2_X1 U374 ( .A(n319), .B(n318), .Z(n336) );
  XOR2_X1 U375 ( .A(G204GAT), .B(G148GAT), .Z(n370) );
  XNOR2_X1 U376 ( .A(G71GAT), .B(G57GAT), .ZN(n320) );
  XNOR2_X1 U377 ( .A(n320), .B(KEYINPUT13), .ZN(n346) );
  XNOR2_X1 U378 ( .A(n370), .B(n346), .ZN(n321) );
  AND2_X1 U379 ( .A1(G230GAT), .A2(G233GAT), .ZN(n322) );
  NAND2_X1 U380 ( .A1(n321), .A2(n322), .ZN(n326) );
  INV_X1 U381 ( .A(n321), .ZN(n324) );
  INV_X1 U382 ( .A(n322), .ZN(n323) );
  NAND2_X1 U383 ( .A1(n324), .A2(n323), .ZN(n325) );
  NAND2_X1 U384 ( .A1(n326), .A2(n325), .ZN(n327) );
  XOR2_X1 U385 ( .A(n327), .B(KEYINPUT77), .Z(n331) );
  XOR2_X1 U386 ( .A(G92GAT), .B(G85GAT), .Z(n329) );
  XNOR2_X1 U387 ( .A(G99GAT), .B(G106GAT), .ZN(n328) );
  XNOR2_X1 U388 ( .A(n329), .B(n328), .ZN(n448) );
  XNOR2_X1 U389 ( .A(n448), .B(KEYINPUT75), .ZN(n330) );
  XNOR2_X1 U390 ( .A(n331), .B(n330), .ZN(n334) );
  XOR2_X1 U391 ( .A(G176GAT), .B(G64GAT), .Z(n400) );
  XOR2_X1 U392 ( .A(G120GAT), .B(G78GAT), .Z(n332) );
  XNOR2_X1 U393 ( .A(n336), .B(n335), .ZN(n583) );
  NOR2_X1 U394 ( .A1(n535), .A2(n583), .ZN(n493) );
  XOR2_X1 U395 ( .A(KEYINPUT83), .B(G64GAT), .Z(n338) );
  XNOR2_X1 U396 ( .A(G22GAT), .B(G127GAT), .ZN(n337) );
  XNOR2_X1 U397 ( .A(n338), .B(n337), .ZN(n351) );
  XNOR2_X1 U398 ( .A(G8GAT), .B(G183GAT), .ZN(n339) );
  XNOR2_X1 U399 ( .A(n294), .B(n339), .ZN(n391) );
  XOR2_X1 U400 ( .A(G155GAT), .B(G78GAT), .Z(n369) );
  XOR2_X1 U401 ( .A(n391), .B(n369), .Z(n341) );
  NAND2_X1 U402 ( .A1(G231GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U403 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U404 ( .A(KEYINPUT82), .B(KEYINPUT12), .Z(n343) );
  XNOR2_X1 U405 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n342) );
  XNOR2_X1 U406 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U407 ( .A(n345), .B(n344), .Z(n349) );
  XNOR2_X1 U408 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U409 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U410 ( .A(n351), .B(n350), .ZN(n587) );
  XNOR2_X1 U411 ( .A(KEYINPUT94), .B(KEYINPUT26), .ZN(n388) );
  XOR2_X1 U412 ( .A(G71GAT), .B(G176GAT), .Z(n358) );
  XOR2_X1 U413 ( .A(G190GAT), .B(G99GAT), .Z(n353) );
  NAND2_X1 U414 ( .A1(G227GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U415 ( .A(n353), .B(n352), .ZN(n356) );
  XOR2_X1 U416 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n355) );
  XNOR2_X1 U417 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n354) );
  XNOR2_X1 U418 ( .A(n355), .B(n354), .ZN(n393) );
  XNOR2_X1 U419 ( .A(n356), .B(n393), .ZN(n357) );
  XNOR2_X1 U420 ( .A(n358), .B(n357), .ZN(n368) );
  XOR2_X1 U421 ( .A(KEYINPUT0), .B(KEYINPUT85), .Z(n360) );
  XNOR2_X1 U422 ( .A(G134GAT), .B(KEYINPUT84), .ZN(n359) );
  XNOR2_X1 U423 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U424 ( .A(n361), .B(G127GAT), .Z(n363) );
  XNOR2_X1 U425 ( .A(G113GAT), .B(G120GAT), .ZN(n362) );
  XNOR2_X1 U426 ( .A(n363), .B(n362), .ZN(n415) );
  XOR2_X1 U427 ( .A(G183GAT), .B(KEYINPUT20), .Z(n365) );
  XNOR2_X1 U428 ( .A(G43GAT), .B(G15GAT), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U430 ( .A(n415), .B(n366), .ZN(n367) );
  XOR2_X1 U431 ( .A(n370), .B(n369), .Z(n373) );
  XOR2_X1 U432 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n425) );
  XNOR2_X1 U433 ( .A(n371), .B(n425), .ZN(n372) );
  XOR2_X1 U434 ( .A(n373), .B(n372), .Z(n386) );
  XOR2_X1 U435 ( .A(G197GAT), .B(KEYINPUT21), .Z(n401) );
  XOR2_X1 U436 ( .A(n401), .B(G211GAT), .Z(n375) );
  NAND2_X1 U437 ( .A1(G228GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U438 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U439 ( .A(KEYINPUT78), .B(G162GAT), .Z(n439) );
  XOR2_X1 U440 ( .A(n376), .B(n439), .Z(n384) );
  XOR2_X1 U441 ( .A(KEYINPUT86), .B(G106GAT), .Z(n378) );
  XNOR2_X1 U442 ( .A(G50GAT), .B(G218GAT), .ZN(n377) );
  XNOR2_X1 U443 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U444 ( .A(KEYINPUT22), .B(KEYINPUT87), .Z(n380) );
  XNOR2_X1 U445 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n379) );
  XNOR2_X1 U446 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U447 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U448 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U449 ( .A(n386), .B(n385), .ZN(n480) );
  NOR2_X1 U450 ( .A1(n404), .A2(n480), .ZN(n387) );
  XNOR2_X1 U451 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U452 ( .A(KEYINPUT93), .B(n389), .Z(n576) );
  XOR2_X1 U453 ( .A(G190GAT), .B(G218GAT), .Z(n438) );
  XOR2_X1 U454 ( .A(n392), .B(KEYINPUT90), .Z(n399) );
  XNOR2_X1 U455 ( .A(n393), .B(KEYINPUT91), .ZN(n397) );
  XOR2_X1 U456 ( .A(KEYINPUT92), .B(G92GAT), .Z(n395) );
  XNOR2_X1 U457 ( .A(G36GAT), .B(G204GAT), .ZN(n394) );
  XNOR2_X1 U458 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U459 ( .A(n401), .B(n400), .Z(n402) );
  XNOR2_X1 U460 ( .A(n403), .B(n402), .ZN(n497) );
  XOR2_X1 U461 ( .A(n497), .B(KEYINPUT27), .Z(n432) );
  NAND2_X1 U462 ( .A1(n576), .A2(n432), .ZN(n552) );
  XNOR2_X1 U463 ( .A(KEYINPUT95), .B(n552), .ZN(n410) );
  INV_X1 U464 ( .A(n480), .ZN(n406) );
  INV_X1 U465 ( .A(n404), .ZN(n483) );
  NOR2_X1 U466 ( .A1(n497), .A2(n483), .ZN(n405) );
  NOR2_X1 U467 ( .A1(n406), .A2(n405), .ZN(n407) );
  XOR2_X1 U468 ( .A(KEYINPUT96), .B(n407), .Z(n408) );
  XNOR2_X1 U469 ( .A(KEYINPUT25), .B(n408), .ZN(n409) );
  NOR2_X1 U470 ( .A1(n410), .A2(n409), .ZN(n411) );
  XNOR2_X1 U471 ( .A(n411), .B(KEYINPUT97), .ZN(n431) );
  XOR2_X1 U472 ( .A(G57GAT), .B(KEYINPUT89), .Z(n413) );
  XNOR2_X1 U473 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n412) );
  XNOR2_X1 U474 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U475 ( .A(n415), .B(n414), .ZN(n429) );
  XOR2_X1 U476 ( .A(G85GAT), .B(G155GAT), .Z(n417) );
  XNOR2_X1 U477 ( .A(G29GAT), .B(G162GAT), .ZN(n416) );
  XNOR2_X1 U478 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U479 ( .A(KEYINPUT88), .B(G148GAT), .Z(n419) );
  XNOR2_X1 U480 ( .A(G141GAT), .B(G1GAT), .ZN(n418) );
  XNOR2_X1 U481 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U482 ( .A(n421), .B(n420), .Z(n427) );
  XOR2_X1 U483 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n423) );
  NAND2_X1 U484 ( .A1(G225GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U485 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U486 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U487 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U488 ( .A(n429), .B(n428), .ZN(n555) );
  XOR2_X1 U489 ( .A(n480), .B(KEYINPUT28), .Z(n531) );
  INV_X1 U490 ( .A(n432), .ZN(n433) );
  NOR2_X1 U491 ( .A1(n531), .A2(n433), .ZN(n434) );
  NAND2_X1 U492 ( .A1(n555), .A2(n434), .ZN(n536) );
  NOR2_X1 U493 ( .A1(n404), .A2(n536), .ZN(n435) );
  NOR2_X1 U494 ( .A1(n295), .A2(n435), .ZN(n492) );
  XOR2_X1 U495 ( .A(KEYINPUT79), .B(KEYINPUT64), .Z(n437) );
  XNOR2_X1 U496 ( .A(KEYINPUT9), .B(KEYINPUT80), .ZN(n436) );
  XNOR2_X1 U497 ( .A(n437), .B(n436), .ZN(n443) );
  XOR2_X1 U498 ( .A(KEYINPUT65), .B(KEYINPUT11), .Z(n441) );
  XNOR2_X1 U499 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U500 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U501 ( .A(n443), .B(n442), .Z(n445) );
  NAND2_X1 U502 ( .A1(G232GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U503 ( .A(n445), .B(n444), .ZN(n447) );
  INV_X1 U504 ( .A(KEYINPUT10), .ZN(n446) );
  XNOR2_X1 U505 ( .A(n447), .B(n446), .ZN(n450) );
  XNOR2_X1 U506 ( .A(G134GAT), .B(n448), .ZN(n449) );
  XNOR2_X1 U507 ( .A(n450), .B(n449), .ZN(n453) );
  INV_X1 U508 ( .A(n451), .ZN(n452) );
  INV_X1 U509 ( .A(n571), .ZN(n564) );
  XNOR2_X1 U510 ( .A(n564), .B(KEYINPUT36), .ZN(n590) );
  NOR2_X1 U511 ( .A1(n492), .A2(n590), .ZN(n454) );
  NAND2_X1 U512 ( .A1(n587), .A2(n454), .ZN(n455) );
  XNOR2_X1 U513 ( .A(n455), .B(KEYINPUT37), .ZN(n523) );
  NAND2_X1 U514 ( .A1(n493), .A2(n523), .ZN(n456) );
  XNOR2_X1 U515 ( .A(n457), .B(n456), .ZN(n458) );
  XOR2_X1 U516 ( .A(KEYINPUT101), .B(n458), .Z(n508) );
  NAND2_X1 U517 ( .A1(n508), .A2(n404), .ZN(n461) );
  XOR2_X1 U518 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n459) );
  XNOR2_X1 U519 ( .A(n583), .B(KEYINPUT41), .ZN(n484) );
  NOR2_X1 U520 ( .A1(n484), .A2(n578), .ZN(n463) );
  XOR2_X1 U521 ( .A(KEYINPUT46), .B(KEYINPUT110), .Z(n462) );
  XNOR2_X1 U522 ( .A(n463), .B(n462), .ZN(n465) );
  XNOR2_X1 U523 ( .A(KEYINPUT109), .B(n587), .ZN(n568) );
  NOR2_X1 U524 ( .A1(n568), .A2(n571), .ZN(n464) );
  NAND2_X1 U525 ( .A1(n465), .A2(n464), .ZN(n466) );
  XNOR2_X1 U526 ( .A(KEYINPUT47), .B(n466), .ZN(n467) );
  XNOR2_X1 U527 ( .A(n467), .B(KEYINPUT111), .ZN(n473) );
  INV_X1 U528 ( .A(KEYINPUT45), .ZN(n469) );
  NOR2_X1 U529 ( .A1(n587), .A2(n590), .ZN(n468) );
  XNOR2_X1 U530 ( .A(n469), .B(n468), .ZN(n470) );
  NOR2_X1 U531 ( .A1(n583), .A2(n470), .ZN(n471) );
  NAND2_X1 U532 ( .A1(n471), .A2(n535), .ZN(n472) );
  NAND2_X1 U533 ( .A1(n473), .A2(n472), .ZN(n475) );
  XOR2_X1 U534 ( .A(KEYINPUT112), .B(KEYINPUT48), .Z(n474) );
  XNOR2_X1 U535 ( .A(n475), .B(n474), .ZN(n553) );
  NOR2_X1 U536 ( .A1(n553), .A2(n497), .ZN(n478) );
  XNOR2_X1 U537 ( .A(KEYINPUT121), .B(KEYINPUT54), .ZN(n476) );
  NOR2_X1 U538 ( .A1(n555), .A2(n479), .ZN(n577) );
  NAND2_X1 U539 ( .A1(n577), .A2(n480), .ZN(n482) );
  XOR2_X1 U540 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n481) );
  XNOR2_X1 U541 ( .A(n482), .B(n481), .ZN(n572) );
  INV_X1 U542 ( .A(n484), .ZN(n540) );
  NAND2_X1 U543 ( .A1(n569), .A2(n540), .ZN(n489) );
  XOR2_X1 U544 ( .A(KEYINPUT125), .B(KEYINPUT124), .Z(n486) );
  XNOR2_X1 U545 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U547 ( .A(KEYINPUT34), .B(KEYINPUT98), .Z(n495) );
  NOR2_X1 U548 ( .A1(n571), .A2(n587), .ZN(n490) );
  XOR2_X1 U549 ( .A(KEYINPUT16), .B(n490), .Z(n491) );
  NOR2_X1 U550 ( .A1(n492), .A2(n491), .ZN(n511) );
  AND2_X1 U551 ( .A1(n493), .A2(n511), .ZN(n502) );
  NAND2_X1 U552 ( .A1(n502), .A2(n555), .ZN(n494) );
  XNOR2_X1 U553 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U554 ( .A(G1GAT), .B(n496), .Z(G1324GAT) );
  INV_X1 U555 ( .A(n497), .ZN(n527) );
  NAND2_X1 U556 ( .A1(n527), .A2(n502), .ZN(n498) );
  XNOR2_X1 U557 ( .A(n498), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT99), .B(KEYINPUT35), .Z(n500) );
  NAND2_X1 U559 ( .A1(n502), .A2(n404), .ZN(n499) );
  XNOR2_X1 U560 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U561 ( .A(G15GAT), .B(n501), .Z(G1326GAT) );
  NAND2_X1 U562 ( .A1(n502), .A2(n531), .ZN(n503) );
  XNOR2_X1 U563 ( .A(n503), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U564 ( .A1(n555), .A2(n508), .ZN(n505) );
  XOR2_X1 U565 ( .A(G29GAT), .B(KEYINPUT39), .Z(n504) );
  XNOR2_X1 U566 ( .A(n505), .B(n504), .ZN(G1328GAT) );
  XNOR2_X1 U567 ( .A(G36GAT), .B(KEYINPUT102), .ZN(n507) );
  NAND2_X1 U568 ( .A1(n508), .A2(n527), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n507), .B(n506), .ZN(G1329GAT) );
  NAND2_X1 U570 ( .A1(n508), .A2(n531), .ZN(n509) );
  XNOR2_X1 U571 ( .A(n509), .B(KEYINPUT104), .ZN(n510) );
  XNOR2_X1 U572 ( .A(G50GAT), .B(n510), .ZN(G1331GAT) );
  NAND2_X1 U573 ( .A1(n540), .A2(n578), .ZN(n524) );
  INV_X1 U574 ( .A(n511), .ZN(n512) );
  NOR2_X1 U575 ( .A1(n524), .A2(n512), .ZN(n518) );
  NAND2_X1 U576 ( .A1(n555), .A2(n518), .ZN(n513) );
  XNOR2_X1 U577 ( .A(KEYINPUT42), .B(n513), .ZN(n514) );
  XNOR2_X1 U578 ( .A(G57GAT), .B(n514), .ZN(G1332GAT) );
  NAND2_X1 U579 ( .A1(n527), .A2(n518), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n515), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U581 ( .A(G71GAT), .B(KEYINPUT105), .Z(n517) );
  NAND2_X1 U582 ( .A1(n518), .A2(n404), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n517), .B(n516), .ZN(G1334GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n520) );
  NAND2_X1 U585 ( .A1(n518), .A2(n531), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n520), .B(n519), .ZN(n522) );
  XOR2_X1 U587 ( .A(G78GAT), .B(KEYINPUT107), .Z(n521) );
  XNOR2_X1 U588 ( .A(n522), .B(n521), .ZN(G1335GAT) );
  INV_X1 U589 ( .A(n523), .ZN(n525) );
  NOR2_X1 U590 ( .A1(n525), .A2(n524), .ZN(n532) );
  NAND2_X1 U591 ( .A1(n555), .A2(n532), .ZN(n526) );
  XNOR2_X1 U592 ( .A(G85GAT), .B(n526), .ZN(G1336GAT) );
  NAND2_X1 U593 ( .A1(n527), .A2(n532), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n528), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U595 ( .A1(n532), .A2(n404), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n529), .B(KEYINPUT108), .ZN(n530) );
  XNOR2_X1 U597 ( .A(G99GAT), .B(n530), .ZN(G1338GAT) );
  NAND2_X1 U598 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n533), .B(KEYINPUT44), .ZN(n534) );
  XNOR2_X1 U600 ( .A(G106GAT), .B(n534), .ZN(G1339GAT) );
  INV_X1 U601 ( .A(n535), .ZN(n566) );
  NOR2_X1 U602 ( .A1(n553), .A2(n536), .ZN(n537) );
  NAND2_X1 U603 ( .A1(n537), .A2(n404), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n538), .B(KEYINPUT113), .ZN(n548) );
  NAND2_X1 U605 ( .A1(n566), .A2(n548), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n539), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n542) );
  NAND2_X1 U608 ( .A1(n548), .A2(n540), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(n544) );
  XOR2_X1 U610 ( .A(G120GAT), .B(KEYINPUT114), .Z(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(G1341GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n546) );
  NAND2_X1 U613 ( .A1(n548), .A2(n568), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U615 ( .A(G127GAT), .B(n547), .Z(G1342GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U617 ( .A1(n548), .A2(n571), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U619 ( .A(G134GAT), .B(n551), .Z(G1343GAT) );
  NOR2_X1 U620 ( .A1(n553), .A2(n552), .ZN(n554) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n563) );
  NOR2_X1 U622 ( .A1(n578), .A2(n563), .ZN(n557) );
  XNOR2_X1 U623 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U625 ( .A(G141GAT), .B(n558), .ZN(G1344GAT) );
  NOR2_X1 U626 ( .A1(n484), .A2(n563), .ZN(n560) );
  XNOR2_X1 U627 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n559) );
  XNOR2_X1 U628 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U629 ( .A(G148GAT), .B(n561), .ZN(G1345GAT) );
  NOR2_X1 U630 ( .A1(n587), .A2(n563), .ZN(n562) );
  XOR2_X1 U631 ( .A(G155GAT), .B(n562), .Z(G1346GAT) );
  NOR2_X1 U632 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U633 ( .A(G162GAT), .B(n565), .Z(G1347GAT) );
  NAND2_X1 U634 ( .A1(n566), .A2(n569), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n567), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n570), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n574) );
  OR2_X1 U639 ( .A1(n572), .A2(n292), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XOR2_X1 U641 ( .A(G190GAT), .B(n575), .Z(G1351GAT) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n589) );
  NOR2_X1 U643 ( .A1(n589), .A2(n578), .ZN(n582) );
  XOR2_X1 U644 ( .A(KEYINPUT59), .B(KEYINPUT127), .Z(n580) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1352GAT) );
  XOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT61), .Z(n586) );
  INV_X1 U649 ( .A(n589), .ZN(n584) );
  NAND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1353GAT) );
  NOR2_X1 U652 ( .A1(n587), .A2(n589), .ZN(n588) );
  XOR2_X1 U653 ( .A(G211GAT), .B(n588), .Z(G1354GAT) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U655 ( .A(KEYINPUT62), .B(n591), .Z(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

