//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 0 0 0 1 0 0 1 0 0 1 0 1 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0 1 0 1 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1232, new_n1233, new_n1234, new_n1235, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n201), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n206), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n209), .B1(new_n213), .B2(new_n215), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n202), .A2(G68), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n217), .A2(G50), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n238), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(G33), .ZN(new_n245));
  INV_X1    g0045(.A(G41), .ZN(new_n246));
  OAI211_X1 g0046(.A(G1), .B(G13), .C1(new_n245), .C2(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G1), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n248), .B1(G41), .B2(G45), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n250), .A2(new_n218), .ZN(new_n251));
  INV_X1    g0051(.A(G45), .ZN(new_n252));
  AOI21_X1  g0052(.A(G1), .B1(new_n246), .B2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT64), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n253), .A2(new_n254), .A3(G274), .ZN(new_n255));
  OAI211_X1 g0055(.A(new_n248), .B(G274), .C1(G41), .C2(G45), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT64), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT72), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n255), .A2(KEYINPUT72), .A3(new_n257), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n251), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AND2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  OAI211_X1 g0064(.A(G232), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  OAI211_X1 g0066(.A(G226), .B(new_n266), .C1(new_n263), .C2(new_n264), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G97), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT71), .ZN(new_n270));
  AND2_X1   g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(new_n210), .ZN(new_n272));
  AND3_X1   g0072(.A1(new_n269), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n270), .B1(new_n269), .B2(new_n272), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n262), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT13), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT13), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n262), .B(new_n277), .C1(new_n273), .C2(new_n274), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n276), .A2(KEYINPUT73), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT73), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n275), .A2(new_n280), .A3(KEYINPUT13), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(G200), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n210), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT66), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT66), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n283), .A2(new_n286), .A3(new_n210), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n285), .A2(new_n287), .B1(new_n248), .B2(G20), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G68), .ZN(new_n289));
  XOR2_X1   g0089(.A(new_n289), .B(KEYINPUT75), .Z(new_n290));
  INV_X1    g0090(.A(G13), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n291), .A2(new_n211), .A3(G1), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(KEYINPUT76), .A3(new_n217), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT12), .ZN(new_n294));
  AOI21_X1  g0094(.A(KEYINPUT76), .B1(new_n292), .B2(new_n217), .ZN(new_n295));
  XOR2_X1   g0095(.A(new_n294), .B(new_n295), .Z(new_n296));
  INV_X1    g0096(.A(new_n287), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n286), .B1(new_n283), .B2(new_n210), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(G20), .A2(G33), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n300), .A2(G50), .B1(G20), .B2(new_n217), .ZN(new_n301));
  INV_X1    g0101(.A(G77), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n211), .A2(G33), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n299), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g0105(.A(KEYINPUT74), .B(KEYINPUT11), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n305), .B(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n290), .A2(new_n296), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n276), .A2(G190), .A3(new_n278), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n282), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n276), .A2(G179), .A3(new_n278), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G169), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n314), .A2(KEYINPUT77), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n279), .A2(new_n281), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT14), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n279), .A2(KEYINPUT14), .A3(new_n281), .A4(new_n315), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n313), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n311), .B1(new_n320), .B2(new_n309), .ZN(new_n321));
  INV_X1    g0121(.A(G58), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n322), .A2(new_n217), .ZN(new_n323));
  OAI21_X1  g0123(.A(G20), .B1(new_n323), .B2(new_n201), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n300), .A2(G159), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT7), .ZN(new_n328));
  NOR4_X1   g0128(.A1(new_n263), .A2(new_n264), .A3(new_n328), .A4(G20), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT78), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(new_n263), .B2(new_n264), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT3), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n245), .ZN(new_n333));
  NAND2_X1  g0133(.A1(KEYINPUT3), .A2(G33), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n333), .A2(KEYINPUT78), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n331), .A2(new_n335), .A3(new_n211), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n329), .B1(new_n336), .B2(new_n328), .ZN(new_n337));
  OAI211_X1 g0137(.A(KEYINPUT16), .B(new_n327), .C1(new_n337), .C2(new_n217), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT16), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n333), .A2(new_n334), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n328), .B1(new_n340), .B2(G20), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n263), .A2(new_n264), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n217), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n339), .B1(new_n344), .B2(new_n326), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n338), .A2(new_n299), .A3(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT79), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n338), .A2(KEYINPUT79), .A3(new_n299), .A4(new_n345), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n285), .A2(new_n287), .ZN(new_n351));
  INV_X1    g0151(.A(new_n292), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT8), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(new_n322), .B2(KEYINPUT67), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT67), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n356), .A2(KEYINPUT8), .A3(G58), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(G1), .B2(new_n211), .ZN(new_n360));
  OAI22_X1  g0160(.A1(new_n353), .A2(new_n360), .B1(new_n352), .B2(new_n359), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n350), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT18), .ZN(new_n364));
  INV_X1    g0164(.A(G232), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n258), .B1(new_n365), .B2(new_n250), .ZN(new_n366));
  INV_X1    g0166(.A(G226), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(G1698), .ZN(new_n368));
  OAI221_X1 g0168(.A(new_n368), .B1(G223), .B2(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n369));
  NAND2_X1  g0169(.A1(G33), .A2(G87), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n247), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OR2_X1    g0171(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n314), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT80), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n366), .A2(new_n371), .ZN(new_n375));
  INV_X1    g0175(.A(G179), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n375), .A2(new_n374), .A3(new_n376), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n363), .A2(new_n364), .A3(new_n380), .ZN(new_n381));
  NOR3_X1   g0181(.A1(new_n366), .A2(G190), .A3(new_n371), .ZN(new_n382));
  INV_X1    g0182(.A(G200), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n382), .B1(new_n383), .B2(new_n372), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n350), .A2(new_n362), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT17), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n361), .B1(new_n348), .B2(new_n349), .ZN(new_n389));
  INV_X1    g0189(.A(new_n379), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(new_n377), .B2(new_n373), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT18), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n389), .A2(KEYINPUT17), .A3(new_n385), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n381), .A2(new_n388), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n250), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n395), .A2(G226), .B1(new_n255), .B2(new_n257), .ZN(new_n396));
  OAI211_X1 g0196(.A(G222), .B(new_n266), .C1(new_n263), .C2(new_n264), .ZN(new_n397));
  OAI211_X1 g0197(.A(G223), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n397), .B(new_n398), .C1(new_n302), .C2(new_n340), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n272), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n396), .A2(new_n400), .A3(KEYINPUT65), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT65), .B1(new_n396), .B2(new_n400), .ZN(new_n402));
  OAI21_X1  g0202(.A(G190), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n203), .A2(G20), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n300), .A2(G150), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n404), .B(new_n405), .C1(new_n358), .C2(new_n303), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n299), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT68), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n352), .A2(G50), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n410), .B1(new_n288), .B2(G50), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n406), .A2(KEYINPUT68), .A3(new_n299), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n409), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT9), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n409), .A2(new_n411), .A3(KEYINPUT9), .A4(new_n412), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n403), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NOR3_X1   g0218(.A1(new_n401), .A2(new_n402), .A3(new_n383), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT10), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT69), .ZN(new_n421));
  AND2_X1   g0221(.A1(KEYINPUT69), .A2(KEYINPUT70), .ZN(new_n422));
  OAI22_X1  g0222(.A1(new_n419), .A2(new_n421), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n418), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n419), .B1(new_n417), .B2(KEYINPUT70), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n424), .B1(new_n425), .B2(new_n420), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n401), .A2(new_n402), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n314), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n428), .B(new_n413), .C1(G179), .C2(new_n427), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G20), .A2(G77), .ZN(new_n431));
  XNOR2_X1  g0231(.A(KEYINPUT15), .B(G87), .ZN(new_n432));
  INV_X1    g0232(.A(new_n300), .ZN(new_n433));
  XNOR2_X1  g0233(.A(KEYINPUT8), .B(G58), .ZN(new_n434));
  OAI221_X1 g0234(.A(new_n431), .B1(new_n432), .B2(new_n303), .C1(new_n433), .C2(new_n434), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n435), .A2(new_n299), .B1(new_n302), .B2(new_n292), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n288), .A2(G77), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(G244), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n258), .B1(new_n439), .B2(new_n250), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n340), .A2(G232), .A3(new_n266), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n340), .A2(G238), .A3(G1698), .ZN(new_n442));
  INV_X1    g0242(.A(G107), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n441), .B(new_n442), .C1(new_n443), .C2(new_n340), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n440), .B1(new_n272), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n438), .B1(new_n445), .B2(G190), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(new_n383), .B2(new_n445), .ZN(new_n447));
  OR2_X1    g0247(.A1(new_n445), .A2(G169), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n445), .A2(new_n376), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(new_n438), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  NOR4_X1   g0251(.A1(new_n321), .A2(new_n394), .A3(new_n430), .A4(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G33), .A2(G283), .ZN(new_n454));
  INV_X1    g0254(.A(G97), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n454), .B(new_n211), .C1(G33), .C2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(G116), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G20), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n456), .A2(new_n284), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT20), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n456), .A2(new_n284), .A3(KEYINPUT20), .A4(new_n458), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n248), .A2(G33), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n351), .A2(G116), .A3(new_n352), .A4(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n291), .A2(G1), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(G20), .A3(new_n457), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n463), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n248), .A2(G45), .ZN(new_n469));
  OR2_X1    g0269(.A1(KEYINPUT5), .A2(G41), .ZN(new_n470));
  NAND2_X1  g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n472), .A2(KEYINPUT81), .A3(G274), .A4(new_n247), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT81), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n252), .A2(G1), .ZN(new_n475));
  INV_X1    g0275(.A(new_n471), .ZN(new_n476));
  NOR2_X1   g0276(.A1(KEYINPUT5), .A2(G41), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(G274), .B1(new_n271), .B2(new_n210), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n474), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n473), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(G264), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n482));
  OAI211_X1 g0282(.A(G257), .B(new_n266), .C1(new_n263), .C2(new_n264), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n333), .A2(G303), .A3(new_n334), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n272), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n472), .A2(new_n272), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G270), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n481), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n468), .A2(new_n489), .A3(G169), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT21), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n489), .A2(G200), .ZN(new_n493));
  INV_X1    g0293(.A(new_n468), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n481), .A2(new_n486), .A3(new_n488), .A4(G190), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n481), .A2(new_n486), .A3(new_n488), .A4(G179), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n468), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n468), .A2(new_n489), .A3(KEYINPUT21), .A4(G169), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n492), .A2(new_n496), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n211), .B(G87), .C1(new_n263), .C2(new_n264), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT22), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT22), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n340), .A2(new_n504), .A3(new_n211), .A4(G87), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT24), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G116), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n508), .A2(G20), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT23), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(new_n211), .B2(G107), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n443), .A2(KEYINPUT23), .A3(G20), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n509), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AND3_X1   g0313(.A1(new_n506), .A2(new_n507), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n507), .B1(new_n506), .B2(new_n513), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n299), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n351), .A2(new_n352), .A3(new_n464), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n517), .A2(new_n443), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n292), .A2(new_n443), .ZN(new_n519));
  XNOR2_X1  g0319(.A(new_n519), .B(KEYINPUT25), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(G250), .B(new_n266), .C1(new_n263), .C2(new_n264), .ZN(new_n522));
  OAI211_X1 g0322(.A(G257), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G294), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n272), .ZN(new_n526));
  AND2_X1   g0326(.A1(new_n481), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n478), .A2(G264), .A3(new_n247), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT82), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n478), .A2(KEYINPUT82), .A3(new_n247), .A4(G264), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(G200), .B1(new_n527), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n481), .A2(new_n526), .A3(new_n528), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n534), .A2(G190), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n516), .B(new_n521), .C1(new_n533), .C2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(G169), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n532), .A2(G179), .A3(new_n481), .A4(new_n526), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n515), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n506), .A2(new_n507), .A3(new_n513), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n351), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n521), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n539), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n536), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n475), .A2(G274), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n469), .A2(G250), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n546), .B1(new_n272), .B2(new_n547), .ZN(new_n548));
  OAI211_X1 g0348(.A(G238), .B(new_n266), .C1(new_n263), .C2(new_n264), .ZN(new_n549));
  OAI211_X1 g0349(.A(G244), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n549), .A2(new_n550), .A3(new_n508), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n548), .B1(new_n551), .B2(new_n272), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n552), .A2(new_n383), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n351), .A2(G87), .A3(new_n352), .A4(new_n464), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT19), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n211), .B1(new_n268), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(G97), .A2(G107), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n219), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n211), .B(G68), .C1(new_n263), .C2(new_n264), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n555), .B1(new_n303), .B2(new_n455), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n299), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n432), .A2(new_n292), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n554), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n553), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n552), .A2(G190), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n551), .A2(new_n272), .ZN(new_n568));
  INV_X1    g0368(.A(new_n548), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n568), .A2(G179), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(new_n314), .B2(new_n552), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n563), .B(new_n564), .C1(new_n517), .C2(new_n432), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n566), .A2(new_n567), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(KEYINPUT7), .B1(new_n342), .B2(new_n211), .ZN(new_n574));
  OAI21_X1  g0374(.A(G107), .B1(new_n574), .B2(new_n329), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT6), .ZN(new_n576));
  AND2_X1   g0376(.A1(G97), .A2(G107), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n576), .B1(new_n577), .B2(new_n557), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n443), .A2(KEYINPUT6), .A3(G97), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n580), .A2(G20), .B1(G77), .B2(new_n300), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n351), .B1(new_n575), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n517), .A2(new_n455), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n352), .A2(G97), .ZN(new_n584));
  NOR3_X1   g0384(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(G244), .B(new_n266), .C1(new_n263), .C2(new_n264), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT4), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n340), .A2(KEYINPUT4), .A3(G244), .A4(new_n266), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n340), .A2(G250), .A3(G1698), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n454), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n272), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n473), .A2(new_n480), .B1(new_n487), .B2(G257), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G200), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n592), .A2(new_n593), .A3(G190), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n585), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n594), .A2(new_n314), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n580), .A2(G20), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n300), .A2(G77), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n443), .B1(new_n341), .B2(new_n343), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n299), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n517), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(G97), .ZN(new_n605));
  INV_X1    g0405(.A(new_n584), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n603), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n592), .A2(new_n593), .A3(new_n376), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n598), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n573), .A2(new_n597), .A3(new_n609), .ZN(new_n610));
  NOR4_X1   g0410(.A1(new_n453), .A2(new_n501), .A3(new_n545), .A4(new_n610), .ZN(G372));
  AOI21_X1  g0411(.A(new_n364), .B1(new_n363), .B2(new_n380), .ZN(new_n612));
  NOR3_X1   g0412(.A1(new_n389), .A2(KEYINPUT18), .A3(new_n391), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n311), .A2(new_n438), .A3(new_n449), .A4(new_n448), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n616), .B1(new_n320), .B2(new_n309), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n389), .A2(KEYINPUT17), .A3(new_n385), .ZN(new_n618));
  AOI21_X1  g0418(.A(KEYINPUT17), .B1(new_n389), .B2(new_n385), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n615), .B1(new_n617), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT85), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n426), .B1(new_n621), .B2(new_n622), .ZN(new_n625));
  OR2_X1    g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n572), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n571), .A2(KEYINPUT83), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT83), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n570), .B(new_n629), .C1(new_n314), .C2(new_n552), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n627), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n566), .A2(new_n567), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n631), .A2(new_n609), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT84), .B1(new_n633), .B2(KEYINPUT26), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n628), .A2(new_n630), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n572), .ZN(new_n636));
  INV_X1    g0436(.A(new_n609), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n566), .A2(new_n567), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT84), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT26), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n637), .A2(KEYINPUT26), .A3(new_n573), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n634), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n536), .A2(new_n609), .A3(new_n597), .A4(new_n638), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n492), .A2(new_n499), .A3(new_n500), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n516), .A2(new_n521), .B1(new_n537), .B2(new_n538), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n649), .A2(new_n631), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n644), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n452), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n626), .A2(new_n429), .A3(new_n652), .ZN(G369));
  NAND2_X1  g0453(.A1(new_n466), .A2(new_n211), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(new_n656), .A3(G213), .ZN(new_n657));
  INV_X1    g0457(.A(G343), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n646), .A2(new_n468), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n659), .ZN(new_n661));
  OAI22_X1  g0461(.A1(new_n501), .A2(KEYINPUT86), .B1(new_n494), .B2(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n501), .A2(KEYINPUT86), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n660), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(G330), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n527), .A2(new_n532), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n383), .ZN(new_n668));
  INV_X1    g0468(.A(new_n535), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n542), .A2(new_n543), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n647), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n671), .B2(new_n661), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n544), .B2(new_n661), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n666), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n646), .A2(new_n661), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  AOI22_X1  g0477(.A1(new_n677), .A2(new_n672), .B1(new_n647), .B2(new_n661), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n675), .A2(new_n678), .ZN(G399));
  INV_X1    g0479(.A(new_n207), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(G41), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n558), .A2(G116), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G1), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n215), .B2(new_n682), .ZN(new_n685));
  XOR2_X1   g0485(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n686));
  XNOR2_X1  g0486(.A(new_n685), .B(new_n686), .ZN(new_n687));
  AOI211_X1 g0487(.A(KEYINPUT29), .B(new_n659), .C1(new_n644), .C2(new_n650), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n637), .A2(new_n641), .A3(new_n573), .ZN(new_n689));
  OAI211_X1 g0489(.A(new_n636), .B(new_n689), .C1(new_n645), .C2(new_n648), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n633), .A2(new_n641), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n661), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n692), .A2(KEYINPUT29), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n688), .A2(new_n693), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n573), .A2(new_n597), .A3(new_n609), .ZN(new_n695));
  INV_X1    g0495(.A(new_n501), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n695), .A2(new_n672), .A3(new_n696), .A4(new_n661), .ZN(new_n697));
  AND3_X1   g0497(.A1(new_n594), .A2(new_n376), .A3(new_n489), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n552), .A2(KEYINPUT88), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n552), .A2(KEYINPUT88), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n698), .A2(new_n667), .A3(new_n699), .A4(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT30), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n532), .A2(new_n526), .A3(new_n552), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n703), .A2(new_n497), .ZN(new_n704));
  OAI211_X1 g0504(.A(KEYINPUT89), .B(new_n702), .C1(new_n704), .C2(new_n594), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT89), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n594), .A2(new_n703), .A3(new_n497), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n706), .B1(new_n707), .B2(KEYINPUT30), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n707), .A2(KEYINPUT30), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n701), .B(new_n705), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  AOI22_X1  g0510(.A1(new_n697), .A2(KEYINPUT31), .B1(new_n659), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n659), .A2(KEYINPUT31), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n707), .B(new_n702), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n712), .B1(new_n713), .B2(new_n701), .ZN(new_n714));
  OAI21_X1  g0514(.A(G330), .B1(new_n711), .B2(new_n714), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n694), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n687), .B1(new_n716), .B2(G1), .ZN(G364));
  NOR2_X1   g0517(.A1(new_n291), .A2(G20), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n248), .B1(new_n718), .B2(G45), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n681), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n666), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n722), .B1(G330), .B2(new_n664), .ZN(new_n723));
  INV_X1    g0523(.A(new_n721), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n210), .B1(G20), .B2(new_n314), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n211), .A2(G190), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OR3_X1    g0528(.A1(KEYINPUT92), .A2(G179), .A3(G200), .ZN(new_n729));
  OAI21_X1  g0529(.A(KEYINPUT92), .B1(G179), .B2(G200), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G159), .ZN(new_n732));
  XOR2_X1   g0532(.A(new_n732), .B(KEYINPUT32), .Z(new_n733));
  INV_X1    g0533(.A(G190), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n211), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n376), .A2(new_n383), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n383), .A2(G179), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n727), .A2(new_n738), .ZN(new_n739));
  OAI22_X1  g0539(.A1(new_n737), .A2(new_n202), .B1(new_n739), .B2(new_n443), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n735), .A2(new_n738), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n376), .A2(G200), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n727), .A2(new_n742), .ZN(new_n743));
  OAI22_X1  g0543(.A1(new_n741), .A2(new_n219), .B1(new_n743), .B2(new_n302), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n736), .A2(new_n727), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n340), .B1(new_n745), .B2(new_n217), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n740), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n734), .B1(new_n729), .B2(new_n730), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n211), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n455), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n735), .A2(new_n742), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT91), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n752), .A2(new_n753), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G58), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n733), .A2(new_n747), .A3(new_n751), .A4(new_n759), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n758), .A2(G322), .B1(G329), .B2(new_n731), .ZN(new_n761));
  INV_X1    g0561(.A(new_n749), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G294), .ZN(new_n763));
  XOR2_X1   g0563(.A(KEYINPUT33), .B(G317), .Z(new_n764));
  INV_X1    g0564(.A(G303), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n764), .A2(new_n745), .B1(new_n741), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G326), .ZN(new_n767));
  INV_X1    g0567(.A(G311), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n737), .A2(new_n767), .B1(new_n743), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n739), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n340), .B1(new_n771), .B2(G283), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n761), .A2(new_n763), .A3(new_n770), .A4(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n726), .B1(new_n760), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n680), .A2(new_n342), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n775), .A2(G355), .B1(new_n457), .B2(new_n680), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n331), .A2(new_n335), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n680), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(G45), .B2(new_n215), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n243), .A2(new_n252), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n776), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OR2_X1    g0581(.A1(new_n781), .A2(KEYINPUT90), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G13), .A2(G33), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(G20), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n785), .B(new_n725), .C1(new_n781), .C2(KEYINPUT90), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n724), .B(new_n774), .C1(new_n782), .C2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n785), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n787), .B1(new_n664), .B2(new_n788), .ZN(new_n789));
  AND2_X1   g0589(.A1(new_n723), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(G396));
  AOI21_X1  g0591(.A(new_n659), .B1(new_n644), .B2(new_n650), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n450), .A2(new_n659), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n438), .A2(new_n659), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n447), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n793), .B1(new_n795), .B2(new_n450), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n792), .B(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n721), .B1(new_n797), .B2(new_n715), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(new_n715), .B2(new_n797), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n725), .A2(new_n783), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n724), .B1(new_n302), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n737), .ZN(new_n802));
  INV_X1    g0602(.A(new_n745), .ZN(new_n803));
  AOI22_X1  g0603(.A1(G137), .A2(new_n802), .B1(new_n803), .B2(G150), .ZN(new_n804));
  INV_X1    g0604(.A(G159), .ZN(new_n805));
  INV_X1    g0605(.A(G143), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n804), .B1(new_n805), .B2(new_n743), .C1(new_n757), .C2(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT34), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n739), .A2(new_n217), .ZN(new_n809));
  INV_X1    g0609(.A(new_n741), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n809), .B1(G50), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G132), .ZN(new_n812));
  INV_X1    g0612(.A(new_n731), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n811), .B(new_n777), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G58), .B2(new_n762), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n739), .A2(new_n219), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(new_n731), .B2(G311), .ZN(new_n817));
  XOR2_X1   g0617(.A(new_n817), .B(KEYINPUT93), .Z(new_n818));
  INV_X1    g0618(.A(G294), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n757), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n743), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G107), .A2(new_n810), .B1(new_n821), .B2(G116), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n765), .B2(new_n737), .ZN(new_n823));
  INV_X1    g0623(.A(G283), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n342), .B1(new_n745), .B2(new_n824), .ZN(new_n825));
  NOR4_X1   g0625(.A1(new_n820), .A2(new_n823), .A3(new_n750), .A4(new_n825), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n808), .A2(new_n815), .B1(new_n818), .B2(new_n826), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n801), .B1(new_n726), .B2(new_n827), .C1(new_n796), .C2(new_n784), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n799), .A2(new_n828), .ZN(G384));
  AOI211_X1 g0629(.A(new_n457), .B(new_n213), .C1(new_n580), .C2(KEYINPUT35), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(KEYINPUT35), .B2(new_n580), .ZN(new_n831));
  XOR2_X1   g0631(.A(new_n831), .B(KEYINPUT36), .Z(new_n832));
  OR3_X1    g0632(.A1(new_n215), .A2(new_n302), .A3(new_n323), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n248), .B(G13), .C1(new_n833), .C2(new_n239), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(G330), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n386), .B1(new_n389), .B2(new_n391), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n657), .B1(new_n350), .B2(new_n362), .ZN(new_n838));
  OAI21_X1  g0638(.A(KEYINPUT37), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n363), .A2(new_n380), .ZN(new_n840));
  INV_X1    g0640(.A(new_n657), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n363), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT37), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n840), .A2(new_n842), .A3(new_n843), .A4(new_n386), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n839), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n394), .A2(new_n838), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g0647(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n327), .B1(new_n337), .B2(new_n217), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n849), .A2(new_n339), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n338), .A2(new_n299), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n841), .B1(new_n852), .B2(new_n361), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n380), .A2(new_n841), .B1(new_n852), .B2(new_n361), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n386), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(KEYINPUT37), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n394), .A2(new_n854), .B1(new_n844), .B2(new_n857), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n847), .A2(new_n848), .B1(new_n858), .B2(KEYINPUT38), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n308), .A2(new_n659), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n311), .B(new_n860), .C1(new_n320), .C2(new_n309), .ZN(new_n861));
  OR2_X1    g0661(.A1(new_n320), .A2(new_n860), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n796), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n697), .A2(KEYINPUT31), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n710), .A2(new_n659), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n710), .A2(KEYINPUT31), .A3(new_n659), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n864), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n863), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT40), .B1(new_n859), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT38), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n853), .B1(new_n614), .B2(new_n620), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n843), .B1(new_n855), .B2(new_n386), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n389), .A2(new_n391), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n361), .B(new_n384), .C1(new_n348), .C2(new_n349), .ZN(new_n876));
  NOR3_X1   g0676(.A1(new_n875), .A2(new_n838), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n874), .B1(new_n877), .B2(new_n843), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n872), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n394), .A2(new_n854), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n844), .A2(new_n857), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n880), .A2(KEYINPUT38), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n868), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n796), .B1(new_n711), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(new_n861), .B2(new_n862), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT40), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n883), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n871), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n889), .B(KEYINPUT96), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n867), .A2(new_n868), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n452), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n836), .B1(new_n890), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n893), .B2(new_n890), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n614), .A2(new_n841), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n793), .B(KEYINPUT94), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n792), .B2(new_n796), .ZN(new_n899));
  INV_X1    g0699(.A(new_n863), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n896), .B1(new_n901), .B2(new_n883), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n844), .A2(new_n839), .B1(new_n394), .B2(new_n838), .ZN(new_n903));
  INV_X1    g0703(.A(new_n848), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n882), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT39), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n320), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(new_n308), .A3(new_n661), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n879), .A2(KEYINPUT39), .A3(new_n882), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n907), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n902), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n452), .B1(new_n688), .B2(new_n693), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n914), .B(new_n429), .C1(new_n624), .C2(new_n625), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n913), .B(new_n915), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n895), .A2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT97), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI221_X1 g0719(.A(new_n919), .B1(new_n248), .B2(new_n718), .C1(new_n916), .C2(new_n895), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n917), .A2(new_n918), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n835), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n922), .B(KEYINPUT98), .Z(G367));
  NOR2_X1   g0723(.A1(new_n785), .A2(new_n725), .ZN(new_n924));
  INV_X1    g0724(.A(new_n778), .ZN(new_n925));
  OAI221_X1 g0725(.A(new_n924), .B1(new_n207), .B2(new_n432), .C1(new_n925), .C2(new_n234), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT100), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n927), .A2(new_n724), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n737), .A2(new_n768), .B1(new_n745), .B2(new_n819), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n771), .A2(G97), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n824), .B2(new_n743), .ZN(new_n931));
  AOI211_X1 g0731(.A(new_n929), .B(new_n931), .C1(G317), .C2(new_n731), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n758), .A2(G303), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n762), .A2(G107), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n810), .A2(G116), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT46), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n331), .B(new_n335), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n936), .B2(new_n935), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n932), .A2(new_n933), .A3(new_n934), .A4(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n739), .A2(new_n302), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(G50), .B2(new_n821), .ZN(new_n941));
  OAI221_X1 g0741(.A(new_n941), .B1(new_n322), .B2(new_n741), .C1(new_n806), .C2(new_n737), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n340), .B1(new_n745), .B2(new_n805), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(G150), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n757), .A2(new_n945), .B1(new_n217), .B2(new_n749), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT101), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(G137), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n944), .B(new_n948), .C1(new_n949), .C2(new_n813), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n946), .A2(new_n947), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n939), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT47), .Z(new_n953));
  OAI21_X1  g0753(.A(new_n928), .B1(new_n953), .B2(new_n726), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n565), .A2(new_n659), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n636), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n631), .A2(new_n632), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n956), .B1(new_n957), .B2(new_n955), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n954), .B1(new_n785), .B2(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT102), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n597), .B(new_n609), .C1(new_n585), .C2(new_n661), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n637), .A2(new_n659), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n678), .A2(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT45), .Z(new_n965));
  NOR2_X1   g0765(.A1(new_n678), .A2(new_n963), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT44), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n675), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n968), .B(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n677), .A2(new_n672), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n674), .B2(new_n677), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(new_n666), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n716), .A2(new_n973), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n970), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n716), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n681), .B(KEYINPUT41), .Z(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n720), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n963), .A2(new_n672), .A3(new_n677), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT42), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n609), .B1(new_n961), .B2(new_n544), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n982), .A2(new_n661), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT43), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n981), .A2(new_n983), .B1(new_n984), .B2(new_n958), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n958), .A2(new_n984), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n985), .B(new_n986), .Z(new_n987));
  NAND3_X1  g0787(.A1(new_n969), .A2(KEYINPUT99), .A3(new_n963), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(KEYINPUT99), .B1(new_n969), .B2(new_n963), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n989), .B(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n960), .B1(new_n979), .B2(new_n991), .ZN(G387));
  INV_X1    g0792(.A(new_n683), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n993), .A2(new_n775), .B1(new_n443), .B2(new_n680), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n231), .A2(new_n252), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n434), .A2(G50), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT50), .Z(new_n997));
  OAI211_X1 g0797(.A(new_n683), .B(new_n252), .C1(new_n217), .C2(new_n302), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n778), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n994), .B1(new_n995), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n724), .B1(new_n1000), .B2(new_n924), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n674), .B2(new_n788), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n777), .B1(new_n358), .B2(new_n745), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n930), .B1(new_n217), .B2(new_n743), .C1(new_n805), .C2(new_n737), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n1003), .B(new_n1004), .C1(G50), .C2(new_n758), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n749), .A2(new_n432), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(KEYINPUT103), .B(G150), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n813), .A2(new_n1007), .B1(new_n302), .B2(new_n741), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT104), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1005), .A2(new_n1006), .A3(new_n1009), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n762), .A2(G283), .B1(G294), .B2(new_n810), .ZN(new_n1011));
  INV_X1    g0811(.A(G317), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n757), .A2(new_n1012), .B1(new_n765), .B2(new_n743), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1013), .A2(KEYINPUT105), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(KEYINPUT105), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G322), .A2(new_n802), .B1(new_n803), .B2(G311), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT48), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1011), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT106), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1020), .A2(KEYINPUT49), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n777), .B1(G116), .B2(new_n771), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1022), .B(new_n1023), .C1(new_n767), .C2(new_n813), .ZN(new_n1024));
  AOI21_X1  g0824(.A(KEYINPUT49), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1010), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1002), .B1(new_n1026), .B2(new_n725), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n720), .B2(new_n973), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n974), .A2(new_n681), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n716), .A2(new_n973), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1028), .B1(new_n1029), .B2(new_n1030), .ZN(G393));
  NOR2_X1   g0831(.A1(new_n963), .A2(new_n788), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT107), .Z(new_n1033));
  OAI22_X1  g0833(.A1(new_n741), .A2(new_n217), .B1(new_n743), .B2(new_n434), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n816), .B(new_n1034), .C1(G50), .C2(new_n803), .ZN(new_n1035));
  AND2_X1   g0835(.A1(new_n1035), .A2(new_n777), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1036), .B1(new_n302), .B2(new_n749), .C1(new_n806), .C2(new_n813), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n757), .A2(new_n805), .B1(new_n945), .B2(new_n737), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(KEYINPUT108), .B(KEYINPUT51), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1038), .B(new_n1039), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n757), .A2(new_n768), .B1(new_n1012), .B2(new_n737), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT52), .Z(new_n1042));
  NAND2_X1  g0842(.A1(new_n762), .A2(G116), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n731), .A2(G322), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n741), .A2(new_n824), .B1(new_n743), .B2(new_n819), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(G303), .B2(new_n803), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n340), .B1(new_n771), .B2(G107), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1043), .A2(new_n1044), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n1037), .A2(new_n1040), .B1(new_n1042), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n725), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n924), .B1(new_n455), .B2(new_n207), .C1(new_n925), .C2(new_n238), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1033), .A2(new_n721), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n970), .B2(new_n719), .ZN(new_n1053));
  AND2_X1   g0853(.A1(new_n975), .A2(new_n681), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n970), .A2(new_n974), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1053), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(G390));
  NAND3_X1  g0857(.A1(new_n869), .A2(new_n863), .A3(G330), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n659), .B(new_n864), .C1(new_n644), .C2(new_n650), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n863), .B1(new_n1060), .B2(new_n898), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n907), .A2(new_n911), .B1(new_n1061), .B2(new_n909), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n897), .B1(new_n692), .B2(new_n864), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(KEYINPUT109), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT109), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1065), .B(new_n897), .C1(new_n692), .C2(new_n864), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(new_n863), .A3(new_n1066), .ZN(new_n1067));
  AND3_X1   g0867(.A1(new_n1067), .A2(new_n909), .A3(new_n905), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1059), .B1(new_n1062), .B2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n859), .A2(KEYINPUT39), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n911), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n1070), .A2(new_n1071), .B1(new_n901), .B2(new_n910), .ZN(new_n1072));
  OAI211_X1 g0872(.A(G330), .B(new_n796), .C1(new_n711), .C2(new_n714), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n863), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1067), .A2(new_n909), .A3(new_n905), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1072), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1069), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT110), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n1074), .B2(new_n863), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n900), .A2(KEYINPUT110), .A3(new_n1073), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1080), .A2(new_n1081), .A3(new_n1058), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n899), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1084), .A2(new_n1075), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n900), .B1(new_n836), .B2(new_n885), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1082), .A2(new_n1083), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n893), .A2(G330), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n626), .A2(new_n1088), .A3(new_n429), .A4(new_n914), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(KEYINPUT111), .B1(new_n1078), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1069), .A2(new_n1077), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n915), .B1(G330), .B2(new_n893), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1086), .A2(new_n1084), .A3(new_n1075), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT111), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1092), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1077), .A2(new_n1069), .A3(new_n1093), .A4(new_n1096), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1091), .A2(new_n681), .A3(new_n1099), .A4(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n783), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n724), .B1(new_n358), .B2(new_n800), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n340), .B(new_n809), .C1(G87), .C2(new_n810), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n457), .B2(new_n757), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G107), .A2(new_n803), .B1(new_n821), .B2(G97), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n824), .B2(new_n737), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT113), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1107), .A2(new_n1108), .B1(G77), .B2(new_n762), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n1108), .B2(new_n1107), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n1105), .B(new_n1110), .C1(G294), .C2(new_n731), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  AND2_X1   g0912(.A1(new_n1112), .A2(KEYINPUT114), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1112), .A2(KEYINPUT114), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n741), .A2(new_n1007), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT53), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT54), .B(G143), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT112), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n758), .A2(G132), .B1(new_n821), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n762), .A2(G159), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n340), .B1(new_n739), .B2(new_n202), .ZN(new_n1121));
  INV_X1    g0921(.A(G128), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n737), .A2(new_n1122), .B1(new_n745), .B2(new_n949), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n1121), .B(new_n1123), .C1(G125), .C2(new_n731), .ZN(new_n1124));
  AND4_X1   g0924(.A1(new_n1116), .A2(new_n1119), .A3(new_n1120), .A4(new_n1124), .ZN(new_n1125));
  NOR3_X1   g0925(.A1(new_n1113), .A2(new_n1114), .A3(new_n1125), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1102), .B(new_n1103), .C1(new_n726), .C2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n1092), .B2(new_n719), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT115), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  OAI211_X1 g0930(.A(KEYINPUT115), .B(new_n1127), .C1(new_n1092), .C2(new_n719), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1101), .A2(new_n1132), .ZN(G378));
  INV_X1    g0933(.A(KEYINPUT119), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n413), .A2(new_n841), .ZN(new_n1135));
  XOR2_X1   g0935(.A(new_n1135), .B(KEYINPUT55), .Z(new_n1136));
  INV_X1    g0936(.A(KEYINPUT117), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n426), .A2(new_n1137), .A3(new_n429), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1137), .B1(new_n426), .B2(new_n429), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1136), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n430), .A2(KEYINPUT117), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1136), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1142), .A2(new_n1143), .A3(new_n1138), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n1141), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1145), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n880), .A2(KEYINPUT38), .A3(new_n881), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n904), .B1(new_n845), .B2(new_n846), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n863), .B(new_n869), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(KEYINPUT40), .B1(new_n879), .B2(new_n882), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1151), .A2(KEYINPUT40), .B1(new_n1152), .B2(new_n886), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1148), .B1(new_n1153), .B2(new_n836), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n902), .A2(new_n912), .ZN(new_n1155));
  OR2_X1    g0955(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n889), .A2(G330), .A3(new_n1156), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n1154), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1155), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1134), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NOR3_X1   g0960(.A1(new_n1153), .A2(new_n836), .A3(new_n1148), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1156), .B1(new_n889), .B2(G330), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n913), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1154), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1163), .A2(KEYINPUT119), .A3(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1160), .A2(new_n720), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n724), .B1(new_n202), .B2(new_n800), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n777), .A2(G41), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1168), .B1(new_n824), .B2(new_n813), .C1(new_n757), .C2(new_n443), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n749), .A2(new_n217), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n741), .A2(new_n302), .B1(new_n743), .B2(new_n432), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(G116), .A2(new_n802), .B1(new_n803), .B2(G97), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n322), .B2(new_n739), .ZN(new_n1173));
  NOR4_X1   g0973(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .A4(new_n1173), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1174), .B(KEYINPUT58), .Z(new_n1175));
  OAI21_X1  g0975(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n802), .A2(G125), .B1(new_n821), .B2(G137), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n812), .B2(new_n745), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n810), .B2(new_n1118), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n1122), .B2(new_n757), .C1(new_n945), .C2(new_n749), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1180), .A2(KEYINPUT59), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(KEYINPUT59), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n245), .B(new_n246), .C1(new_n739), .C2(new_n805), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(G124), .B2(new_n731), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1175), .B1(new_n1168), .B2(new_n1176), .C1(new_n1181), .C2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1186), .A2(KEYINPUT116), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(KEYINPUT116), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n725), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1167), .B1(new_n1187), .B2(new_n1189), .C1(new_n1156), .C2(new_n784), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1166), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT57), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n1100), .B2(new_n1093), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT120), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1196));
  AND2_X1   g0996(.A1(new_n1164), .A2(new_n1195), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1194), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1198), .A2(KEYINPUT121), .A3(new_n681), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1100), .A2(new_n1093), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1160), .A2(new_n1200), .A3(new_n1165), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n1193), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1199), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(KEYINPUT121), .B1(new_n1198), .B2(new_n681), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1192), .B1(new_n1203), .B2(new_n1204), .ZN(G375));
  OAI21_X1  g1005(.A(KEYINPUT122), .B1(new_n1087), .B2(new_n719), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT122), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1096), .A2(new_n1207), .A3(new_n720), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(G116), .A2(new_n803), .B1(new_n821), .B2(G107), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n819), .B2(new_n737), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT123), .ZN(new_n1211));
  OR2_X1    g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1212), .A2(new_n1006), .A3(new_n1213), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n340), .B(new_n940), .C1(G97), .C2(new_n810), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1215), .B1(new_n824), .B2(new_n757), .C1(new_n765), .C2(new_n813), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n1118), .A2(new_n803), .B1(G128), .B2(new_n731), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n949), .B2(new_n757), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n762), .A2(G50), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(G159), .A2(new_n810), .B1(new_n771), .B2(G58), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n802), .A2(G132), .B1(new_n821), .B2(G150), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1219), .A2(new_n777), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n1214), .A2(new_n1216), .B1(new_n1218), .B2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n725), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n724), .B1(new_n217), .B2(new_n800), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1224), .B(new_n1225), .C1(new_n863), .C2(new_n784), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1206), .A2(new_n1208), .A3(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1097), .A2(new_n1229), .A3(new_n978), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1228), .A2(new_n1230), .ZN(G381));
  OAI211_X1 g1031(.A(new_n1056), .B(new_n960), .C1(new_n991), .C2(new_n979), .ZN(new_n1232));
  OR4_X1    g1032(.A1(G396), .A2(new_n1232), .A3(G384), .A4(G393), .ZN(new_n1233));
  INV_X1    g1033(.A(G378), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1234), .B(new_n1192), .C1(new_n1203), .C2(new_n1204), .ZN(new_n1235));
  OR3_X1    g1035(.A1(new_n1233), .A2(new_n1235), .A3(G381), .ZN(G407));
  OAI211_X1 g1036(.A(G407), .B(G213), .C1(G343), .C2(new_n1235), .ZN(G409));
  OAI21_X1  g1037(.A(new_n720), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1101), .A2(new_n1132), .A3(new_n1238), .A4(new_n1190), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1201), .A2(new_n977), .ZN(new_n1240));
  INV_X1    g1040(.A(G213), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n1239), .A2(new_n1240), .B1(new_n1241), .B2(G343), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(KEYINPUT120), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1164), .A2(new_n1195), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n682), .B1(new_n1246), .B2(new_n1194), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1247), .A2(KEYINPUT121), .B1(new_n1193), .B2(new_n1201), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1204), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1191), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1243), .B1(new_n1250), .B2(new_n1234), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT124), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1241), .A2(G343), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(G2897), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1087), .A2(new_n1089), .A3(KEYINPUT60), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n681), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1097), .A2(KEYINPUT60), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1257), .B1(new_n1229), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(G384), .ZN(new_n1260));
  NOR3_X1   g1060(.A1(new_n1259), .A2(new_n1260), .A3(new_n1227), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT60), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1229), .B1(new_n1090), .B2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1263), .A2(new_n681), .A3(new_n1256), .ZN(new_n1264));
  AOI21_X1  g1064(.A(G384), .B1(new_n1264), .B2(new_n1228), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1252), .B(new_n1255), .C1(new_n1261), .C2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1252), .B1(new_n1261), .B2(new_n1265), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1260), .B1(new_n1259), .B2(new_n1227), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1264), .A2(G384), .A3(new_n1228), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1269), .A2(new_n1270), .A3(KEYINPUT124), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1255), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1267), .B1(new_n1268), .B2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT61), .B1(new_n1251), .B2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(G375), .A2(G378), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1261), .A2(new_n1265), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1275), .A2(new_n1243), .A3(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT63), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT125), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G387), .A2(G390), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1280), .B1(new_n1281), .B2(new_n1232), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  XNOR2_X1  g1083(.A(G393), .B(new_n790), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1281), .A2(new_n1232), .A3(new_n1280), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1283), .A2(new_n1285), .A3(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1285), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1282), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1242), .B1(G375), .B2(G378), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1292), .A2(KEYINPUT63), .A3(new_n1276), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1274), .A2(new_n1279), .A3(new_n1291), .A4(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT61), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1272), .A2(new_n1268), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1266), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1295), .B1(new_n1292), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT62), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1277), .A2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1292), .A2(KEYINPUT62), .A3(new_n1276), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1298), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT126), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1290), .A2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1287), .A2(KEYINPUT126), .A3(new_n1289), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1294), .B1(new_n1302), .B2(new_n1306), .ZN(G405));
  INV_X1    g1107(.A(KEYINPUT127), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1275), .A2(new_n1235), .A3(new_n1276), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1276), .B1(new_n1275), .B2(new_n1235), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1290), .B(new_n1308), .C1(new_n1310), .C2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1311), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1290), .A2(new_n1308), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1287), .A2(KEYINPUT127), .A3(new_n1289), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1313), .A2(new_n1314), .A3(new_n1309), .A4(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1312), .A2(new_n1316), .ZN(G402));
endmodule


