//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1 0 0 0 1 0 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0 0 1 1 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1305, new_n1306, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380, new_n1381, new_n1382, new_n1383,
    new_n1384, new_n1385, new_n1386, new_n1387, new_n1388;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G77), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT65), .Z(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G250), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G257), .ZN(new_n210));
  INV_X1    g0010(.A(G264), .ZN(new_n211));
  AOI211_X1 g0011(.A(new_n206), .B(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NOR2_X1   g0015(.A1(G58), .A2(G68), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(new_n212), .A2(KEYINPUT0), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n220), .B1(KEYINPUT0), .B2(new_n212), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT66), .Z(new_n222));
  XNOR2_X1  g0022(.A(KEYINPUT68), .B(G244), .ZN(new_n223));
  XNOR2_X1  g0023(.A(KEYINPUT67), .B(G68), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(new_n223), .B1(new_n224), .B2(G238), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n228));
  NAND4_X1  g0028(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(new_n207), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT69), .ZN(new_n231));
  INV_X1    g0031(.A(KEYINPUT1), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AND2_X1   g0033(.A1(new_n231), .A2(new_n232), .ZN(new_n234));
  NOR3_X1   g0034(.A1(new_n222), .A2(new_n233), .A3(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT2), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT70), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G1), .A3(G13), .ZN(new_n254));
  MUX2_X1   g0054(.A(G222), .B(G223), .S(G1698), .Z(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT3), .B(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G77), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n257), .B1(new_n258), .B2(new_n256), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n254), .B1(new_n259), .B2(KEYINPUT71), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n260), .B1(KEYINPUT71), .B2(new_n259), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n254), .A2(G274), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n263), .B1(G41), .B2(G45), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n254), .A2(new_n264), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n265), .B1(G226), .B2(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G190), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n202), .A2(G20), .ZN(new_n270));
  INV_X1    g0070(.A(G150), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G20), .A2(G33), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT8), .B(G58), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT72), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT72), .ZN(new_n276));
  INV_X1    g0076(.A(G58), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(new_n277), .A3(KEYINPUT8), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G33), .ZN(new_n280));
  OAI21_X1  g0080(.A(KEYINPUT73), .B1(new_n280), .B2(G20), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT73), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(new_n214), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  OAI221_X1 g0085(.A(new_n270), .B1(new_n271), .B2(new_n273), .C1(new_n279), .C2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n213), .B1(new_n207), .B2(new_n280), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n263), .A2(G13), .A3(G20), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT74), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n263), .A2(KEYINPUT74), .A3(G13), .A4(G20), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n287), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G50), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n297), .B1(new_n263), .B2(G20), .ZN(new_n298));
  INV_X1    g0098(.A(new_n293), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n296), .A2(new_n298), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n288), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT9), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n288), .A2(KEYINPUT9), .A3(new_n300), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n261), .A2(new_n267), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G200), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n269), .A2(new_n303), .A3(new_n304), .A4(new_n306), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n307), .B(KEYINPUT10), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT3), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G33), .ZN(new_n310));
  INV_X1    g0110(.A(G226), .ZN(new_n311));
  INV_X1    g0111(.A(G1698), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n280), .A2(KEYINPUT3), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n237), .A2(G1698), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n310), .A2(new_n313), .A3(new_n314), .A4(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G33), .A2(G97), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n254), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n264), .ZN(new_n320));
  INV_X1    g0120(.A(G274), .ZN(new_n321));
  AND2_X1   g0121(.A1(G1), .A2(G13), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n321), .B1(new_n322), .B2(new_n253), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n266), .A2(G238), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  AND4_X1   g0124(.A1(KEYINPUT79), .A2(new_n319), .A3(new_n324), .A4(KEYINPUT13), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n319), .A2(new_n324), .B1(KEYINPUT79), .B2(KEYINPUT13), .ZN(new_n326));
  OAI21_X1  g0126(.A(G179), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n319), .A2(new_n324), .A3(KEYINPUT13), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT13), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n323), .A2(new_n320), .ZN(new_n330));
  INV_X1    g0130(.A(G238), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n254), .A2(new_n264), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n329), .B1(new_n333), .B2(new_n318), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n328), .A2(new_n334), .A3(G169), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT14), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT14), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n328), .A2(new_n334), .A3(new_n337), .A4(G169), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n327), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n224), .A2(new_n214), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n258), .B1(new_n281), .B2(new_n283), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT80), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(KEYINPUT80), .B1(new_n340), .B2(new_n341), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n272), .A2(G50), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n287), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT11), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n342), .A2(new_n343), .B1(G50), .B2(new_n272), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n294), .B1(new_n351), .B2(new_n345), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT11), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT76), .ZN(new_n354));
  AND3_X1   g0154(.A1(new_n291), .A2(new_n354), .A3(new_n292), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n354), .B1(new_n291), .B2(new_n292), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AND2_X1   g0157(.A1(KEYINPUT67), .A2(G68), .ZN(new_n358));
  NOR2_X1   g0158(.A1(KEYINPUT67), .A2(G68), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n357), .A2(KEYINPUT12), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G68), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n362), .B1(new_n263), .B2(G20), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n294), .B(new_n363), .C1(new_n355), .C2(new_n356), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT12), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(new_n293), .B2(G68), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n361), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n350), .A2(new_n353), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n339), .A2(new_n369), .ZN(new_n370));
  XOR2_X1   g0170(.A(KEYINPUT8), .B(G58), .Z(new_n371));
  AOI22_X1  g0171(.A1(new_n371), .A2(new_n272), .B1(G20), .B2(G77), .ZN(new_n372));
  XNOR2_X1  g0172(.A(KEYINPUT15), .B(G87), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n284), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n258), .A2(new_n357), .B1(new_n376), .B2(new_n287), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n293), .A2(KEYINPUT76), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n291), .A2(new_n354), .A3(new_n292), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n287), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n258), .B1(new_n263), .B2(G20), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT77), .ZN(new_n384));
  INV_X1    g0184(.A(G200), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n265), .B1(new_n223), .B2(new_n266), .ZN(new_n386));
  NOR2_X1   g0186(.A1(G232), .A2(G1698), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n312), .A2(G238), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n256), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n254), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n389), .B(new_n390), .C1(G107), .C2(new_n256), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n385), .B1(new_n386), .B2(new_n391), .ZN(new_n392));
  OR3_X1    g0192(.A1(new_n383), .A2(new_n384), .A3(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n384), .B1(new_n383), .B2(new_n392), .ZN(new_n394));
  INV_X1    g0194(.A(G190), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n386), .A2(new_n391), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n393), .B(new_n394), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n367), .B1(new_n352), .B2(KEYINPUT11), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n328), .A2(new_n334), .A3(G200), .ZN(new_n399));
  OAI21_X1  g0199(.A(G190), .B1(new_n325), .B2(new_n326), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n398), .A2(new_n350), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n396), .A2(G179), .ZN(new_n402));
  XNOR2_X1  g0202(.A(new_n402), .B(KEYINPUT78), .ZN(new_n403));
  INV_X1    g0203(.A(G169), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n396), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(new_n383), .A3(new_n405), .ZN(new_n406));
  AND4_X1   g0206(.A1(new_n370), .A2(new_n397), .A3(new_n401), .A4(new_n406), .ZN(new_n407));
  OR2_X1    g0207(.A1(G223), .A2(G1698), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n311), .A2(G1698), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n310), .A2(new_n408), .A3(new_n314), .A4(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G33), .A2(G87), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n254), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n266), .A2(G232), .B1(new_n320), .B2(new_n323), .ZN(new_n414));
  INV_X1    g0214(.A(G179), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT83), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n413), .A2(new_n414), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n404), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT83), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n413), .A2(new_n414), .A3(new_n420), .A4(new_n415), .ZN(new_n421));
  AND3_X1   g0221(.A1(new_n417), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  XOR2_X1   g0222(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n423));
  INV_X1    g0223(.A(KEYINPUT82), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(new_n280), .B2(KEYINPUT3), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n309), .A2(KEYINPUT82), .A3(G33), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n425), .A2(new_n314), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT7), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(G20), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n428), .B1(new_n256), .B2(G20), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n360), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n216), .B1(new_n224), .B2(G58), .ZN(new_n433));
  INV_X1    g0233(.A(G159), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n433), .A2(new_n214), .B1(new_n434), .B2(new_n273), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n423), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  NOR3_X1   g0236(.A1(new_n256), .A2(new_n428), .A3(G20), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n310), .A2(new_n314), .ZN(new_n438));
  AOI21_X1  g0238(.A(KEYINPUT7), .B1(new_n438), .B2(new_n214), .ZN(new_n439));
  OAI21_X1  g0239(.A(G68), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n217), .B1(new_n360), .B2(new_n277), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n441), .A2(G20), .B1(G159), .B2(new_n272), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n440), .A2(new_n442), .A3(KEYINPUT16), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n436), .A2(new_n287), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n279), .B1(new_n263), .B2(G20), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n445), .A2(new_n296), .B1(new_n299), .B2(new_n279), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT18), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n422), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n448), .B1(new_n422), .B2(new_n447), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n330), .B1(new_n237), .B2(new_n332), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n385), .B1(new_n452), .B2(new_n412), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n453), .B1(new_n418), .B2(G190), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n444), .A2(new_n446), .A3(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT17), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n444), .A2(KEYINPUT17), .A3(new_n446), .A4(new_n454), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n451), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT75), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n305), .A2(new_n463), .A3(G179), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT75), .B1(new_n268), .B2(new_n415), .ZN(new_n465));
  OAI221_X1 g0265(.A(new_n301), .B1(G169), .B2(new_n268), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n308), .A2(new_n407), .A3(new_n462), .A4(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G116), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n378), .A2(new_n468), .A3(new_n379), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G283), .ZN(new_n470));
  INV_X1    g0270(.A(G97), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n470), .B(new_n214), .C1(G33), .C2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n468), .A2(G20), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(new_n287), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT20), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n472), .A2(new_n287), .A3(KEYINPUT20), .A4(new_n473), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n469), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT87), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n263), .A2(G33), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(new_n468), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n481), .B1(new_n380), .B2(new_n484), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n294), .B(new_n484), .C1(new_n355), .C2(new_n356), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(KEYINPUT87), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n480), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G45), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(G1), .ZN(new_n490));
  AND2_X1   g0290(.A1(KEYINPUT5), .A2(G41), .ZN(new_n491));
  NOR2_X1   g0291(.A1(KEYINPUT5), .A2(G41), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n262), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n493), .A2(new_n254), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n494), .B1(new_n495), .B2(G270), .ZN(new_n496));
  INV_X1    g0296(.A(G303), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n438), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(G257), .A2(G1698), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n499), .B1(new_n211), .B2(G1698), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n498), .B(new_n390), .C1(new_n438), .C2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G169), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n488), .A2(KEYINPUT21), .A3(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT21), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n486), .A2(KEYINPUT87), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n378), .A2(new_n379), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n508), .A2(new_n481), .A3(new_n294), .A4(new_n484), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n479), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n506), .B1(new_n510), .B2(new_n503), .ZN(new_n511));
  OR2_X1    g0311(.A1(new_n262), .A2(new_n493), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n493), .A2(G270), .A3(new_n254), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n501), .A2(G179), .A3(new_n512), .A4(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n488), .A2(new_n515), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n496), .A2(new_n501), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G190), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n502), .A2(G200), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n510), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n505), .A2(new_n511), .A3(new_n516), .A4(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(G244), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n522), .A2(G1698), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n523), .A2(new_n310), .A3(new_n314), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT4), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n256), .A2(KEYINPUT4), .A3(new_n523), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n310), .A2(new_n314), .A3(G250), .A4(G1698), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n526), .A2(new_n527), .A3(new_n470), .A4(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n390), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n495), .A2(G257), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n530), .A2(G190), .A3(new_n512), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT84), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n530), .A2(new_n512), .A3(new_n531), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G200), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n299), .A2(new_n471), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n293), .A2(new_n294), .A3(G97), .A4(new_n482), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT6), .ZN(new_n539));
  AND2_X1   g0339(.A1(G97), .A2(G107), .ZN(new_n540));
  NOR2_X1   g0340(.A1(G97), .A2(G107), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(G107), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n543), .A2(KEYINPUT6), .A3(G97), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n545), .A2(G20), .B1(G77), .B2(new_n272), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n438), .A2(new_n214), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n547), .A2(new_n428), .B1(new_n427), .B2(new_n429), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n546), .B1(new_n548), .B2(new_n543), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n538), .B1(new_n549), .B2(new_n287), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n529), .A2(new_n390), .B1(G257), .B2(new_n495), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT84), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n551), .A2(new_n552), .A3(G190), .A4(new_n512), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n533), .A2(new_n535), .A3(new_n550), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n549), .A2(new_n287), .ZN(new_n555));
  INV_X1    g0355(.A(new_n538), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n534), .A2(new_n404), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n551), .A2(new_n415), .A3(new_n512), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n554), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n310), .A2(new_n314), .A3(new_n214), .A4(G87), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT22), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT22), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n256), .A2(new_n564), .A3(new_n214), .A4(G87), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT24), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n280), .A2(new_n468), .A3(G20), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT23), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n214), .B2(G107), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n543), .A2(KEYINPUT23), .A3(G20), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n568), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n566), .A2(new_n567), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n567), .B1(new_n566), .B2(new_n572), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n287), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n295), .A2(new_n483), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n299), .A2(KEYINPUT25), .A3(new_n543), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT25), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n293), .B2(G107), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n576), .A2(G107), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n493), .A2(G264), .A3(new_n254), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n206), .A2(new_n312), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n210), .A2(G1698), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n310), .A2(new_n583), .A3(new_n314), .A4(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(G294), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n280), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n254), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(KEYINPUT88), .B1(new_n582), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT88), .ZN(new_n591));
  NOR2_X1   g0391(.A1(G250), .A2(G1698), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n592), .B1(new_n210), .B2(G1698), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n587), .B1(new_n593), .B2(new_n256), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n591), .B(new_n581), .C1(new_n594), .C2(new_n254), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n590), .A2(G179), .A3(new_n512), .A4(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n512), .B(new_n581), .C1(new_n254), .C2(new_n594), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(G169), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n575), .A2(new_n580), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n575), .A2(new_n580), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n590), .A2(new_n512), .A3(new_n595), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n385), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(G190), .B2(new_n597), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n599), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n310), .A2(new_n314), .A3(new_n214), .A4(G68), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT19), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n214), .B1(new_n317), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(G87), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n541), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n471), .B1(new_n281), .B2(new_n283), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n606), .B(new_n611), .C1(new_n612), .C2(KEYINPUT19), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n357), .A2(new_n373), .B1(new_n613), .B2(new_n287), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT85), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n331), .A2(new_n312), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n522), .A2(G1698), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n310), .A2(new_n616), .A3(new_n314), .A4(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n280), .A2(new_n468), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n254), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n254), .A2(G274), .A3(new_n490), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n206), .B1(new_n263), .B2(G45), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n254), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(G200), .B1(new_n621), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n293), .A2(new_n294), .A3(G87), .A4(new_n482), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n614), .A2(new_n615), .A3(new_n626), .A4(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT19), .B1(new_n284), .B2(G97), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n611), .A2(new_n606), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n287), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n378), .A2(new_n379), .A3(new_n373), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n626), .A2(new_n631), .A3(new_n632), .A4(new_n627), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(KEYINPUT85), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n323), .A2(new_n490), .B1(new_n254), .B2(new_n623), .ZN(new_n635));
  NOR2_X1   g0435(.A1(G238), .A2(G1698), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n636), .B1(new_n522), .B2(G1698), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n619), .B1(new_n637), .B2(new_n256), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n635), .B(G190), .C1(new_n638), .C2(new_n254), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT86), .ZN(new_n640));
  INV_X1    g0440(.A(new_n621), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT86), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n641), .A2(new_n642), .A3(G190), .A4(new_n635), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n628), .A2(new_n634), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n576), .A2(new_n374), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n614), .A2(new_n646), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n621), .A2(new_n625), .A3(G179), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n621), .A2(new_n625), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n648), .B1(new_n650), .B2(new_n404), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n645), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n561), .A2(new_n605), .A3(new_n653), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n467), .A2(new_n521), .A3(new_n654), .ZN(G372));
  INV_X1    g0455(.A(new_n401), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n370), .B1(new_n656), .B2(new_n406), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n657), .A2(new_n460), .ZN(new_n658));
  INV_X1    g0458(.A(new_n451), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n308), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT90), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT89), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n618), .A2(new_n620), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n662), .B1(new_n663), .B2(new_n390), .ZN(new_n664));
  AOI211_X1 g0464(.A(KEYINPUT89), .B(new_n254), .C1(new_n618), .C2(new_n620), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n635), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n404), .ZN(new_n667));
  INV_X1    g0467(.A(new_n648), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n661), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  AOI211_X1 g0469(.A(KEYINPUT90), .B(new_n648), .C1(new_n666), .C2(new_n404), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n647), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n614), .A2(new_n627), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n666), .A2(G200), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(new_n639), .A3(new_n673), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n596), .A2(new_n598), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n600), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n505), .A2(new_n677), .A3(new_n511), .A4(new_n516), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n581), .B1(new_n594), .B2(new_n254), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n494), .B1(new_n679), .B2(KEYINPUT88), .ZN(new_n680));
  AOI21_X1  g0480(.A(G200), .B1(new_n680), .B2(new_n595), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n597), .A2(G190), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n575), .B(new_n580), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n683), .A2(new_n560), .A3(new_n554), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n675), .A2(new_n678), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT26), .ZN(new_n686));
  INV_X1    g0486(.A(new_n560), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n671), .A2(new_n686), .A3(new_n687), .A4(new_n674), .ZN(new_n688));
  AOI22_X1  g0488(.A1(new_n555), .A2(new_n556), .B1(new_n534), .B2(new_n404), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n645), .A2(new_n559), .A3(new_n689), .A4(new_n652), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT26), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n688), .A2(new_n671), .A3(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n685), .A2(new_n692), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n660), .B(new_n466), .C1(new_n467), .C2(new_n693), .ZN(G369));
  NAND3_X1  g0494(.A1(new_n505), .A2(new_n511), .A3(new_n516), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n263), .A2(new_n214), .A3(G13), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G213), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(G343), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n510), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n695), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n521), .B2(new_n703), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n705), .A2(G330), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n605), .B1(new_n601), .B2(new_n702), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n677), .B2(new_n702), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n695), .A2(new_n702), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n605), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n599), .A2(new_n702), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n709), .A2(new_n714), .ZN(G399));
  NOR2_X1   g0515(.A1(new_n209), .A2(G41), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n610), .A2(G116), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(G1), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n218), .B2(new_n717), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT28), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n702), .B1(new_n685), .B2(new_n692), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT29), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n671), .A2(KEYINPUT26), .A3(new_n687), .A4(new_n674), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT93), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n690), .A2(new_n727), .A3(new_n686), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n727), .B1(new_n690), .B2(new_n686), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n671), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n685), .B1(new_n731), .B2(KEYINPUT94), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT94), .ZN(new_n733));
  OAI211_X1 g0533(.A(new_n733), .B(new_n671), .C1(new_n729), .C2(new_n730), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n701), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n725), .B1(new_n735), .B2(new_n724), .ZN(new_n736));
  INV_X1    g0536(.A(G330), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n683), .A2(new_n677), .A3(new_n652), .A4(new_n645), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n521), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n739), .A2(new_n740), .A3(new_n561), .A4(new_n702), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT92), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n554), .A2(new_n560), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n738), .A2(new_n521), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(KEYINPUT92), .A3(new_n702), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT30), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n514), .B(KEYINPUT91), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n680), .A2(new_n551), .A3(new_n649), .A4(new_n595), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT91), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n514), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n551), .A2(new_n649), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n602), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n753), .A2(new_n755), .A3(KEYINPUT30), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n517), .A2(G179), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n757), .A2(new_n534), .A3(new_n602), .A4(new_n666), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n751), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n701), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT31), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n759), .A2(KEYINPUT31), .A3(new_n701), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n737), .B1(new_n747), .B2(new_n764), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n736), .A2(new_n765), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n766), .A2(KEYINPUT95), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(KEYINPUT95), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n721), .B1(new_n769), .B2(G1), .ZN(G364));
  NOR2_X1   g0570(.A1(new_n705), .A2(G330), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n214), .A2(G13), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n263), .B1(new_n773), .B2(G45), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n771), .B(new_n706), .C1(new_n717), .C2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n774), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n716), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n256), .A2(new_n208), .ZN(new_n778));
  INV_X1    g0578(.A(G355), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n778), .A2(new_n779), .B1(G116), .B2(new_n208), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n209), .A2(new_n256), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(new_n489), .B2(new_n219), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n251), .A2(G45), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n780), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(G13), .A2(G33), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(G20), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n213), .B1(G20), .B2(new_n404), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n777), .B1(new_n785), .B2(new_n791), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n214), .A2(new_n385), .A3(G179), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n793), .A2(new_n395), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n794), .A2(KEYINPUT96), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(KEYINPUT96), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G283), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n214), .A2(new_n415), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n800), .A2(G190), .A3(new_n385), .ZN(new_n801));
  INV_X1    g0601(.A(G322), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(G190), .A2(G200), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G311), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n438), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n804), .A2(G20), .A3(new_n415), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n803), .B(new_n807), .C1(G329), .C2(new_n809), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n395), .A2(G179), .A3(G200), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n214), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n800), .A2(G200), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(G190), .ZN(new_n815));
  XNOR2_X1  g0615(.A(KEYINPUT33), .B(G317), .ZN(new_n816));
  AOI22_X1  g0616(.A1(G294), .A2(new_n813), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n793), .A2(G190), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n814), .A2(new_n395), .ZN(new_n820));
  XOR2_X1   g0620(.A(KEYINPUT97), .B(G326), .Z(new_n821));
  AOI22_X1  g0621(.A1(G303), .A2(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n810), .A2(new_n817), .A3(new_n822), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n256), .B1(new_n805), .B2(new_n258), .C1(new_n277), .C2(new_n801), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n808), .A2(new_n434), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT32), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n818), .A2(new_n609), .ZN(new_n828));
  NOR3_X1   g0628(.A1(new_n824), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n812), .A2(new_n471), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(G68), .B2(new_n815), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n820), .A2(G50), .B1(new_n825), .B2(new_n826), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n829), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n797), .A2(new_n543), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n799), .A2(new_n823), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT98), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n789), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(new_n835), .B2(new_n836), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n792), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n788), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n840), .B1(new_n705), .B2(new_n841), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT99), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n775), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(G396));
  NAND2_X1  g0645(.A1(new_n383), .A2(new_n701), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n406), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n397), .A2(new_n406), .A3(new_n846), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n722), .B(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(KEYINPUT92), .B1(new_n745), .B2(new_n702), .ZN(new_n851));
  NOR4_X1   g0651(.A1(new_n654), .A2(new_n742), .A3(new_n521), .A4(new_n701), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n764), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(G330), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n777), .B1(new_n850), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n854), .B2(new_n850), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n838), .A2(new_n787), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n777), .B1(G77), .B2(new_n857), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n815), .A2(KEYINPUT100), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n815), .A2(KEYINPUT100), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(G283), .ZN(new_n863));
  INV_X1    g0663(.A(new_n797), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(G87), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n801), .A2(new_n586), .B1(new_n805), .B2(new_n468), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n256), .B(new_n866), .C1(G311), .C2(new_n809), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n818), .A2(new_n543), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n830), .B(new_n868), .C1(G303), .C2(new_n820), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n863), .A2(new_n865), .A3(new_n867), .A4(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n438), .B1(new_n809), .B2(G132), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n297), .B2(new_n818), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n797), .A2(new_n362), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n872), .B(new_n873), .C1(G58), .C2(new_n813), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n875), .A2(KEYINPUT101), .ZN(new_n876));
  INV_X1    g0676(.A(new_n801), .ZN(new_n877));
  INV_X1    g0677(.A(new_n805), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n877), .A2(G143), .B1(new_n878), .B2(G159), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n815), .A2(G150), .ZN(new_n880));
  INV_X1    g0680(.A(G137), .ZN(new_n881));
  INV_X1    g0681(.A(new_n820), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n879), .B(new_n880), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT34), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT101), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n884), .B1(new_n874), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n870), .B1(new_n876), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n858), .B1(new_n887), .B2(new_n789), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n847), .A2(new_n848), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n888), .B1(new_n889), .B2(new_n787), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n856), .A2(new_n890), .ZN(G384));
  OR2_X1    g0691(.A1(new_n545), .A2(KEYINPUT35), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n545), .A2(KEYINPUT35), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n892), .A2(G116), .A3(new_n215), .A4(new_n893), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n894), .B(KEYINPUT36), .Z(new_n895));
  OAI211_X1 g0695(.A(new_n219), .B(G77), .C1(new_n277), .C2(new_n360), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n297), .A2(G68), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n263), .B(G13), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n659), .A2(new_n699), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n406), .A2(new_n701), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n722), .B2(new_n849), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n369), .A2(new_n701), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n370), .A2(new_n401), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT102), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT102), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n370), .A2(new_n401), .A3(new_n904), .A4(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n904), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n339), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n903), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT38), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n422), .A2(new_n447), .ZN(new_n915));
  INV_X1    g0715(.A(new_n699), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n447), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n915), .A2(new_n917), .A3(new_n455), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n918), .A2(KEYINPUT37), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n417), .A2(new_n419), .A3(new_n421), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n438), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n362), .B1(new_n431), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n423), .B1(new_n435), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n923), .A2(new_n443), .A3(new_n287), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n920), .B1(new_n924), .B2(new_n446), .ZN(new_n925));
  INV_X1    g0725(.A(new_n455), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT103), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT103), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n924), .A2(new_n446), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n928), .B(new_n455), .C1(new_n929), .C2(new_n920), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n929), .A2(new_n699), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n927), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n919), .B1(new_n933), .B2(KEYINPUT37), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n932), .B1(new_n451), .B2(new_n460), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n914), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n461), .A2(new_n931), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT37), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n455), .B1(new_n929), .B2(new_n920), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n931), .B1(new_n939), .B2(KEYINPUT103), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n938), .B1(new_n940), .B2(new_n930), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n937), .B(KEYINPUT38), .C1(new_n941), .C2(new_n919), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n936), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n900), .B1(new_n913), .B2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n917), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n457), .A2(KEYINPUT104), .A3(new_n458), .ZN(new_n947));
  INV_X1    g0747(.A(new_n450), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n422), .A2(new_n447), .A3(new_n448), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(KEYINPUT104), .B1(new_n457), .B2(new_n458), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n946), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n918), .A2(KEYINPUT37), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n918), .A2(KEYINPUT37), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(KEYINPUT38), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n933), .A2(KEYINPUT37), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n935), .B1(new_n957), .B2(new_n953), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n956), .A2(KEYINPUT105), .B1(new_n958), .B2(KEYINPUT38), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT105), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT104), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n459), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n962), .A2(new_n451), .A3(new_n947), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n963), .A2(new_n946), .B1(new_n953), .B2(new_n954), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n960), .B1(new_n964), .B2(KEYINPUT38), .ZN(new_n965));
  AOI21_X1  g0765(.A(KEYINPUT39), .B1(new_n959), .B2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT39), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n943), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n370), .A2(new_n701), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n945), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n660), .A2(new_n466), .ZN(new_n972));
  INV_X1    g0772(.A(new_n467), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n972), .B1(new_n736), .B2(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n971), .B(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT40), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n952), .A2(new_n955), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n977), .A2(KEYINPUT105), .A3(new_n914), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n965), .A2(new_n978), .A3(new_n942), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n762), .A2(new_n763), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n980), .B1(new_n743), .B2(new_n746), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n912), .A2(new_n889), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n976), .B1(new_n979), .B2(new_n983), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n906), .A2(new_n908), .B1(new_n339), .B2(new_n910), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n985), .A2(new_n849), .ZN(new_n986));
  AND4_X1   g0786(.A1(new_n976), .A2(new_n943), .A3(new_n853), .A4(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n467), .B2(new_n981), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n983), .A2(new_n976), .A3(new_n943), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n853), .A2(new_n986), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(new_n965), .B2(new_n959), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n990), .B1(new_n992), .B2(new_n976), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n993), .A2(new_n973), .A3(new_n853), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n989), .A2(new_n994), .A3(G330), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n975), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n263), .B2(new_n773), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n975), .A2(new_n995), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n899), .B1(new_n997), .B2(new_n998), .ZN(G367));
  OAI21_X1  g0799(.A(new_n561), .B1(new_n550), .B2(new_n702), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n687), .A2(new_n701), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n714), .A2(KEYINPUT45), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT45), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1002), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1004), .B1(new_n713), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g0807(.A(KEYINPUT108), .B(KEYINPUT44), .C1(new_n714), .C2(new_n1002), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1002), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1010), .A2(new_n713), .A3(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1007), .A2(new_n1008), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n709), .ZN(new_n1014));
  OAI21_X1  g0814(.A(KEYINPUT109), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1013), .A2(KEYINPUT109), .A3(new_n1014), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n711), .B1(new_n708), .B2(new_n710), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(new_n706), .Z(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n1020), .A2(new_n1023), .B1(new_n767), .B2(new_n768), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n716), .B(KEYINPUT41), .Z(new_n1025));
  OAI21_X1  g0825(.A(new_n774), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1005), .A2(new_n711), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1027), .A2(KEYINPUT42), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(KEYINPUT42), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n560), .B1(new_n1000), .B2(new_n677), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n1028), .A2(new_n1029), .B1(new_n702), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT106), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n672), .A2(new_n702), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1033), .B(new_n647), .C1(new_n669), .C2(new_n670), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n671), .A2(new_n674), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1032), .B(new_n1034), .C1(new_n1035), .C2(new_n1033), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT43), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1037), .B(new_n1038), .ZN(new_n1039));
  OR3_X1    g0839(.A1(new_n1031), .A2(KEYINPUT107), .A3(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(KEYINPUT107), .B1(new_n1031), .B2(new_n1039), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1031), .A2(new_n1038), .A3(new_n1037), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n709), .A2(new_n1005), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1043), .B(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1026), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n862), .A2(G294), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n864), .A2(G97), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n882), .A2(new_n806), .B1(new_n543), .B2(new_n812), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n438), .B1(new_n801), .B2(new_n497), .ZN(new_n1050));
  INV_X1    g0850(.A(G317), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n805), .A2(new_n798), .B1(new_n808), .B2(new_n1051), .ZN(new_n1052));
  NOR3_X1   g0852(.A1(new_n1049), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n819), .A2(G116), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT46), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1047), .A2(new_n1048), .A3(new_n1053), .A4(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(G143), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n882), .A2(new_n1057), .B1(new_n277), .B2(new_n818), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n877), .A2(G150), .B1(G137), .B2(new_n809), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n297), .B2(new_n805), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n1058), .B(new_n1060), .C1(G68), .C2(new_n813), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n864), .A2(G77), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1062), .A2(KEYINPUT110), .A3(new_n256), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1061), .B(new_n1063), .C1(new_n434), .C2(new_n861), .ZN(new_n1064));
  AOI21_X1  g0864(.A(KEYINPUT110), .B1(new_n1062), .B2(new_n256), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1056), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT47), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n789), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1037), .A2(new_n788), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n791), .B1(new_n209), .B2(new_n374), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n243), .A2(new_n781), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n716), .B(new_n776), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  AND3_X1   g0872(.A1(new_n1068), .A2(new_n1069), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1046), .A2(new_n1074), .ZN(G387));
  OAI21_X1  g0875(.A(KEYINPUT112), .B1(new_n769), .B2(new_n1023), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1022), .B1(new_n767), .B2(new_n768), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT112), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n767), .A2(new_n1079), .A3(new_n768), .A4(new_n1022), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1076), .A2(new_n1078), .A3(new_n716), .A4(new_n1080), .ZN(new_n1081));
  OR2_X1    g0881(.A1(new_n708), .A2(new_n841), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n778), .A2(new_n718), .B1(G107), .B2(new_n208), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n240), .A2(new_n489), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n718), .ZN(new_n1085));
  AOI211_X1 g0885(.A(G45), .B(new_n1085), .C1(G68), .C2(G77), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n274), .A2(G50), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT50), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n782), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1083), .B1(new_n1084), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n777), .B1(new_n1090), .B2(new_n791), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT111), .Z(new_n1092));
  AOI22_X1  g0892(.A1(new_n877), .A2(G317), .B1(new_n878), .B2(G303), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1093), .B1(new_n802), .B2(new_n882), .C1(new_n861), .C2(new_n806), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT48), .ZN(new_n1095));
  OR2_X1    g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n819), .A2(G294), .B1(new_n813), .B2(G283), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT49), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n864), .A2(G116), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n256), .B1(new_n809), .B2(new_n821), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n812), .A2(new_n373), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n818), .A2(new_n258), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1106), .B(new_n1107), .C1(G159), .C2(new_n820), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n279), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n815), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n801), .A2(new_n297), .B1(new_n805), .B2(new_n362), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n438), .B(new_n1111), .C1(G150), .C2(new_n809), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1048), .A2(new_n1108), .A3(new_n1110), .A4(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1105), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1092), .B1(new_n1114), .B2(new_n789), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1023), .A2(new_n776), .B1(new_n1082), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1081), .A2(new_n1116), .ZN(G393));
  XNOR2_X1  g0917(.A(new_n1013), .B(new_n709), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n776), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n248), .A2(new_n782), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n790), .B1(new_n471), .B2(new_n208), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n777), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(G317), .A2(new_n820), .B1(new_n877), .B2(G311), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT52), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n438), .B1(new_n805), .B2(new_n586), .C1(new_n812), .C2(new_n468), .ZN(new_n1125));
  OR3_X1    g0925(.A1(new_n1124), .A2(new_n834), .A3(new_n1125), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n818), .A2(new_n798), .B1(new_n802), .B2(new_n808), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n862), .A2(G303), .B1(KEYINPUT113), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(KEYINPUT113), .B2(new_n1127), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(G150), .A2(new_n820), .B1(new_n877), .B2(G159), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT51), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n862), .A2(G50), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n256), .B1(new_n808), .B2(new_n1057), .C1(new_n805), .C2(new_n274), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n812), .A2(new_n258), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(new_n224), .B2(new_n819), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1132), .A2(new_n865), .A3(new_n1134), .A4(new_n1136), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n1126), .A2(new_n1129), .B1(new_n1131), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1122), .B1(new_n1138), .B2(new_n789), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n1002), .B2(new_n841), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1119), .A2(new_n1140), .ZN(new_n1141));
  OR2_X1    g0941(.A1(new_n1077), .A2(new_n1118), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n717), .B1(new_n1077), .B2(new_n1020), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1141), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(G390));
  OAI21_X1  g0945(.A(new_n777), .B1(new_n1109), .B2(new_n857), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n873), .B1(G107), .B2(new_n862), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n801), .A2(new_n468), .B1(new_n586), .B2(new_n808), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n256), .B(new_n1148), .C1(G97), .C2(new_n878), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n1135), .B(new_n828), .C1(G283), .C2(new_n820), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1147), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n818), .A2(new_n271), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT53), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n438), .B1(new_n809), .B2(G125), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(KEYINPUT54), .B(G143), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n877), .A2(G132), .B1(new_n878), .B2(new_n1156), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(G159), .A2(new_n813), .B1(new_n820), .B2(G128), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1153), .A2(new_n1154), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n861), .A2(new_n881), .B1(new_n797), .B2(new_n297), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1151), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1146), .B1(new_n1161), .B2(new_n789), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n969), .B2(new_n787), .ZN(new_n1163));
  NOR4_X1   g0963(.A1(new_n981), .A2(new_n737), .A3(new_n849), .A4(new_n985), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n970), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n979), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n731), .A2(KEYINPUT94), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n685), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1167), .A2(new_n1168), .A3(new_n734), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1169), .A2(new_n702), .A3(new_n889), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n902), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1166), .B1(new_n1171), .B2(new_n912), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n979), .A2(new_n967), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n944), .A2(KEYINPUT39), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n1173), .A2(new_n1174), .B1(new_n1165), .B2(new_n913), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1164), .B1(new_n1172), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n970), .B1(new_n959), .B2(new_n965), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n901), .B1(new_n735), .B2(new_n889), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1177), .B1(new_n1178), .B2(new_n985), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n913), .A2(new_n1165), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n966), .B2(new_n968), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n853), .A2(G330), .A3(new_n889), .A4(new_n912), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1179), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1176), .A2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1163), .B1(new_n1184), .B2(new_n774), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n1172), .A2(new_n1175), .A3(new_n1164), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1182), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT115), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n854), .A2(new_n467), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n972), .B(new_n1190), .C1(new_n736), .C2(new_n973), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n912), .B1(new_n765), .B2(new_n889), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n903), .B1(new_n1192), .B2(new_n1164), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n853), .A2(G330), .A3(new_n889), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n985), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1195), .A2(new_n902), .A3(new_n1170), .A4(new_n1182), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT114), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1193), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1178), .A2(KEYINPUT114), .A3(new_n1182), .A4(new_n1195), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n1191), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1188), .A2(new_n1189), .A3(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1191), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1202));
  OAI21_X1  g1002(.A(KEYINPUT115), .B1(new_n1184), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1201), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n717), .B1(new_n1184), .B2(new_n1202), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1185), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(G378));
  NAND2_X1  g1007(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n900), .B1(new_n944), .B2(new_n913), .C1(new_n1208), .C2(new_n1165), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n301), .A2(new_n916), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n308), .A2(new_n466), .A3(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1212), .B1(new_n308), .B2(new_n466), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1211), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1215), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1217), .A2(new_n1213), .A3(new_n1210), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n993), .B2(G330), .ZN(new_n1220));
  OAI211_X1 g1020(.A(G330), .B(new_n1219), .C1(new_n984), .C2(new_n987), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1209), .B1(new_n1220), .B2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1219), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n988), .B2(new_n737), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1225), .A2(new_n971), .A3(new_n1221), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1223), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n776), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n777), .B1(G50), .B2(new_n857), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n256), .A2(G41), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(G33), .A2(G41), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n1230), .A2(G50), .A3(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n864), .A2(G58), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1230), .B1(new_n373), .B2(new_n805), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n801), .A2(new_n543), .B1(new_n798), .B2(new_n808), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1107), .B1(G68), .B2(new_n813), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n815), .A2(G97), .B1(new_n820), .B2(G116), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1233), .A2(new_n1236), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  XOR2_X1   g1039(.A(new_n1239), .B(KEYINPUT116), .Z(new_n1240));
  INV_X1    g1040(.A(KEYINPUT58), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1232), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  XOR2_X1   g1042(.A(new_n1242), .B(KEYINPUT117), .Z(new_n1243));
  INV_X1    g1043(.A(G128), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n801), .A2(new_n1244), .B1(new_n805), .B2(new_n881), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n819), .A2(new_n1156), .B1(new_n815), .B2(G132), .ZN(new_n1246));
  INV_X1    g1046(.A(G125), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1246), .B1(new_n1247), .B2(new_n882), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1245), .B(new_n1248), .C1(G150), .C2(new_n813), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT59), .ZN(new_n1250));
  OR2_X1    g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n809), .A2(G124), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1231), .B(new_n1252), .C1(new_n797), .C2(new_n434), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT118), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1256));
  OR2_X1    g1056(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1251), .A2(new_n1255), .A3(new_n1256), .A4(new_n1257), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1243), .B(new_n1258), .C1(new_n1241), .C2(new_n1240), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1229), .B1(new_n1259), .B2(new_n789), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n1219), .B2(new_n787), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1228), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1189), .B1(new_n1188), .B2(new_n1200), .ZN(new_n1264));
  NOR3_X1   g1064(.A1(new_n1184), .A2(new_n1202), .A3(KEYINPUT115), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1191), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(KEYINPUT57), .B1(new_n1266), .B2(new_n1227), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1191), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT119), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1223), .A2(new_n1270), .A3(new_n1226), .ZN(new_n1271));
  OAI211_X1 g1071(.A(KEYINPUT119), .B(new_n1209), .C1(new_n1220), .C2(new_n1222), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1271), .A2(KEYINPUT57), .A3(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n716), .B1(new_n1269), .B2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1263), .B1(new_n1267), .B2(new_n1274), .ZN(G375));
  NAND2_X1  g1075(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1268), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1025), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1277), .A2(new_n1278), .A3(new_n1202), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1198), .A2(new_n776), .A3(new_n1199), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n777), .B1(G68), .B2(new_n857), .ZN(new_n1281));
  OAI221_X1 g1081(.A(new_n438), .B1(new_n805), .B2(new_n543), .C1(new_n798), .C2(new_n801), .ZN(new_n1282));
  AOI211_X1 g1082(.A(new_n1106), .B(new_n1282), .C1(G294), .C2(new_n820), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n862), .A2(G116), .ZN(new_n1284));
  OAI22_X1  g1084(.A1(new_n818), .A2(new_n471), .B1(new_n497), .B2(new_n808), .ZN(new_n1285));
  XOR2_X1   g1085(.A(new_n1285), .B(KEYINPUT120), .Z(new_n1286));
  NAND4_X1  g1086(.A1(new_n1283), .A2(new_n1284), .A3(new_n1062), .A4(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n256), .B1(new_n808), .B2(new_n1244), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1288), .B1(G150), .B2(new_n878), .ZN(new_n1289));
  AOI22_X1  g1089(.A1(new_n819), .A2(G159), .B1(new_n813), .B2(G50), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1233), .A2(new_n1289), .A3(new_n1290), .ZN(new_n1291));
  XOR2_X1   g1091(.A(new_n1291), .B(KEYINPUT121), .Z(new_n1292));
  AOI22_X1  g1092(.A1(G132), .A2(new_n820), .B1(new_n877), .B2(G137), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1293), .B1(new_n861), .B2(new_n1155), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1287), .B1(new_n1292), .B2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1281), .B1(new_n1295), .B2(new_n789), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1296), .B1(new_n912), .B2(new_n787), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1279), .A2(new_n1280), .A3(new_n1297), .ZN(G381));
  NOR3_X1   g1098(.A1(G390), .A2(G384), .A3(G381), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1073), .B1(new_n1026), .B2(new_n1045), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1081), .A2(new_n844), .A3(new_n1116), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1299), .A2(new_n1300), .A3(new_n1206), .A4(new_n1302), .ZN(new_n1303));
  OR2_X1    g1103(.A1(new_n1303), .A2(G375), .ZN(G407));
  NAND2_X1  g1104(.A1(new_n700), .A2(G213), .ZN(new_n1305));
  OR3_X1    g1105(.A1(G375), .A2(G378), .A3(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(G407), .A2(G213), .A3(new_n1306), .ZN(G409));
  NAND2_X1  g1107(.A1(G387), .A2(new_n1144), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(G390), .A2(new_n1300), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(G393), .A2(G396), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n1301), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1310), .A2(new_n1312), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1308), .A2(new_n1309), .A3(new_n1301), .A4(new_n1311), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT125), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT61), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n700), .A2(G213), .A3(G2897), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT60), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1277), .B1(new_n1200), .B2(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1276), .A2(new_n1268), .A3(KEYINPUT60), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1320), .A2(new_n716), .A3(new_n1321), .ZN(new_n1322));
  OR2_X1    g1122(.A1(G384), .A2(KEYINPUT122), .ZN(new_n1323));
  AND3_X1   g1123(.A1(new_n1323), .A2(new_n1280), .A3(new_n1297), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1322), .A2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1325), .A2(KEYINPUT122), .A3(G384), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(G384), .A2(KEYINPUT122), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1322), .A2(new_n1324), .A3(new_n1327), .ZN(new_n1328));
  AOI211_X1 g1128(.A(KEYINPUT123), .B(new_n1318), .C1(new_n1326), .C2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1318), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1326), .A2(new_n1328), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT123), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1330), .B1(new_n1331), .B2(new_n1332), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1326), .A2(KEYINPUT123), .A3(new_n1328), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1329), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  OAI211_X1 g1135(.A(G378), .B(new_n1263), .C1(new_n1267), .C2(new_n1274), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1227), .ZN(new_n1337));
  NOR3_X1   g1137(.A1(new_n1269), .A2(new_n1025), .A3(new_n1337), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1271), .A2(new_n776), .A3(new_n1272), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1339), .A2(new_n1261), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1206), .B1(new_n1338), .B2(new_n1340), .ZN(new_n1341));
  AOI22_X1  g1141(.A1(new_n1336), .A2(new_n1341), .B1(G213), .B2(new_n700), .ZN(new_n1342));
  OAI211_X1 g1142(.A(new_n1316), .B(new_n1317), .C1(new_n1335), .C2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1342), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1331), .ZN(new_n1345));
  OAI21_X1  g1145(.A(KEYINPUT62), .B1(new_n1344), .B2(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT62), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1342), .A2(new_n1347), .A3(new_n1331), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1343), .A2(new_n1346), .A3(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1350), .A2(new_n1318), .A3(new_n1334), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1329), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1351), .A2(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1353), .A2(new_n1344), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1316), .B1(new_n1354), .B2(new_n1317), .ZN(new_n1355));
  OAI21_X1  g1155(.A(new_n1315), .B1(new_n1349), .B2(new_n1355), .ZN(new_n1356));
  NOR2_X1   g1156(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1357));
  OR2_X1    g1157(.A1(new_n1357), .A2(KEYINPUT63), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1313), .A2(new_n1317), .A3(new_n1314), .ZN(new_n1359));
  XNOR2_X1  g1159(.A(new_n1359), .B(KEYINPUT124), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1357), .A2(KEYINPUT63), .ZN(new_n1361));
  NAND4_X1  g1161(.A1(new_n1358), .A2(new_n1360), .A3(new_n1354), .A4(new_n1361), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1356), .A2(new_n1362), .ZN(G405));
  INV_X1    g1163(.A(KEYINPUT127), .ZN(new_n1364));
  AND3_X1   g1164(.A1(new_n1271), .A2(KEYINPUT57), .A3(new_n1272), .ZN(new_n1365));
  AOI21_X1  g1165(.A(new_n717), .B1(new_n1266), .B2(new_n1365), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT57), .ZN(new_n1367));
  OAI21_X1  g1167(.A(new_n1367), .B1(new_n1269), .B2(new_n1337), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1366), .A2(new_n1368), .ZN(new_n1369));
  AOI21_X1  g1169(.A(G378), .B1(new_n1369), .B2(new_n1263), .ZN(new_n1370));
  AOI211_X1 g1170(.A(new_n1206), .B(new_n1262), .C1(new_n1366), .C2(new_n1368), .ZN(new_n1371));
  OAI21_X1  g1171(.A(new_n1331), .B1(new_n1370), .B2(new_n1371), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(G375), .A2(new_n1206), .ZN(new_n1373));
  NAND3_X1  g1173(.A1(new_n1373), .A2(new_n1336), .A3(new_n1345), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1372), .A2(new_n1374), .ZN(new_n1375));
  AOI21_X1  g1175(.A(new_n1364), .B1(new_n1375), .B2(KEYINPUT126), .ZN(new_n1376));
  INV_X1    g1176(.A(KEYINPUT126), .ZN(new_n1377));
  AOI211_X1 g1177(.A(new_n1377), .B(KEYINPUT127), .C1(new_n1372), .C2(new_n1374), .ZN(new_n1378));
  NAND3_X1  g1178(.A1(new_n1372), .A2(new_n1377), .A3(new_n1374), .ZN(new_n1379));
  INV_X1    g1179(.A(new_n1315), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1379), .A2(new_n1380), .ZN(new_n1381));
  NOR3_X1   g1181(.A1(new_n1376), .A2(new_n1378), .A3(new_n1381), .ZN(new_n1382));
  AND3_X1   g1182(.A1(new_n1373), .A2(new_n1336), .A3(new_n1345), .ZN(new_n1383));
  AOI21_X1  g1183(.A(new_n1345), .B1(new_n1373), .B2(new_n1336), .ZN(new_n1384));
  OAI21_X1  g1184(.A(KEYINPUT126), .B1(new_n1383), .B2(new_n1384), .ZN(new_n1385));
  NAND2_X1  g1185(.A1(new_n1385), .A2(KEYINPUT127), .ZN(new_n1386));
  NAND3_X1  g1186(.A1(new_n1375), .A2(KEYINPUT126), .A3(new_n1364), .ZN(new_n1387));
  AOI22_X1  g1187(.A1(new_n1386), .A2(new_n1387), .B1(new_n1380), .B2(new_n1379), .ZN(new_n1388));
  NOR2_X1   g1188(.A1(new_n1382), .A2(new_n1388), .ZN(G402));
endmodule


