//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 1 1 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n554, new_n555, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n571, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n615, new_n617, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1234, new_n1235, new_n1236;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT64), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT65), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(new_n466), .A3(G125), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n460), .B1(new_n462), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n469));
  NAND2_X1  g044(.A1(G101), .A2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT3), .B(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n471), .B1(new_n472), .B2(G137), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n469), .B1(new_n473), .B2(G2105), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n464), .A2(new_n466), .A3(G137), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(new_n470), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n476), .A2(KEYINPUT66), .A3(new_n460), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n468), .B1(new_n474), .B2(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n464), .A2(new_n466), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(new_n460), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(new_n481), .A2(KEYINPUT68), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(KEYINPUT68), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n479), .A2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT67), .ZN(new_n487));
  NOR2_X1   g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT69), .ZN(new_n489));
  INV_X1    g064(.A(G112), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n463), .B1(new_n490), .B2(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n484), .A2(new_n487), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  NAND4_X1  g069(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n460), .ZN(new_n495));
  XOR2_X1   g070(.A(KEYINPUT70), .B(KEYINPUT4), .Z(new_n496));
  AND2_X1   g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AND3_X1   g072(.A1(KEYINPUT70), .A2(KEYINPUT4), .A3(G138), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(new_n464), .A3(new_n466), .ZN(new_n499));
  NAND2_X1  g074(.A1(G102), .A2(G2104), .ZN(new_n500));
  AOI21_X1  g075(.A(G2105), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n464), .A2(new_n466), .A3(G126), .ZN(new_n502));
  NAND2_X1  g077(.A1(G114), .A2(G2104), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n460), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR3_X1   g079(.A1(new_n497), .A2(new_n501), .A3(new_n504), .ZN(G164));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT71), .B1(new_n506), .B2(KEYINPUT6), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n508), .A2(new_n509), .A3(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n506), .A2(KEYINPUT6), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  AND3_X1   g094(.A1(new_n511), .A2(G543), .A3(new_n512), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n519), .A2(G88), .B1(new_n520), .B2(G50), .ZN(new_n521));
  NAND2_X1  g096(.A1(G75), .A2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G62), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n522), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G651), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT72), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n524), .A2(KEYINPUT72), .A3(G651), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n521), .A2(new_n527), .A3(new_n528), .ZN(G166));
  XNOR2_X1  g104(.A(KEYINPUT73), .B(KEYINPUT7), .ZN(new_n530));
  AND3_X1   g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n530), .B(new_n531), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n507), .A2(new_n510), .B1(KEYINPUT6), .B2(new_n506), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n533), .A2(G51), .A3(G543), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n533), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n535));
  OAI211_X1 g110(.A(new_n532), .B(new_n534), .C1(new_n535), .C2(new_n518), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n518), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G651), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n515), .A2(new_n517), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n533), .A2(G90), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n533), .A2(G52), .A3(G543), .ZN(new_n544));
  AND3_X1   g119(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(G171));
  NAND2_X1  g120(.A1(G68), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G56), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n518), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G651), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n533), .A2(G43), .A3(G543), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n533), .A2(G81), .A3(new_n542), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n551), .A2(G860), .A3(new_n552), .ZN(G153));
  AND3_X1   g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(new_n555));
  XOR2_X1   g130(.A(new_n555), .B(KEYINPUT74), .Z(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n554), .A2(new_n558), .ZN(G188));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n518), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n519), .A2(G91), .B1(G651), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n511), .A2(G543), .A3(new_n512), .ZN(new_n565));
  INV_X1    g140(.A(G53), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n520), .A2(KEYINPUT9), .A3(G53), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n563), .A2(new_n567), .A3(new_n568), .ZN(G299));
  NAND3_X1  g144(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(G301));
  AND2_X1   g145(.A1(new_n527), .A2(new_n528), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(new_n521), .ZN(G303));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n573));
  OAI211_X1 g148(.A(new_n573), .B(G651), .C1(new_n542), .C2(G74), .ZN(new_n574));
  AOI21_X1  g149(.A(G74), .B1(new_n515), .B2(new_n517), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT75), .B1(new_n575), .B2(new_n506), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n533), .A2(G87), .A3(new_n542), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n533), .A2(G49), .A3(G543), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G288));
  INV_X1    g155(.A(G48), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT77), .B1(new_n565), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n533), .A2(G86), .A3(new_n542), .ZN(new_n583));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT76), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n515), .A2(new_n517), .A3(G61), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G651), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT77), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n533), .A2(new_n589), .A3(G48), .A4(G543), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n582), .A2(new_n583), .A3(new_n588), .A4(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n542), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n592), .A2(new_n506), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n519), .A2(G85), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n520), .A2(G47), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n519), .A2(new_n598), .A3(G92), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n518), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n520), .A2(G54), .B1(G651), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n533), .A2(new_n542), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(KEYINPUT10), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n599), .A2(new_n603), .A3(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n597), .B1(new_n608), .B2(G868), .ZN(G284));
  OAI21_X1  g184(.A(new_n597), .B1(new_n608), .B2(G868), .ZN(G321));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(G299), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(new_n611), .B2(G168), .ZN(G297));
  OAI21_X1  g188(.A(new_n612), .B1(new_n611), .B2(G168), .ZN(G280));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n608), .B1(new_n615), .B2(G860), .ZN(G148));
  NAND3_X1  g191(.A1(new_n549), .A2(new_n552), .A3(new_n550), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n608), .A2(new_n615), .ZN(new_n618));
  MUX2_X1   g193(.A(new_n617), .B(new_n618), .S(G868), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT78), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n485), .A2(G2104), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT12), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  XOR2_X1   g199(.A(KEYINPUT79), .B(G2100), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n480), .A2(G123), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n485), .A2(G135), .ZN(new_n628));
  NOR2_X1   g203(.A1(G99), .A2(G2105), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(new_n460), .B2(G111), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n627), .B(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT80), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2096), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n626), .A2(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2435), .ZN(new_n636));
  XOR2_X1   g211(.A(G2427), .B(G2438), .Z(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n636), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(new_n640), .A3(KEYINPUT14), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2451), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2454), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n643), .A2(new_n647), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G1341), .B(G1348), .Z(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  OAI21_X1  g227(.A(KEYINPUT82), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(G14), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n654), .B1(new_n650), .B2(new_n652), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT82), .ZN(new_n656));
  NAND4_X1  g231(.A1(new_n648), .A2(new_n649), .A3(new_n656), .A4(new_n651), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n653), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(G401));
  XOR2_X1   g234(.A(G2072), .B(G2078), .Z(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2067), .B(G2678), .Z(new_n663));
  OR2_X1    g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT83), .B(KEYINPUT18), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n660), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT84), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2096), .B(G2100), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT17), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(new_n662), .B2(new_n663), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n665), .B1(new_n664), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n669), .B(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G227));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT85), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT19), .Z(new_n677));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  AND2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT20), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n678), .A2(new_n679), .ZN(new_n683));
  AOI22_X1  g258(.A1(new_n681), .A2(new_n682), .B1(new_n677), .B2(new_n683), .ZN(new_n684));
  OR3_X1    g259(.A1(new_n677), .A2(new_n680), .A3(new_n683), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n684), .B(new_n685), .C1(new_n682), .C2(new_n681), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT21), .B(G1986), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n688), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT22), .B(G1981), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n691), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(G229));
  INV_X1    g270(.A(G29), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G27), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G164), .B2(new_n696), .ZN(new_n698));
  INV_X1    g273(.A(G2078), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT92), .B(G28), .ZN(new_n701));
  AOI21_X1  g276(.A(G29), .B1(new_n701), .B2(KEYINPUT30), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT93), .Z(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(KEYINPUT30), .B2(new_n701), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  MUX2_X1   g280(.A(G19), .B(new_n617), .S(G16), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G1341), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT27), .B(G1996), .Z(new_n708));
  NAND2_X1  g283(.A1(new_n472), .A2(G2105), .ZN(new_n709));
  INV_X1    g284(.A(G129), .ZN(new_n710));
  OR3_X1    g285(.A1(new_n709), .A2(KEYINPUT91), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(KEYINPUT91), .B1(new_n709), .B2(new_n710), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n472), .A2(G141), .B1(G105), .B2(G2104), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n714), .A2(G2105), .ZN(new_n715));
  NAND3_X1  g290(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT26), .Z(new_n717));
  NAND3_X1  g292(.A1(new_n713), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G29), .ZN(new_n720));
  OR2_X1    g295(.A1(G29), .A2(G32), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n708), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NOR3_X1   g297(.A1(new_n705), .A2(new_n707), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(G160), .A2(G29), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT24), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n696), .B1(new_n725), .B2(G34), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n726), .A2(KEYINPUT90), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n725), .A2(G34), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n726), .A2(KEYINPUT90), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n724), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G2084), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OR2_X1    g308(.A1(G5), .A2(G16), .ZN(new_n734));
  INV_X1    g309(.A(G16), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(G301), .B2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G1961), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n721), .B(new_n708), .C1(new_n718), .C2(new_n696), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n733), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT94), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n733), .A2(new_n739), .A3(KEYINPUT94), .A4(new_n738), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G2067), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT28), .ZN(new_n746));
  INV_X1    g321(.A(G26), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n746), .B1(new_n747), .B2(G29), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n747), .A2(G29), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n480), .A2(KEYINPUT88), .A3(G128), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT88), .ZN(new_n751));
  INV_X1    g326(.A(G128), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n751), .B1(new_n709), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n485), .A2(G140), .ZN(new_n754));
  OR2_X1    g329(.A1(G104), .A2(G2105), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n755), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n750), .A2(new_n753), .A3(new_n754), .A4(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n749), .B1(new_n757), .B2(G29), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n745), .B(new_n748), .C1(new_n758), .C2(new_n746), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n748), .B1(new_n758), .B2(new_n746), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(G2067), .ZN(new_n761));
  OR2_X1    g336(.A1(G16), .A2(G21), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G286), .B2(new_n735), .ZN(new_n763));
  INV_X1    g338(.A(G1966), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n736), .A2(new_n737), .ZN(new_n766));
  AND4_X1   g341(.A1(new_n759), .A2(new_n761), .A3(new_n765), .A4(new_n766), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n631), .A2(new_n696), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n723), .A2(new_n744), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  OR2_X1    g344(.A1(G4), .A2(G16), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n607), .B2(new_n735), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT87), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G1348), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n696), .A2(G33), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT25), .Z(new_n776));
  NAND2_X1  g351(.A1(new_n485), .A2(G139), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n472), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n776), .B(new_n777), .C1(new_n460), .C2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n774), .B1(new_n779), .B2(G29), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT89), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n781), .A2(G2072), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n763), .A2(new_n764), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n781), .A2(G2072), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n769), .A2(new_n773), .A3(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT34), .ZN(new_n787));
  OR2_X1    g362(.A1(G16), .A2(G23), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G288), .B2(new_n735), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT33), .B(G1976), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n735), .B1(new_n571), .B2(new_n521), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n735), .A2(G22), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(G1971), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(G1971), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n796), .B(new_n793), .C1(G166), .C2(new_n735), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n791), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n735), .A2(G6), .ZN(new_n799));
  INV_X1    g374(.A(G305), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n735), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT32), .B(G1981), .Z(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n801), .B(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n787), .B1(new_n798), .B2(new_n804), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n795), .A2(new_n797), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n801), .B(new_n802), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n806), .A2(new_n807), .A3(KEYINPUT34), .A4(new_n791), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT86), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT36), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n735), .A2(G24), .ZN(new_n813));
  INV_X1    g388(.A(G290), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(new_n735), .ZN(new_n815));
  INV_X1    g390(.A(G1986), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n696), .A2(G25), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n480), .A2(G119), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n485), .A2(G131), .ZN(new_n820));
  OR2_X1    g395(.A1(G95), .A2(G2105), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n821), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n819), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n818), .B1(new_n824), .B2(new_n696), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT35), .B(G1991), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n809), .A2(new_n812), .A3(new_n817), .A4(new_n827), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n696), .A2(G35), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(new_n493), .B2(G29), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT29), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n482), .A2(new_n483), .B1(new_n491), .B2(new_n489), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n696), .B1(new_n833), .B2(new_n487), .ZN(new_n834));
  OAI21_X1  g409(.A(KEYINPUT29), .B1(new_n834), .B2(new_n829), .ZN(new_n835));
  AND3_X1   g410(.A1(new_n832), .A2(new_n835), .A3(G2090), .ZN(new_n836));
  AOI21_X1  g411(.A(G2090), .B1(new_n832), .B2(new_n835), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  AND3_X1   g414(.A1(new_n786), .A2(new_n828), .A3(new_n839), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT31), .B(G11), .Z(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n724), .A2(G2084), .A3(new_n730), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n809), .A2(new_n817), .A3(new_n827), .ZN(new_n844));
  INV_X1    g419(.A(new_n812), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n810), .A2(new_n811), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n840), .A2(new_n842), .A3(new_n843), .A4(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(G299), .A2(G16), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n735), .A2(KEYINPUT23), .A3(G20), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT23), .ZN(new_n851));
  INV_X1    g426(.A(G20), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n851), .B1(new_n852), .B2(G16), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n849), .A2(new_n850), .A3(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(G1956), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n848), .A2(new_n855), .ZN(G311));
  INV_X1    g431(.A(KEYINPUT95), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n848), .B2(new_n855), .ZN(new_n858));
  NOR4_X1   g433(.A1(new_n769), .A2(new_n773), .A3(new_n838), .A4(new_n785), .ZN(new_n859));
  AND4_X1   g434(.A1(new_n843), .A2(new_n847), .A3(new_n859), .A4(new_n828), .ZN(new_n860));
  INV_X1    g435(.A(new_n855), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n860), .A2(KEYINPUT95), .A3(new_n861), .A4(new_n842), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n858), .A2(new_n862), .ZN(G150));
  NOR2_X1   g438(.A1(new_n607), .A2(new_n615), .ZN(new_n864));
  XNOR2_X1  g439(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(G80), .A2(G543), .ZN(new_n867));
  INV_X1    g442(.A(G67), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n867), .B1(new_n518), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(G651), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n533), .A2(G93), .A3(new_n542), .ZN(new_n871));
  INV_X1    g446(.A(G55), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n870), .B(new_n871), .C1(new_n872), .C2(new_n565), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n873), .A2(new_n551), .A3(new_n552), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n520), .A2(G55), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n617), .A2(new_n871), .A3(new_n870), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n866), .B(new_n877), .Z(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(KEYINPUT39), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT97), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n879), .B(new_n880), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n878), .A2(KEYINPUT39), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n882), .A2(G860), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n873), .A2(G860), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(KEYINPUT37), .Z(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT98), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n884), .A2(KEYINPUT98), .A3(new_n886), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(G145));
  XNOR2_X1  g466(.A(new_n493), .B(new_n631), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(G160), .ZN(new_n893));
  INV_X1    g468(.A(G130), .ZN(new_n894));
  OR3_X1    g469(.A1(new_n709), .A2(KEYINPUT99), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(KEYINPUT99), .B1(new_n709), .B2(new_n894), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n485), .A2(G142), .ZN(new_n897));
  OR2_X1    g472(.A1(G106), .A2(G2105), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n898), .B(G2104), .C1(G118), .C2(new_n460), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n895), .A2(new_n896), .A3(new_n897), .A4(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(new_n823), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT100), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n901), .A2(new_n902), .ZN(new_n904));
  INV_X1    g479(.A(new_n623), .ZN(new_n905));
  OR3_X1    g480(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n905), .B1(new_n903), .B2(new_n904), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(KEYINPUT101), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n499), .A2(new_n500), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n460), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n502), .A2(new_n503), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(G2105), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n495), .A2(new_n496), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n910), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n757), .B(new_n914), .ZN(new_n915));
  OR2_X1    g490(.A1(new_n915), .A2(new_n779), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n779), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(new_n718), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n908), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n908), .A2(new_n919), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n893), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G37), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n906), .A2(new_n907), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(new_n919), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n922), .B(new_n923), .C1(new_n893), .C2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g502(.A(new_n618), .B(new_n877), .Z(new_n928));
  OR2_X1    g503(.A1(G299), .A2(new_n607), .ZN(new_n929));
  NAND2_X1  g504(.A1(G299), .A2(new_n607), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(KEYINPUT41), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT41), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n933), .B1(new_n937), .B2(new_n928), .ZN(new_n938));
  OR2_X1    g513(.A1(new_n938), .A2(KEYINPUT42), .ZN(new_n939));
  NAND2_X1  g514(.A1(G166), .A2(G290), .ZN(new_n940));
  NAND2_X1  g515(.A1(G303), .A2(new_n814), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(new_n941), .A3(G288), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(G288), .B1(new_n940), .B2(new_n941), .ZN(new_n944));
  OAI21_X1  g519(.A(G305), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n940), .A2(new_n941), .ZN(new_n946));
  INV_X1    g521(.A(G288), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n948), .A2(new_n800), .A3(new_n942), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n945), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n938), .A2(KEYINPUT42), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n939), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n950), .B1(new_n939), .B2(new_n951), .ZN(new_n953));
  OAI21_X1  g528(.A(G868), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n873), .A2(new_n611), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(G295));
  NAND2_X1  g531(.A1(new_n954), .A2(new_n955), .ZN(G331));
  NAND2_X1  g532(.A1(G63), .A2(G651), .ZN(new_n958));
  INV_X1    g533(.A(G89), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n958), .B1(new_n513), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n542), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n961), .A2(G301), .A3(new_n534), .A4(new_n532), .ZN(new_n962));
  NAND2_X1  g537(.A1(G286), .A2(G171), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n877), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT103), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n874), .A2(new_n962), .A3(new_n963), .A4(new_n876), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n964), .A2(new_n877), .A3(KEYINPUT103), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n937), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT102), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n965), .A2(new_n972), .A3(new_n967), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n964), .A2(new_n877), .A3(KEYINPUT102), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n931), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n949), .B(new_n945), .C1(new_n971), .C2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n970), .A2(new_n932), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT104), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n934), .A2(new_n936), .A3(new_n974), .A4(new_n973), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n970), .A2(KEYINPUT104), .A3(new_n932), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n979), .A2(new_n950), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n976), .A2(new_n923), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT43), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n923), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT104), .B1(new_n970), .B2(new_n932), .ZN(new_n986));
  AOI211_X1 g561(.A(new_n978), .B(new_n931), .C1(new_n968), .C2(new_n969), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n950), .B1(new_n988), .B2(new_n980), .ZN(new_n989));
  OR2_X1    g564(.A1(new_n985), .A2(new_n989), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n984), .B(KEYINPUT44), .C1(new_n990), .C2(KEYINPUT43), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT105), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT43), .B1(new_n985), .B2(new_n989), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT43), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n976), .A2(new_n982), .A3(new_n994), .A4(new_n923), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT44), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n992), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AOI211_X1 g573(.A(KEYINPUT105), .B(KEYINPUT44), .C1(new_n993), .C2(new_n995), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n991), .B1(new_n998), .B2(new_n999), .ZN(G397));
  XNOR2_X1  g575(.A(KEYINPUT106), .B(G1384), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n501), .A2(new_n504), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1001), .B1(new_n1002), .B2(new_n913), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n462), .A2(new_n467), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(G2105), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT66), .B1(new_n476), .B2(new_n460), .ZN(new_n1006));
  AOI211_X1 g581(.A(new_n469), .B(G2105), .C1(new_n475), .C2(new_n470), .ZN(new_n1007));
  OAI211_X1 g582(.A(G40), .B(new_n1005), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n1003), .A2(new_n1008), .A3(KEYINPUT45), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n757), .B(G2067), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n1010), .B(KEYINPUT107), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1996), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n718), .B(new_n1013), .ZN(new_n1014));
  XOR2_X1   g589(.A(new_n823), .B(new_n826), .Z(new_n1015));
  XNOR2_X1  g590(.A(new_n1015), .B(KEYINPUT108), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1012), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(G290), .B(G1986), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1009), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1001), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n914), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT45), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT109), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT109), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1003), .A2(new_n1025), .A3(KEYINPUT45), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1028), .A2(G2078), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1008), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1027), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT121), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G1384), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n914), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1008), .B1(new_n1035), .B2(new_n1023), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1025), .B1(new_n1003), .B2(KEYINPUT45), .ZN(new_n1037));
  NOR4_X1   g612(.A1(G164), .A2(KEYINPUT109), .A3(new_n1023), .A4(new_n1001), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1036), .B(new_n699), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n1028), .ZN(new_n1040));
  INV_X1    g615(.A(G40), .ZN(new_n1041));
  AOI211_X1 g616(.A(new_n1041), .B(new_n468), .C1(new_n474), .C2(new_n477), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT50), .ZN(new_n1043));
  NOR3_X1   g618(.A1(G164), .A2(new_n1043), .A3(G1384), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT50), .B1(new_n914), .B2(new_n1034), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1042), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n737), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1027), .A2(KEYINPUT121), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1033), .A2(new_n1040), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(G171), .ZN(new_n1050));
  AOI22_X1  g625(.A1(new_n1039), .A2(new_n1028), .B1(new_n737), .B2(new_n1046), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n914), .A2(KEYINPUT45), .A3(new_n1034), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1036), .A2(new_n1029), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(G301), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1020), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1051), .A2(G301), .A3(new_n1053), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT122), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1049), .A2(G171), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT122), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1051), .A2(new_n1059), .A3(G301), .A4(new_n1053), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1057), .A2(new_n1058), .A3(KEYINPUT54), .A4(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT51), .ZN(new_n1062));
  XNOR2_X1  g637(.A(KEYINPUT111), .B(G8), .ZN(new_n1063));
  NAND2_X1  g638(.A1(G286), .A2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1043), .B1(G164), .B2(G1384), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n914), .A2(KEYINPUT50), .A3(new_n1034), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1008), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1023), .B1(G164), .B2(G1384), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1068), .A2(new_n1042), .A3(new_n1052), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n732), .A2(new_n1067), .B1(new_n1069), .B2(new_n764), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1063), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1062), .B(new_n1064), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G8), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1069), .A2(new_n764), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n732), .B(new_n1042), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1073), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1064), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT51), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n1077), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1072), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  XNOR2_X1  g658(.A(KEYINPUT110), .B(KEYINPUT55), .ZN(new_n1084));
  NAND3_X1  g659(.A1(G303), .A2(G8), .A3(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(G166), .A2(new_n1073), .ZN(new_n1086));
  AND2_X1   g661(.A1(KEYINPUT110), .A2(KEYINPUT55), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1036), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1090));
  INV_X1    g665(.A(G2090), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1090), .A2(new_n796), .B1(new_n1091), .B2(new_n1067), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1089), .B1(new_n1092), .B2(new_n1071), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1067), .A2(new_n1091), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(G1971), .B1(new_n1027), .B2(new_n1036), .ZN(new_n1096));
  OAI211_X1 g671(.A(G8), .B(new_n1088), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(G1384), .B1(new_n1002), .B2(new_n913), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1042), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G1976), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT52), .B1(G288), .B2(new_n1100), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n577), .A2(G1976), .A3(new_n578), .A4(new_n579), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1099), .A2(new_n1101), .A3(new_n1063), .A4(new_n1102), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1063), .B(new_n1102), .C1(new_n1035), .C2(new_n1008), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT52), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT112), .ZN(new_n1107));
  NAND2_X1  g682(.A1(G305), .A2(G1981), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n506), .B1(new_n585), .B2(new_n586), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1109), .B1(new_n519), .B2(G86), .ZN(new_n1110));
  INV_X1    g685(.A(G1981), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1110), .A2(new_n1111), .A3(new_n582), .A4(new_n590), .ZN(new_n1112));
  AND4_X1   g687(.A1(new_n1107), .A2(new_n1108), .A3(new_n1112), .A4(KEYINPUT49), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT49), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1114), .A2(KEYINPUT112), .ZN(new_n1115));
  AOI22_X1  g690(.A1(G305), .A2(G1981), .B1(KEYINPUT112), .B2(new_n1114), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1115), .B1(new_n1116), .B2(new_n1112), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1071), .B1(new_n1042), .B2(new_n1098), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1106), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1093), .A2(new_n1097), .A3(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1055), .A2(new_n1061), .A3(new_n1083), .A4(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT117), .ZN(new_n1123));
  INV_X1    g698(.A(G1348), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n1035), .A2(new_n1008), .A3(G2067), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT116), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n1046), .A2(new_n1124), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1098), .A2(G40), .A3(G160), .A4(new_n745), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT116), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1123), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1042), .A2(new_n1126), .A3(new_n745), .A4(new_n1098), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1129), .B(new_n1131), .C1(new_n1067), .C2(G1348), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1132), .A2(KEYINPUT117), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT60), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1134), .A2(KEYINPUT120), .A3(new_n607), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT60), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1132), .A2(KEYINPUT117), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1046), .A2(new_n1124), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1140), .A2(new_n1123), .A3(new_n1129), .A4(new_n1131), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1137), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT120), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n608), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AOI211_X1 g719(.A(KEYINPUT120), .B(new_n1137), .C1(new_n1139), .C2(new_n1141), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1135), .B(new_n1138), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(KEYINPUT56), .B(G2072), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1036), .B(new_n1147), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT114), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  OR2_X1    g725(.A1(new_n1067), .A2(G1956), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1027), .A2(KEYINPUT114), .A3(new_n1036), .A4(new_n1147), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT57), .ZN(new_n1153));
  XNOR2_X1  g728(.A(G299), .B(new_n1153), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .A4(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT115), .ZN(new_n1156));
  OR2_X1    g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1159));
  XNOR2_X1  g734(.A(G299), .B(KEYINPUT57), .ZN(new_n1160));
  AOI21_X1  g735(.A(KEYINPUT61), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1157), .A2(new_n1158), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT118), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1154), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1160), .A2(KEYINPUT118), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1159), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(new_n1155), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(KEYINPUT61), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1162), .A2(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g745(.A(KEYINPUT119), .B(G1996), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1027), .A2(new_n1036), .A3(new_n1171), .ZN(new_n1172));
  XOR2_X1   g747(.A(KEYINPUT58), .B(G1341), .Z(new_n1173));
  NAND2_X1  g748(.A1(new_n1099), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n617), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  XOR2_X1   g750(.A(new_n1175), .B(KEYINPUT59), .Z(new_n1176));
  NAND3_X1  g751(.A1(new_n1146), .A2(new_n1170), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1136), .A2(new_n608), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(new_n1167), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1179), .A2(new_n1158), .A3(new_n1157), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1122), .B1(new_n1177), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT62), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1082), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT123), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1183), .A2(new_n1184), .A3(new_n1121), .A4(new_n1054), .ZN(new_n1185));
  OAI211_X1 g760(.A(new_n1080), .B(KEYINPUT51), .C1(new_n1077), .C2(new_n1076), .ZN(new_n1186));
  AOI21_X1  g761(.A(KEYINPUT62), .B1(new_n1186), .B2(new_n1072), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1054), .A2(new_n1093), .A3(new_n1097), .A4(new_n1120), .ZN(new_n1188));
  OAI21_X1  g763(.A(KEYINPUT123), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  OR3_X1    g764(.A1(new_n1082), .A2(KEYINPUT124), .A3(new_n1182), .ZN(new_n1190));
  OAI21_X1  g765(.A(KEYINPUT124), .B1(new_n1082), .B2(new_n1182), .ZN(new_n1191));
  NAND4_X1  g766(.A1(new_n1185), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1070), .A2(G286), .A3(new_n1071), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1090), .A2(new_n796), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1073), .B1(new_n1194), .B2(new_n1094), .ZN(new_n1195));
  OAI211_X1 g770(.A(new_n1120), .B(new_n1193), .C1(new_n1195), .C2(new_n1088), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1196), .A2(KEYINPUT63), .ZN(new_n1197));
  XOR2_X1   g772(.A(new_n1112), .B(KEYINPUT113), .Z(new_n1198));
  NAND2_X1  g773(.A1(new_n1198), .A2(new_n1119), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1201));
  NOR4_X1   g776(.A1(new_n1070), .A2(KEYINPUT63), .A3(G286), .A4(new_n1071), .ZN(new_n1202));
  AOI22_X1  g777(.A1(new_n1093), .A2(new_n1202), .B1(new_n1195), .B2(new_n1088), .ZN(new_n1203));
  OAI22_X1  g778(.A1(new_n1203), .A2(new_n1106), .B1(G288), .B2(new_n1104), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1200), .B1(new_n1201), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1192), .A2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1019), .B1(new_n1181), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT47), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1009), .B1(new_n1011), .B2(new_n718), .ZN(new_n1209));
  AND2_X1   g784(.A1(new_n1009), .A2(new_n1013), .ZN(new_n1210));
  OR2_X1    g785(.A1(new_n1210), .A2(KEYINPUT46), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1210), .A2(KEYINPUT46), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1209), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1213), .A2(KEYINPUT125), .ZN(new_n1214));
  INV_X1    g789(.A(new_n1214), .ZN(new_n1215));
  NOR2_X1   g790(.A1(new_n1213), .A2(KEYINPUT125), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n1208), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g792(.A(new_n1216), .ZN(new_n1218));
  NAND3_X1  g793(.A1(new_n1218), .A2(KEYINPUT47), .A3(new_n1214), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n824), .A2(new_n826), .ZN(new_n1221));
  OAI22_X1  g796(.A1(new_n1220), .A2(new_n1221), .B1(G2067), .B2(new_n757), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1017), .A2(new_n1009), .ZN(new_n1223));
  NAND3_X1  g798(.A1(new_n1009), .A2(new_n816), .A3(new_n814), .ZN(new_n1224));
  XNOR2_X1  g799(.A(new_n1224), .B(KEYINPUT48), .ZN(new_n1225));
  AOI22_X1  g800(.A1(new_n1222), .A2(new_n1009), .B1(new_n1223), .B2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g801(.A1(new_n1217), .A2(new_n1219), .A3(new_n1226), .ZN(new_n1227));
  INV_X1    g802(.A(KEYINPUT126), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NAND4_X1  g804(.A1(new_n1217), .A2(new_n1219), .A3(KEYINPUT126), .A4(new_n1226), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n1207), .A2(new_n1231), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g807(.A1(new_n658), .A2(G319), .A3(new_n673), .ZN(new_n1234));
  INV_X1    g808(.A(KEYINPUT127), .ZN(new_n1235));
  XNOR2_X1  g809(.A(new_n1234), .B(new_n1235), .ZN(new_n1236));
  AND4_X1   g810(.A1(new_n694), .A2(new_n1236), .A3(new_n926), .A4(new_n996), .ZN(G308));
  NAND4_X1  g811(.A1(new_n694), .A2(new_n1236), .A3(new_n926), .A4(new_n996), .ZN(G225));
endmodule


