//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 0 0 0 1 0 1 1 0 0 1 1 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n814, new_n816, new_n817, new_n819, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937;
  INV_X1    g000(.A(KEYINPUT87), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT86), .ZN(new_n204));
  INV_X1    g003(.A(G1gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AND2_X1   g005(.A1(new_n205), .A2(KEYINPUT16), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n206), .B1(new_n204), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G8gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n208), .A2(G8gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n202), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n208), .A2(G8gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n213), .A2(KEYINPUT87), .A3(new_n209), .ZN(new_n214));
  XOR2_X1   g013(.A(KEYINPUT85), .B(KEYINPUT17), .Z(new_n215));
  INV_X1    g014(.A(G36gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT14), .ZN(new_n217));
  INV_X1    g016(.A(G29gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n217), .B(new_n218), .ZN(new_n219));
  XOR2_X1   g018(.A(G43gat), .B(G50gat), .Z(new_n220));
  INV_X1    g019(.A(KEYINPUT15), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT83), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT14), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n223), .B1(new_n224), .B2(G36gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n219), .A2(new_n222), .A3(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n220), .A2(new_n221), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT84), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n226), .A2(new_n227), .ZN(new_n231));
  NOR3_X1   g030(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n226), .A2(new_n227), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT84), .B1(new_n233), .B2(new_n228), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n215), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n227), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n226), .B(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT17), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n212), .A2(new_n214), .A3(new_n235), .A4(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G229gat), .A2(G233gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n210), .A2(new_n211), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n232), .A2(new_n234), .ZN(new_n242));
  NOR3_X1   g041(.A1(new_n241), .A2(new_n242), .A3(KEYINPUT88), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT88), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n213), .A2(new_n209), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n237), .A2(KEYINPUT84), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n230), .B1(new_n229), .B2(new_n231), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n244), .B1(new_n245), .B2(new_n248), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n239), .B(new_n240), .C1(new_n243), .C2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT18), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  OAI22_X1  g051(.A1(new_n243), .A2(new_n249), .B1(new_n245), .B2(new_n248), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n240), .B(KEYINPUT13), .Z(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(KEYINPUT88), .B1(new_n241), .B2(new_n242), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n245), .A2(new_n248), .A3(new_n244), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n258), .A2(KEYINPUT18), .A3(new_n240), .A4(new_n239), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n252), .A2(new_n255), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT82), .ZN(new_n261));
  XNOR2_X1  g060(.A(G113gat), .B(G141gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(G197gat), .ZN(new_n263));
  XOR2_X1   g062(.A(KEYINPUT11), .B(G169gat), .Z(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n265), .B(KEYINPUT12), .Z(new_n266));
  NAND2_X1  g065(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n266), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n260), .A2(KEYINPUT82), .A3(new_n268), .ZN(new_n269));
  AND2_X1   g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G78gat), .B(G106gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT31), .B(G50gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT3), .ZN(new_n276));
  XNOR2_X1  g075(.A(G197gat), .B(G204gat), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT22), .ZN(new_n278));
  INV_X1    g077(.A(G211gat), .ZN(new_n279));
  INV_X1    g078(.A(G218gat), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  XOR2_X1   g081(.A(G211gat), .B(G218gat), .Z(new_n283));
  OR2_X1    g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n283), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n284), .A2(KEYINPUT67), .A3(new_n285), .ZN(new_n286));
  OR2_X1    g085(.A1(new_n285), .A2(KEYINPUT67), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n276), .B1(new_n288), .B2(KEYINPUT29), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT69), .ZN(new_n290));
  AND2_X1   g089(.A1(G141gat), .A2(G148gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(G141gat), .A2(G148gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G155gat), .B(G162gat), .ZN(new_n294));
  INV_X1    g093(.A(G155gat), .ZN(new_n295));
  INV_X1    g094(.A(G162gat), .ZN(new_n296));
  OAI21_X1  g095(.A(KEYINPUT2), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n293), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n294), .B1(new_n293), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n290), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n292), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT2), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT68), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT68), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT2), .ZN(new_n306));
  NAND2_X1  g105(.A1(G141gat), .A2(G148gat), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n302), .A2(new_n304), .A3(new_n306), .A4(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n294), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n293), .A2(new_n294), .A3(new_n297), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n310), .A2(KEYINPUT69), .A3(new_n311), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n301), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n289), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G228gat), .ZN(new_n315));
  INV_X1    g114(.A(G233gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT29), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n310), .A2(new_n311), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n318), .B1(new_n319), .B2(KEYINPUT3), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n288), .A2(KEYINPUT75), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n288), .A2(new_n320), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT75), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n314), .A2(new_n317), .A3(new_n321), .A4(new_n324), .ZN(new_n325));
  XOR2_X1   g124(.A(KEYINPUT76), .B(G22gat), .Z(new_n326));
  INV_X1    g125(.A(new_n322), .ZN(new_n327));
  INV_X1    g126(.A(new_n319), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n284), .A2(new_n285), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n318), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n328), .B1(new_n330), .B2(new_n276), .ZN(new_n331));
  OAI22_X1  g130(.A1(new_n327), .A2(new_n331), .B1(new_n315), .B2(new_n316), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n325), .A2(new_n326), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n326), .B1(new_n325), .B2(new_n332), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n275), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n325), .A2(new_n332), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(G22gat), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n325), .A2(KEYINPUT77), .A3(new_n326), .A4(new_n332), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n338), .A3(new_n274), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n333), .A2(KEYINPUT77), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n335), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(G169gat), .A2(G176gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(G169gat), .A2(G176gat), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT26), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AOI22_X1  g144(.A1(new_n345), .A2(KEYINPUT65), .B1(new_n344), .B2(new_n343), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT65), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n347), .B(new_n342), .C1(new_n343), .C2(new_n344), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT27), .B(G183gat), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT28), .ZN(new_n351));
  INV_X1    g150(.A(G190gat), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(G183gat), .A2(G190gat), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n350), .A2(new_n352), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n355), .B1(new_n356), .B2(KEYINPUT28), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n349), .A2(new_n353), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT64), .ZN(new_n359));
  OAI21_X1  g158(.A(KEYINPUT25), .B1(new_n342), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n360), .B1(new_n359), .B2(new_n342), .ZN(new_n361));
  AND2_X1   g160(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(G190gat), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n363), .B1(new_n365), .B2(new_n355), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n343), .A2(KEYINPUT23), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT23), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n368), .B1(G169gat), .B2(G176gat), .ZN(new_n369));
  AND2_X1   g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n361), .A2(new_n366), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT25), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n367), .A2(new_n369), .A3(new_n342), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n354), .A2(new_n364), .B1(new_n362), .B2(G190gat), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n358), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G113gat), .B(G120gat), .ZN(new_n378));
  OR2_X1    g177(.A1(KEYINPUT66), .A2(KEYINPUT1), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G127gat), .B(G134gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n381), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n383), .B1(new_n378), .B2(new_n379), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n377), .A2(new_n385), .ZN(new_n386));
  AND2_X1   g185(.A1(new_n382), .A2(new_n384), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n358), .A2(new_n376), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(G227gat), .A2(G233gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT34), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT34), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n386), .A2(new_n393), .A3(new_n390), .A4(new_n388), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  XOR2_X1   g194(.A(G15gat), .B(G43gat), .Z(new_n396));
  XNOR2_X1  g195(.A(G71gat), .B(G99gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n396), .B(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n389), .A2(new_n391), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT33), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n395), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n400), .A2(KEYINPUT32), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n390), .B1(new_n386), .B2(new_n388), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n398), .B1(new_n406), .B2(KEYINPUT33), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(new_n392), .A3(new_n394), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n403), .A2(new_n405), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n405), .B1(new_n403), .B2(new_n408), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n341), .A2(new_n411), .A3(KEYINPUT81), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT35), .ZN(new_n413));
  AND2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT30), .ZN(new_n415));
  INV_X1    g214(.A(new_n288), .ZN(new_n416));
  NAND2_X1  g215(.A1(G226gat), .A2(G233gat), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n418), .B1(new_n377), .B2(new_n318), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n417), .B1(new_n358), .B2(new_n376), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n416), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n420), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT29), .B1(new_n358), .B2(new_n376), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n422), .B(new_n288), .C1(new_n418), .C2(new_n423), .ZN(new_n424));
  AND2_X1   g223(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(G8gat), .B(G36gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(G64gat), .B(G92gat), .ZN(new_n427));
  XOR2_X1   g226(.A(new_n426), .B(new_n427), .Z(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n415), .B1(new_n425), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n425), .A2(new_n429), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n429), .B1(new_n421), .B2(new_n424), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT30), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n430), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT5), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n387), .A2(new_n328), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT4), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(G225gat), .A2(G233gat), .ZN(new_n439));
  XOR2_X1   g238(.A(new_n439), .B(KEYINPUT72), .Z(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n387), .A2(KEYINPUT4), .A3(new_n328), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n438), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n301), .A2(KEYINPUT3), .A3(new_n312), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT70), .B1(new_n319), .B2(KEYINPUT3), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n301), .A2(KEYINPUT70), .A3(new_n312), .A4(KEYINPUT3), .ZN(new_n448));
  AND4_X1   g247(.A1(KEYINPUT71), .A2(new_n447), .A3(new_n448), .A4(new_n385), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n387), .B1(new_n445), .B2(new_n446), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT71), .B1(new_n450), .B2(new_n448), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n435), .B(new_n444), .C1(new_n449), .C2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n447), .A2(new_n448), .A3(new_n385), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT71), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n450), .A2(KEYINPUT71), .A3(new_n448), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n443), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT73), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n301), .A2(new_n312), .A3(new_n385), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n436), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n458), .B1(new_n460), .B2(new_n441), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n436), .A2(new_n459), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n462), .A2(KEYINPUT73), .A3(new_n440), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n461), .A2(KEYINPUT5), .A3(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n452), .B1(new_n457), .B2(new_n464), .ZN(new_n465));
  XOR2_X1   g264(.A(G1gat), .B(G29gat), .Z(new_n466));
  XNOR2_X1  g265(.A(KEYINPUT74), .B(KEYINPUT0), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n466), .B(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G57gat), .B(G85gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n468), .B(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT6), .ZN(new_n472));
  INV_X1    g271(.A(new_n470), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n452), .B(new_n473), .C1(new_n457), .C2(new_n464), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n471), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n465), .A2(KEYINPUT6), .A3(new_n470), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n434), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n477), .A2(new_n341), .A3(new_n411), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n414), .B(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT80), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT38), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT37), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n421), .A2(new_n424), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n483), .B1(new_n421), .B2(new_n424), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n482), .B(new_n429), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n429), .B1(new_n484), .B2(new_n485), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n432), .B1(new_n487), .B2(KEYINPUT38), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n475), .A2(new_n476), .A3(new_n486), .A4(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n341), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT39), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n491), .B1(new_n460), .B2(new_n441), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n438), .A2(new_n442), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n493), .B1(new_n455), .B2(new_n456), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n492), .B1(new_n494), .B2(new_n441), .ZN(new_n495));
  INV_X1    g294(.A(new_n493), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n496), .B1(new_n449), .B2(new_n451), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(new_n491), .A3(new_n440), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n495), .A2(new_n498), .A3(KEYINPUT40), .A4(new_n473), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n499), .A2(new_n434), .A3(new_n471), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n495), .A2(new_n498), .A3(KEYINPUT78), .A4(new_n473), .ZN(new_n501));
  XOR2_X1   g300(.A(KEYINPUT79), .B(KEYINPUT40), .Z(new_n502));
  AND2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT78), .ZN(new_n504));
  INV_X1    g303(.A(new_n495), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n498), .A2(new_n473), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n500), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n481), .B1(new_n490), .B2(new_n508), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n434), .A2(new_n471), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n498), .A2(new_n473), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT78), .B1(new_n511), .B2(new_n495), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n501), .A2(new_n502), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n510), .B(new_n499), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n514), .A2(KEYINPUT80), .A3(new_n341), .A4(new_n489), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n509), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n410), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n403), .A2(new_n408), .A3(new_n405), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n517), .A2(KEYINPUT36), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT36), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n520), .B1(new_n409), .B2(new_n410), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(new_n477), .B2(new_n341), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n516), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n271), .B1(new_n480), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT8), .ZN(new_n527));
  NAND2_X1  g326(.A1(G99gat), .A2(G106gat), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n527), .B1(new_n528), .B2(KEYINPUT96), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n529), .B1(KEYINPUT96), .B2(new_n528), .ZN(new_n530));
  XNOR2_X1  g329(.A(KEYINPUT97), .B(G85gat), .ZN(new_n531));
  INV_X1    g330(.A(G92gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G85gat), .A2(G92gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n530), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G99gat), .B(G106gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n235), .A2(new_n238), .A3(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT41), .ZN(new_n540));
  INV_X1    g339(.A(G232gat), .ZN(new_n541));
  NOR3_X1   g340(.A1(new_n540), .A2(new_n541), .A3(new_n316), .ZN(new_n542));
  INV_X1    g341(.A(new_n538), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n542), .B1(new_n248), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G190gat), .B(G218gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(KEYINPUT98), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n545), .B(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT95), .ZN(new_n549));
  XNOR2_X1  g348(.A(G134gat), .B(G162gat), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n540), .B1(new_n541), .B2(new_n316), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XOR2_X1   g351(.A(KEYINPUT93), .B(KEYINPUT94), .Z(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n554), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n548), .A2(KEYINPUT95), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT99), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n558), .A2(new_n559), .A3(new_n548), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n555), .A2(KEYINPUT99), .A3(new_n557), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT21), .ZN(new_n563));
  INV_X1    g362(.A(G71gat), .ZN(new_n564));
  INV_X1    g363(.A(G78gat), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(KEYINPUT89), .B1(new_n566), .B2(KEYINPUT9), .ZN(new_n567));
  NOR2_X1   g366(.A1(G71gat), .A2(G78gat), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n567), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(G57gat), .B(G64gat), .Z(new_n570));
  OAI21_X1  g369(.A(new_n570), .B1(KEYINPUT9), .B2(new_n566), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n569), .B(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n241), .B1(new_n563), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n563), .ZN(new_n574));
  XOR2_X1   g373(.A(KEYINPUT91), .B(KEYINPUT19), .Z(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n573), .B(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G127gat), .B(G155gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT20), .ZN(new_n579));
  NAND2_X1  g378(.A1(G231gat), .A2(G233gat), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n580), .B(KEYINPUT90), .Z(new_n581));
  XNOR2_X1  g380(.A(new_n579), .B(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G183gat), .B(G211gat), .Z(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT92), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n582), .B(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n577), .B(new_n585), .Z(new_n586));
  NAND2_X1  g385(.A1(new_n562), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G230gat), .A2(G233gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT103), .ZN(new_n589));
  INV_X1    g388(.A(new_n572), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT100), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n536), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT101), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n537), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT100), .B1(new_n537), .B2(new_n593), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n536), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n590), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT10), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n538), .A2(new_n572), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n543), .A2(KEYINPUT10), .A3(new_n590), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n589), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n589), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n603), .B1(new_n597), .B2(new_n599), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G120gat), .B(G148gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(G176gat), .B(G204gat), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n606), .B(new_n607), .Z(new_n608));
  OR3_X1    g407(.A1(new_n605), .A2(KEYINPUT104), .A3(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(KEYINPUT104), .B1(new_n605), .B2(new_n608), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n600), .A2(new_n601), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT102), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n589), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n600), .A2(KEYINPUT102), .A3(new_n601), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n608), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n604), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n611), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n587), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n526), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n475), .A2(new_n476), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(new_n205), .ZN(G1324gat));
  INV_X1    g424(.A(new_n622), .ZN(new_n626));
  XOR2_X1   g425(.A(KEYINPUT16), .B(G8gat), .Z(new_n627));
  NAND3_X1  g426(.A1(new_n626), .A2(new_n434), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT42), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n434), .ZN(new_n631));
  OAI21_X1  g430(.A(G8gat), .B1(new_n622), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n628), .A2(new_n629), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n630), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT105), .ZN(G1325gat));
  AOI21_X1  g434(.A(G15gat), .B1(new_n626), .B2(new_n411), .ZN(new_n636));
  INV_X1    g435(.A(new_n522), .ZN(new_n637));
  OR2_X1    g436(.A1(new_n637), .A2(KEYINPUT106), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(KEYINPUT106), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(G15gat), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n642), .B(KEYINPUT107), .Z(new_n643));
  AOI21_X1  g442(.A(new_n636), .B1(new_n626), .B2(new_n643), .ZN(G1326gat));
  NOR2_X1   g443(.A1(new_n622), .A2(new_n341), .ZN(new_n645));
  XOR2_X1   g444(.A(KEYINPUT43), .B(G22gat), .Z(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(G1327gat));
  NOR3_X1   g446(.A1(new_n562), .A2(new_n586), .A3(new_n620), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT108), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n526), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n623), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n651), .A2(new_n218), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT45), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n271), .A2(new_n586), .A3(new_n620), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n562), .A2(KEYINPUT44), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n525), .A2(KEYINPUT109), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n523), .B1(new_n509), .B2(new_n515), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT109), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n657), .B1(new_n662), .B2(new_n480), .ZN(new_n663));
  INV_X1    g462(.A(new_n562), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n664), .B1(new_n479), .B2(new_n659), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n665), .A2(KEYINPUT44), .ZN(new_n666));
  OAI211_X1 g465(.A(KEYINPUT110), .B(new_n655), .C1(new_n663), .C2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT110), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n660), .B1(new_n516), .B2(new_n524), .ZN(new_n669));
  AOI211_X1 g468(.A(KEYINPUT109), .B(new_n523), .C1(new_n509), .C2(new_n515), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n480), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AOI22_X1  g470(.A1(new_n671), .A2(new_n656), .B1(KEYINPUT44), .B2(new_n665), .ZN(new_n672));
  INV_X1    g471(.A(new_n655), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n668), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  AND3_X1   g473(.A1(new_n667), .A2(new_n674), .A3(new_n652), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n654), .B1(new_n218), .B2(new_n675), .ZN(G1328gat));
  NAND3_X1  g475(.A1(new_n667), .A2(new_n674), .A3(new_n434), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n216), .B1(new_n677), .B2(KEYINPUT111), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n678), .B1(KEYINPUT111), .B2(new_n677), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n650), .A2(G36gat), .A3(new_n631), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT46), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n681), .ZN(G1329gat));
  OAI21_X1  g481(.A(new_n655), .B1(new_n663), .B2(new_n666), .ZN(new_n683));
  OAI21_X1  g482(.A(G43gat), .B1(new_n683), .B2(new_n522), .ZN(new_n684));
  INV_X1    g483(.A(G43gat), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n651), .A2(new_n685), .A3(new_n411), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n684), .A2(KEYINPUT47), .A3(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n667), .A2(new_n674), .A3(new_n641), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(G43gat), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n689), .A2(new_n686), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n687), .B1(new_n690), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g490(.A(new_n341), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n667), .A2(new_n674), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(G50gat), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT48), .ZN(new_n695));
  INV_X1    g494(.A(G50gat), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n695), .B1(new_n650), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT112), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n672), .A2(new_n673), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n696), .B1(new_n702), .B2(new_n692), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n650), .A2(new_n697), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT48), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n700), .A2(new_n701), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n698), .B1(new_n693), .B2(G50gat), .ZN(new_n707));
  OAI21_X1  g506(.A(G50gat), .B1(new_n683), .B2(new_n341), .ZN(new_n708));
  INV_X1    g507(.A(new_n704), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n695), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(KEYINPUT112), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n706), .A2(new_n711), .ZN(G1331gat));
  INV_X1    g511(.A(new_n619), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n713), .B1(new_n610), .B2(new_n609), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n270), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n671), .A2(new_n586), .A3(new_n562), .A4(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n652), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(G57gat), .ZN(G1332gat));
  XOR2_X1   g518(.A(new_n434), .B(KEYINPUT113), .Z(new_n720));
  NOR2_X1   g519(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n722));
  AND2_X1   g521(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n724), .B1(new_n721), .B2(new_n722), .ZN(G1333gat));
  OAI21_X1  g524(.A(G71gat), .B1(new_n716), .B2(new_n640), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n411), .A2(new_n564), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n726), .B1(new_n716), .B2(new_n727), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n728), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g528(.A1(new_n716), .A2(new_n341), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(new_n565), .ZN(G1335gat));
  INV_X1    g530(.A(KEYINPUT51), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n479), .B1(new_n658), .B2(new_n661), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n562), .A2(new_n586), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n271), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n732), .B1(new_n733), .B2(new_n735), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n671), .A2(KEYINPUT51), .A3(new_n271), .A4(new_n734), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n620), .A2(new_n652), .A3(new_n531), .ZN(new_n740));
  INV_X1    g539(.A(new_n586), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n715), .A2(new_n741), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n672), .A2(new_n623), .A3(new_n742), .ZN(new_n743));
  OAI22_X1  g542(.A1(new_n739), .A2(new_n740), .B1(new_n743), .B2(new_n531), .ZN(G1336gat));
  NOR3_X1   g543(.A1(new_n720), .A2(new_n714), .A3(G92gat), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n738), .A2(new_n745), .ZN(new_n746));
  XOR2_X1   g545(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n747));
  NOR3_X1   g546(.A1(new_n672), .A2(new_n720), .A3(new_n742), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n746), .B(new_n747), .C1(new_n748), .C2(new_n532), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n672), .A2(new_n631), .A3(new_n742), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n746), .B1(new_n532), .B2(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n751), .A2(KEYINPUT114), .A3(KEYINPUT52), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT114), .B1(new_n751), .B2(KEYINPUT52), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n749), .B1(new_n753), .B2(new_n754), .ZN(G1337gat));
  INV_X1    g554(.A(G99gat), .ZN(new_n756));
  INV_X1    g555(.A(new_n411), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n714), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n738), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n672), .A2(new_n640), .A3(new_n742), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n759), .B1(new_n756), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT116), .ZN(G1338gat));
  NOR3_X1   g561(.A1(new_n672), .A2(new_n341), .A3(new_n742), .ZN(new_n763));
  INV_X1    g562(.A(G106gat), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n714), .A2(G106gat), .A3(new_n341), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n767), .B1(new_n736), .B2(new_n737), .ZN(new_n768));
  OAI211_X1 g567(.A(KEYINPUT117), .B(KEYINPUT53), .C1(new_n765), .C2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  OAI22_X1  g569(.A1(new_n739), .A2(new_n767), .B1(new_n763), .B2(new_n764), .ZN(new_n771));
  AOI21_X1  g570(.A(KEYINPUT117), .B1(new_n771), .B2(KEYINPUT53), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT118), .ZN(new_n773));
  NOR4_X1   g572(.A1(new_n765), .A2(new_n773), .A3(new_n768), .A4(KEYINPUT53), .ZN(new_n774));
  INV_X1    g573(.A(new_n742), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n692), .B(new_n775), .C1(new_n663), .C2(new_n666), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n768), .B1(G106gat), .B2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT118), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI22_X1  g578(.A1(new_n770), .A2(new_n772), .B1(new_n774), .B2(new_n779), .ZN(G1339gat));
  AND4_X1   g579(.A1(new_n271), .A2(new_n562), .A3(new_n586), .A4(new_n714), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783));
  OAI21_X1  g582(.A(KEYINPUT54), .B1(new_n612), .B2(new_n603), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n784), .B1(new_n615), .B2(new_n614), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT54), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n608), .B1(new_n602), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n783), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n785), .A2(new_n788), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n713), .B1(new_n790), .B2(KEYINPUT55), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n267), .A2(new_n269), .A3(new_n789), .A4(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT119), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n253), .A2(new_n254), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n240), .B1(new_n258), .B2(new_n239), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n265), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n252), .A2(new_n255), .A3(new_n259), .A4(new_n268), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n793), .B1(new_n714), .B2(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n620), .A2(KEYINPUT119), .A3(new_n796), .A4(new_n797), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n792), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n562), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n789), .A2(new_n796), .A3(new_n797), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n560), .A2(new_n561), .A3(new_n791), .A4(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n802), .A2(KEYINPUT120), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n741), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT120), .B1(new_n802), .B2(new_n804), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n782), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n808), .A2(new_n341), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n809), .A2(new_n652), .A3(new_n411), .A4(new_n720), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n810), .A2(new_n271), .ZN(new_n811));
  INV_X1    g610(.A(G113gat), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n811), .B(new_n812), .ZN(G1340gat));
  NAND4_X1  g612(.A1(new_n809), .A2(new_n652), .A3(new_n720), .A4(new_n758), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(G120gat), .ZN(G1341gat));
  NOR2_X1   g614(.A1(new_n810), .A2(new_n741), .ZN(new_n816));
  INV_X1    g615(.A(G127gat), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n816), .B(new_n817), .ZN(G1342gat));
  NOR4_X1   g617(.A1(new_n562), .A2(G134gat), .A3(new_n434), .A4(new_n757), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n809), .A2(new_n652), .A3(new_n819), .ZN(new_n820));
  XOR2_X1   g619(.A(new_n820), .B(KEYINPUT56), .Z(new_n821));
  OAI21_X1  g620(.A(G134gat), .B1(new_n810), .B2(new_n562), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(G1343gat));
  INV_X1    g622(.A(KEYINPUT57), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n808), .A2(new_n824), .A3(new_n692), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT121), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n614), .A2(new_n615), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n826), .B(new_n787), .C1(new_n827), .C2(new_n784), .ZN(new_n828));
  OAI21_X1  g627(.A(KEYINPUT121), .B1(new_n785), .B2(new_n788), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n828), .A2(new_n829), .A3(new_n783), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n267), .A2(new_n830), .A3(new_n269), .A4(new_n791), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n620), .A2(new_n796), .A3(new_n797), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n562), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT122), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT122), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n833), .A2(new_n562), .A3(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n835), .A2(new_n804), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n781), .B1(new_n838), .B2(new_n741), .ZN(new_n839));
  OAI21_X1  g638(.A(KEYINPUT57), .B1(new_n839), .B2(new_n341), .ZN(new_n840));
  INV_X1    g639(.A(new_n720), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n841), .A2(new_n637), .A3(new_n623), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n825), .A2(new_n840), .A3(new_n270), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(G141gat), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n808), .A2(new_n692), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n641), .A2(new_n623), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n271), .A2(G141gat), .ZN(new_n847));
  XOR2_X1   g646(.A(new_n847), .B(KEYINPUT123), .Z(new_n848));
  NAND4_X1  g647(.A1(new_n845), .A2(new_n720), .A3(new_n846), .A4(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n844), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(KEYINPUT58), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT58), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n844), .A2(new_n852), .A3(new_n849), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(G1344gat));
  NAND2_X1  g653(.A1(new_n845), .A2(new_n846), .ZN(new_n855));
  OR4_X1    g654(.A1(G148gat), .A2(new_n855), .A3(new_n714), .A4(new_n841), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n825), .A2(new_n840), .A3(new_n842), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n857), .A2(new_n714), .ZN(new_n858));
  INV_X1    g657(.A(G148gat), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n858), .A2(KEYINPUT59), .A3(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n808), .A2(new_n692), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(KEYINPUT57), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT124), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n781), .B(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n586), .B1(new_n834), .B2(new_n804), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n824), .B(new_n692), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n863), .A2(new_n620), .A3(new_n842), .A4(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n861), .B1(new_n868), .B2(G148gat), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n856), .B1(new_n860), .B2(new_n869), .ZN(G1345gat));
  NAND4_X1  g669(.A1(new_n825), .A2(new_n840), .A3(new_n586), .A4(new_n842), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(G155gat), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n741), .A2(G155gat), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n845), .A2(new_n720), .A3(new_n846), .A4(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(KEYINPUT125), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT125), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n872), .A2(new_n877), .A3(new_n874), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n878), .ZN(G1346gat));
  OAI21_X1  g678(.A(G162gat), .B1(new_n857), .B2(new_n562), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n664), .A2(new_n296), .A3(new_n631), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n880), .B1(new_n855), .B2(new_n881), .ZN(G1347gat));
  AND2_X1   g681(.A1(new_n808), .A2(new_n623), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n720), .A2(new_n692), .A3(new_n757), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(G169gat), .B1(new_n885), .B2(new_n270), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n623), .A2(new_n434), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n887), .A2(new_n757), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n809), .A2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(G169gat), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n889), .A2(new_n890), .A3(new_n271), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n886), .A2(new_n891), .ZN(G1348gat));
  AOI21_X1  g691(.A(G176gat), .B1(new_n885), .B2(new_n620), .ZN(new_n893));
  INV_X1    g692(.A(G176gat), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n889), .A2(new_n894), .A3(new_n714), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n893), .A2(new_n895), .ZN(G1349gat));
  NAND3_X1  g695(.A1(new_n809), .A2(new_n586), .A3(new_n888), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(G183gat), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT60), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n899), .A2(KEYINPUT126), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n883), .A2(new_n350), .A3(new_n586), .A4(new_n884), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n898), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n900), .B1(new_n898), .B2(new_n901), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n902), .A2(new_n903), .ZN(G1350gat));
  NAND3_X1  g703(.A1(new_n885), .A2(new_n352), .A3(new_n664), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n809), .A2(new_n664), .A3(new_n888), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT61), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n906), .A2(new_n907), .A3(G190gat), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n906), .B2(G190gat), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n905), .B1(new_n908), .B2(new_n909), .ZN(G1351gat));
  NOR3_X1   g709(.A1(new_n641), .A2(new_n341), .A3(new_n720), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n883), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(G197gat), .B1(new_n912), .B2(new_n270), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n863), .A2(new_n867), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n641), .A2(new_n887), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n270), .A2(G197gat), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(G1352gat));
  NAND3_X1  g717(.A1(new_n914), .A2(new_n620), .A3(new_n915), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(G204gat), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n714), .A2(G204gat), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n883), .A2(new_n911), .A3(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n922), .B(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n920), .A2(new_n924), .ZN(G1353gat));
  NAND4_X1  g724(.A1(new_n863), .A2(new_n586), .A3(new_n867), .A4(new_n915), .ZN(new_n926));
  OAI21_X1  g725(.A(G211gat), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n929), .A2(KEYINPUT127), .A3(KEYINPUT63), .ZN(new_n930));
  NAND2_X1  g729(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n926), .A2(new_n928), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n912), .A2(new_n279), .A3(new_n586), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n930), .A2(new_n932), .A3(new_n933), .ZN(G1354gat));
  NAND3_X1  g733(.A1(new_n914), .A2(new_n664), .A3(new_n915), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(G218gat), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n912), .A2(new_n280), .A3(new_n664), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1355gat));
endmodule


