//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 0 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 1 1 1 1 1 0 1 0 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT65), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT0), .Z(new_n213));
  AOI22_X1  g0013(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G58), .ZN(new_n215));
  INV_X1    g0015(.A(G232), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n210), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(G50), .B1(G58), .B2(G68), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT66), .Z(new_n229));
  AOI211_X1 g0029(.A(new_n213), .B(new_n224), .C1(new_n227), .C2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  INV_X1    g0045(.A(KEYINPUT71), .ZN(new_n246));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n225), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  NOR2_X1   g0049(.A1(G20), .A2(G33), .ZN(new_n250));
  AOI22_X1  g0050(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n250), .ZN(new_n251));
  OR3_X1    g0051(.A1(new_n215), .A2(KEYINPUT68), .A3(KEYINPUT8), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n215), .A2(KEYINPUT8), .ZN(new_n253));
  AOI21_X1  g0053(.A(KEYINPUT68), .B1(new_n215), .B2(KEYINPUT8), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n226), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n249), .B1(new_n251), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G13), .A3(G20), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G50), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n249), .B1(G1), .B2(new_n226), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n264), .B1(new_n265), .B2(new_n263), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n259), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G169), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n225), .B1(G33), .B2(G41), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT3), .B(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G1698), .ZN(new_n271));
  XOR2_X1   g0071(.A(KEYINPUT67), .B(G223), .Z(new_n272));
  INV_X1    g0072(.A(G77), .ZN(new_n273));
  OAI22_X1  g0073(.A1(new_n271), .A2(new_n272), .B1(new_n273), .B2(new_n270), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  AND3_X1   g0075(.A1(new_n270), .A2(G222), .A3(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n269), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G41), .ZN(new_n278));
  INV_X1    g0078(.A(G45), .ZN(new_n279));
  AOI21_X1  g0079(.A(G1), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G274), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n269), .A2(new_n280), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n282), .B1(new_n283), .B2(G226), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n277), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n267), .B1(new_n268), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n285), .ZN(new_n287));
  INV_X1    g0087(.A(G179), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  AOI22_X1  g0090(.A1(KEYINPUT9), .A2(new_n267), .B1(new_n287), .B2(G190), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G200), .ZN(new_n293));
  OAI22_X1  g0093(.A1(new_n267), .A2(KEYINPUT9), .B1(new_n287), .B2(new_n293), .ZN(new_n294));
  NOR3_X1   g0094(.A1(new_n292), .A2(new_n294), .A3(KEYINPUT10), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT10), .ZN(new_n296));
  INV_X1    g0096(.A(new_n294), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n296), .B1(new_n297), .B2(new_n291), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n290), .B1(new_n295), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n270), .A2(G232), .A3(new_n275), .ZN(new_n300));
  XOR2_X1   g0100(.A(KEYINPUT69), .B(G107), .Z(new_n301));
  OAI221_X1 g0101(.A(new_n300), .B1(new_n270), .B2(new_n301), .C1(new_n271), .C2(new_n218), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n269), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n283), .A2(G244), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n281), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(KEYINPUT70), .B1(new_n303), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n303), .A2(KEYINPUT70), .A3(new_n306), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n308), .A2(G200), .A3(new_n309), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n303), .A2(KEYINPUT70), .A3(new_n306), .ZN(new_n311));
  OAI21_X1  g0111(.A(G190), .B1(new_n311), .B2(new_n307), .ZN(new_n312));
  AND2_X1   g0112(.A1(new_n215), .A2(KEYINPUT8), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n313), .A2(new_n253), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n315), .A2(new_n250), .B1(G20), .B2(G77), .ZN(new_n316));
  XOR2_X1   g0116(.A(KEYINPUT15), .B(G87), .Z(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n257), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n249), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n262), .A2(new_n273), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(new_n265), .B2(new_n273), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n310), .A2(new_n312), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n308), .A2(new_n268), .A3(new_n309), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n288), .B1(new_n311), .B2(new_n307), .ZN(new_n325));
  INV_X1    g0125(.A(new_n322), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n246), .B1(new_n299), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n290), .ZN(new_n330));
  OAI21_X1  g0130(.A(KEYINPUT10), .B1(new_n292), .B2(new_n294), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n297), .A2(new_n291), .A3(new_n296), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n333), .A2(KEYINPUT71), .A3(new_n323), .A4(new_n327), .ZN(new_n334));
  INV_X1    g0134(.A(G33), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT3), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT3), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G33), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n336), .A2(new_n338), .A3(G226), .A4(G1698), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n336), .A2(new_n338), .A3(G223), .A4(new_n275), .ZN(new_n340));
  NAND2_X1  g0140(.A1(G33), .A2(G87), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n269), .ZN(new_n343));
  NAND2_X1  g0143(.A1(G33), .A2(G41), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n344), .A2(G1), .A3(G13), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n260), .B1(G41), .B2(G45), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(G232), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n281), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n343), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT77), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n348), .B1(new_n342), .B2(new_n269), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT77), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n351), .A2(new_n293), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT79), .ZN(new_n356));
  OR2_X1    g0156(.A1(KEYINPUT78), .A2(G190), .ZN(new_n357));
  NAND2_X1  g0157(.A1(KEYINPUT78), .A2(G190), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n356), .B1(new_n352), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n352), .A2(new_n356), .A3(new_n359), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n355), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT7), .ZN(new_n364));
  NOR3_X1   g0164(.A1(new_n270), .A2(new_n364), .A3(G20), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n336), .A2(new_n338), .ZN(new_n366));
  AOI21_X1  g0166(.A(KEYINPUT7), .B1(new_n366), .B2(new_n226), .ZN(new_n367));
  OAI21_X1  g0167(.A(G68), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n215), .A2(new_n217), .ZN(new_n369));
  OAI21_X1  g0169(.A(G20), .B1(new_n369), .B2(new_n203), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n250), .A2(G159), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n368), .A2(KEYINPUT16), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT16), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n364), .B1(new_n270), .B2(G20), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n366), .A2(KEYINPUT7), .A3(new_n226), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n217), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n375), .B1(new_n378), .B2(new_n372), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n374), .A2(new_n379), .A3(new_n248), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n265), .A2(new_n255), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT76), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n252), .B(new_n261), .C1(new_n253), .C2(new_n254), .ZN(new_n383));
  AND3_X1   g0183(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n382), .B1(new_n381), .B2(new_n383), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n380), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g0187(.A(KEYINPUT80), .B(KEYINPUT17), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n363), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n380), .A2(new_n386), .ZN(new_n390));
  INV_X1    g0190(.A(new_n362), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n391), .A2(new_n360), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n390), .B1(new_n355), .B2(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(KEYINPUT80), .A2(KEYINPUT17), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n389), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT18), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n351), .A2(new_n268), .A3(new_n354), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n350), .A2(G179), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n396), .B1(new_n387), .B2(new_n400), .ZN(new_n401));
  AOI211_X1 g0201(.A(KEYINPUT77), .B(new_n348), .C1(new_n269), .C2(new_n342), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n353), .B1(new_n343), .B2(new_n349), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n398), .B1(new_n404), .B2(new_n268), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n405), .A2(KEYINPUT18), .A3(new_n390), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n401), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n395), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n329), .A2(new_n334), .A3(new_n409), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n257), .A2(G77), .B1(G20), .B2(new_n217), .ZN(new_n411));
  INV_X1    g0211(.A(new_n250), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n411), .B1(new_n263), .B2(new_n412), .ZN(new_n413));
  XOR2_X1   g0213(.A(KEYINPUT74), .B(KEYINPUT11), .Z(new_n414));
  AND3_X1   g0214(.A1(new_n413), .A2(new_n248), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n414), .B1(new_n413), .B2(new_n248), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n262), .A2(KEYINPUT12), .A3(new_n217), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT12), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n261), .B2(G68), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n417), .B(new_n419), .C1(new_n265), .C2(new_n217), .ZN(new_n420));
  NOR3_X1   g0220(.A1(new_n415), .A2(new_n416), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n336), .A2(new_n338), .A3(G232), .A4(G1698), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n336), .A2(new_n338), .A3(G226), .A4(new_n275), .ZN(new_n424));
  NAND2_X1  g0224(.A1(G33), .A2(G97), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n269), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n345), .A2(G238), .A3(new_n346), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n281), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT13), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n429), .B1(new_n426), .B2(new_n269), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT13), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n432), .A2(KEYINPUT72), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT72), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n433), .A2(new_n437), .A3(new_n434), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n436), .A2(G169), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT14), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT14), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n436), .A2(new_n441), .A3(G169), .A4(new_n438), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT73), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n443), .B1(new_n433), .B2(new_n434), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n432), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n431), .A2(new_n443), .A3(KEYINPUT13), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(G179), .ZN(new_n448));
  AND4_X1   g0248(.A1(KEYINPUT75), .A2(new_n440), .A3(new_n442), .A4(new_n448), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n439), .A2(KEYINPUT14), .B1(new_n447), .B2(G179), .ZN(new_n450));
  AOI21_X1  g0250(.A(KEYINPUT75), .B1(new_n450), .B2(new_n442), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n422), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n447), .A2(G190), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n436), .A2(G200), .A3(new_n438), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n453), .A2(new_n454), .A3(new_n421), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  OR2_X1    g0256(.A1(new_n410), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n337), .A2(G33), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n335), .A2(KEYINPUT3), .ZN(new_n459));
  OAI21_X1  g0259(.A(G303), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n336), .A2(new_n338), .A3(G257), .A4(new_n275), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n336), .A2(new_n338), .A3(G264), .A4(G1698), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT83), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n460), .A2(new_n461), .A3(new_n462), .A4(KEYINPUT83), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n465), .A2(new_n269), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT5), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n260), .B(G45), .C1(new_n468), .C2(G41), .ZN(new_n469));
  INV_X1    g0269(.A(G274), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n278), .A2(KEYINPUT5), .ZN(new_n471));
  OR3_X1    g0271(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  OAI211_X1 g0272(.A(G270), .B(new_n345), .C1(new_n469), .C2(new_n471), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n467), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n261), .A2(G116), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n260), .A2(G33), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n249), .A2(new_n261), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(G116), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n247), .A2(new_n225), .B1(G20), .B2(new_n481), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G283), .ZN(new_n485));
  INV_X1    g0285(.A(G97), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n485), .B(new_n226), .C1(G33), .C2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT20), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n484), .A2(KEYINPUT20), .A3(new_n487), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n268), .B1(new_n483), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n476), .A2(new_n492), .A3(KEYINPUT21), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT21), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n345), .B1(new_n463), .B2(new_n464), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n474), .B1(new_n495), .B2(new_n466), .ZN(new_n496));
  AND3_X1   g0296(.A1(new_n484), .A2(KEYINPUT20), .A3(new_n487), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(new_n488), .ZN(new_n498));
  OAI21_X1  g0298(.A(G169), .B1(new_n498), .B2(new_n482), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n494), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n483), .A2(new_n491), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n496), .A2(G179), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n493), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n336), .A2(new_n338), .A3(new_n226), .A4(G87), .ZN(new_n504));
  XNOR2_X1  g0304(.A(new_n504), .B(KEYINPUT22), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT24), .ZN(new_n506));
  XNOR2_X1  g0306(.A(KEYINPUT69), .B(G107), .ZN(new_n507));
  OAI21_X1  g0307(.A(KEYINPUT23), .B1(new_n507), .B2(new_n226), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n226), .A2(KEYINPUT23), .A3(G107), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT84), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G116), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n510), .B1(new_n511), .B2(G20), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n226), .A2(KEYINPUT84), .A3(G33), .A4(G116), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n505), .A2(new_n506), .A3(new_n508), .A4(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT22), .ZN(new_n516));
  XNOR2_X1  g0316(.A(new_n504), .B(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n508), .A2(new_n514), .ZN(new_n518));
  OAI21_X1  g0318(.A(KEYINPUT24), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n515), .B1(new_n519), .B2(KEYINPUT85), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT85), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n505), .A2(new_n508), .A3(new_n514), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n521), .B1(new_n522), .B2(KEYINPUT24), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n248), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(G107), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n262), .A2(new_n525), .ZN(new_n526));
  OR2_X1    g0326(.A1(new_n526), .A2(KEYINPUT25), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(KEYINPUT25), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n527), .B(new_n528), .C1(new_n525), .C2(new_n480), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n524), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(G264), .B(new_n345), .C1(new_n469), .C2(new_n471), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n336), .A2(new_n338), .A3(G250), .A4(new_n275), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n336), .A2(new_n338), .A3(G257), .A4(G1698), .ZN(new_n535));
  INV_X1    g0335(.A(G294), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n534), .B(new_n535), .C1(new_n335), .C2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n533), .B1(new_n537), .B2(new_n269), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n472), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n268), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(G179), .B2(new_n539), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n503), .B1(new_n531), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(G87), .A2(G97), .ZN(new_n544));
  NAND3_X1  g0344(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n301), .A2(new_n544), .B1(new_n226), .B2(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n336), .A2(new_n338), .A3(new_n226), .A4(G68), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n256), .A2(new_n486), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n547), .B1(KEYINPUT19), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n248), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n317), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n262), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n336), .A2(new_n338), .A3(G244), .A4(G1698), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n336), .A2(new_n338), .A3(G238), .A4(new_n275), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(new_n555), .A3(new_n511), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n269), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n260), .A2(G45), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G250), .ZN(new_n559));
  OAI22_X1  g0359(.A1(new_n269), .A2(new_n559), .B1(new_n470), .B2(new_n558), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(G200), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n560), .B1(new_n556), .B2(new_n269), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G190), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n249), .A2(G87), .A3(new_n261), .A4(new_n479), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n553), .A2(new_n563), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n550), .B(new_n552), .C1(new_n551), .C2(new_n480), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n562), .A2(new_n268), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n564), .A2(new_n288), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT6), .ZN(new_n573));
  NAND2_X1  g0373(.A1(G97), .A2(G107), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n207), .A2(KEYINPUT81), .A3(new_n573), .A4(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(KEYINPUT81), .ZN(new_n576));
  INV_X1    g0376(.A(new_n574), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n576), .B1(new_n577), .B2(new_n206), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n486), .A2(KEYINPUT6), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n575), .A2(new_n578), .A3(G20), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n250), .A2(G77), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n507), .B1(new_n365), .B2(new_n367), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT82), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(KEYINPUT82), .B(new_n507), .C1(new_n365), .C2(new_n367), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n249), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n262), .A2(new_n486), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n480), .B2(new_n486), .ZN(new_n589));
  OAI211_X1 g0389(.A(G257), .B(new_n345), .C1(new_n469), .C2(new_n471), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n472), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n336), .A2(new_n338), .A3(G244), .A4(new_n275), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT4), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n270), .A2(KEYINPUT4), .A3(G244), .A4(new_n275), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n270), .A2(G250), .A3(G1698), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n594), .A2(new_n595), .A3(new_n485), .A4(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n591), .B1(new_n597), .B2(new_n269), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n598), .A2(G179), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n598), .A2(new_n268), .ZN(new_n600));
  OAI22_X1  g0400(.A1(new_n587), .A2(new_n589), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n583), .A2(new_n584), .ZN(new_n602));
  INV_X1    g0402(.A(new_n582), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(new_n603), .A3(new_n586), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n248), .ZN(new_n605));
  INV_X1    g0405(.A(new_n589), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n597), .A2(new_n269), .ZN(new_n607));
  INV_X1    g0407(.A(new_n591), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(G200), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n598), .A2(G190), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n605), .A2(new_n606), .A3(new_n610), .A4(new_n611), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n572), .A2(new_n601), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n501), .B1(new_n476), .B2(G200), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n496), .A2(new_n357), .A3(new_n358), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(G190), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n538), .A2(new_n617), .A3(new_n472), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT86), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n538), .A2(KEYINPUT86), .A3(new_n617), .A4(new_n472), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n539), .A2(new_n293), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n524), .A2(new_n530), .A3(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n543), .A2(new_n613), .A3(new_n616), .A4(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n457), .A2(new_n625), .ZN(G372));
  NOR2_X1   g0426(.A1(new_n410), .A2(new_n456), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n624), .A2(new_n572), .A3(new_n601), .A4(new_n612), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT87), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n503), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n493), .A2(new_n500), .A3(KEYINPUT87), .A4(new_n502), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n531), .A2(new_n542), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n628), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n598), .A2(G179), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n268), .B2(new_n598), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT88), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n636), .A2(new_n637), .B1(new_n605), .B2(new_n606), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n635), .B(KEYINPUT88), .C1(new_n268), .C2(new_n598), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n638), .A2(new_n639), .A3(new_n572), .A4(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n567), .A2(new_n571), .ZN(new_n642));
  OAI21_X1  g0442(.A(KEYINPUT26), .B1(new_n601), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n641), .A2(new_n571), .A3(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n627), .B1(new_n634), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n295), .A2(new_n298), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n395), .A2(new_n455), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n440), .A2(new_n442), .A3(new_n448), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT75), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n450), .A2(KEYINPUT75), .A3(new_n442), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n421), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n327), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n648), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n646), .B1(new_n655), .B2(new_n407), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n656), .A2(KEYINPUT89), .A3(new_n330), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT89), .ZN(new_n658));
  INV_X1    g0458(.A(new_n646), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n647), .B1(new_n452), .B2(new_n327), .ZN(new_n660));
  INV_X1    g0460(.A(new_n407), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n658), .B1(new_n662), .B2(new_n290), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n645), .B1(new_n657), .B2(new_n663), .ZN(G369));
  INV_X1    g0464(.A(G13), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n665), .A2(G20), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n260), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(G213), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(G343), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n501), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n503), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n630), .A2(new_n631), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n616), .B(new_n674), .C1(new_n675), .C2(new_n673), .ZN(new_n676));
  INV_X1    g0476(.A(G330), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n633), .A2(new_n624), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n522), .A2(new_n521), .A3(KEYINPUT24), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n519), .A2(KEYINPUT85), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(new_n682), .A3(new_n515), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n529), .B1(new_n683), .B2(new_n248), .ZN(new_n684));
  INV_X1    g0484(.A(new_n672), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n684), .A2(new_n541), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n687), .B1(new_n688), .B2(new_n672), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n679), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n503), .A2(new_n685), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n687), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g0493(.A(new_n672), .B(KEYINPUT90), .Z(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n688), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(KEYINPUT91), .B1(new_n693), .B2(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n693), .A2(KEYINPUT91), .A3(new_n696), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n691), .B1(new_n697), .B2(new_n699), .ZN(G399));
  NAND3_X1  g0500(.A1(new_n301), .A2(new_n481), .A3(new_n544), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n211), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(G41), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(G1), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n228), .B2(new_n705), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT28), .ZN(new_n708));
  INV_X1    g0508(.A(new_n644), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n624), .B(new_n613), .C1(new_n675), .C2(new_n688), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n694), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT29), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n638), .A2(new_n640), .ZN(new_n714));
  OAI21_X1  g0514(.A(KEYINPUT26), .B1(new_n714), .B2(new_n642), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n571), .B(KEYINPUT93), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n601), .A2(new_n642), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n716), .B1(new_n717), .B2(new_n639), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n715), .B(new_n718), .C1(new_n543), .C2(new_n628), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n712), .B1(new_n719), .B2(new_n685), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n713), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n537), .A2(new_n269), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n564), .A2(new_n723), .A3(new_n532), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT92), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT92), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n538), .A2(new_n726), .A3(new_n564), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n725), .A2(new_n598), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n496), .A2(G179), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n722), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n609), .B1(KEYINPUT92), .B2(new_n724), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n476), .A2(new_n288), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n731), .A2(new_n732), .A3(KEYINPUT30), .A4(new_n727), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n598), .A2(G179), .A3(new_n564), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n734), .A2(new_n476), .A3(new_n539), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n730), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(new_n672), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT31), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n736), .A2(KEYINPUT31), .A3(new_n694), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n739), .B(new_n740), .C1(new_n625), .C2(new_n694), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G330), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n721), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n708), .B1(new_n744), .B2(G1), .ZN(G364));
  AOI21_X1  g0545(.A(new_n260), .B1(new_n666), .B2(G45), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n704), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G13), .A2(G33), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  AND2_X1   g0551(.A1(new_n676), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n225), .B1(G20), .B2(new_n268), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n211), .A2(G116), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n703), .A2(new_n270), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n757), .B1(new_n244), .B2(new_n279), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n758), .B1(new_n279), .B2(new_n229), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n703), .A2(new_n366), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT94), .ZN(new_n761));
  AOI211_X1 g0561(.A(new_n756), .B(new_n759), .C1(G355), .C2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n293), .A2(G179), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n226), .A2(G190), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n525), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n226), .A2(new_n288), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G200), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n359), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n766), .B1(G50), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n767), .A2(new_n293), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n359), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n768), .A2(G190), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OAI221_X1 g0575(.A(new_n770), .B1(new_n215), .B2(new_n773), .C1(new_n217), .C2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n771), .A2(G190), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n273), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G179), .A2(G200), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n226), .B1(new_n780), .B2(G190), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n486), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n764), .A2(new_n780), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G159), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT32), .ZN(new_n786));
  NOR4_X1   g0586(.A1(new_n776), .A2(new_n779), .A3(new_n782), .A4(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n763), .A2(G20), .A3(G190), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G87), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(new_n270), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n791), .B(KEYINPUT95), .Z(new_n792));
  INV_X1    g0592(.A(G317), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(KEYINPUT33), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n793), .A2(KEYINPUT33), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n774), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n777), .A2(G311), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n772), .A2(G322), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G303), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n366), .B1(new_n788), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G283), .ZN(new_n802));
  INV_X1    g0602(.A(G329), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n765), .A2(new_n802), .B1(new_n783), .B2(new_n803), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n799), .A2(new_n801), .A3(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n781), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n769), .A2(G326), .B1(G294), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT96), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n787), .A2(new_n792), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n753), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n755), .A2(new_n762), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n748), .B1(new_n752), .B2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n748), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n676), .A2(new_n677), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n814), .B2(new_n678), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT97), .Z(G396));
  AND4_X1   g0617(.A1(new_n326), .A2(new_n324), .A3(new_n325), .A4(new_n685), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT99), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n322), .B2(new_n685), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n326), .A2(KEYINPUT99), .A3(new_n672), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n323), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n818), .B1(new_n822), .B2(new_n327), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n711), .B(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n748), .B1(new_n824), .B2(new_n742), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n742), .B2(new_n824), .ZN(new_n826));
  INV_X1    g0626(.A(new_n765), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n827), .A2(G87), .B1(new_n784), .B2(G311), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT98), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n270), .B(new_n782), .C1(G107), .C2(new_n789), .ZN(new_n830));
  AOI22_X1  g0630(.A1(G283), .A2(new_n774), .B1(new_n772), .B2(G294), .ZN(new_n831));
  AOI22_X1  g0631(.A1(G303), .A2(new_n769), .B1(new_n777), .B2(G116), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n829), .A2(new_n830), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  AOI22_X1  g0633(.A1(G143), .A2(new_n772), .B1(new_n774), .B2(G150), .ZN(new_n834));
  INV_X1    g0634(.A(G137), .ZN(new_n835));
  INV_X1    g0635(.A(new_n769), .ZN(new_n836));
  INV_X1    g0636(.A(G159), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n834), .B1(new_n835), .B2(new_n836), .C1(new_n837), .C2(new_n778), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT34), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n789), .A2(G50), .B1(new_n784), .B2(G132), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n827), .A2(G68), .ZN(new_n842));
  AND3_X1   g0642(.A1(new_n841), .A2(new_n270), .A3(new_n842), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n840), .B(new_n843), .C1(new_n215), .C2(new_n781), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n838), .A2(new_n839), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n833), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n753), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n753), .A2(new_n749), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n813), .B1(new_n273), .B2(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n847), .B(new_n849), .C1(new_n823), .C2(new_n750), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n826), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(G384));
  AND3_X1   g0652(.A1(new_n575), .A2(new_n578), .A3(new_n579), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n853), .A2(KEYINPUT35), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(KEYINPUT35), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n854), .A2(G116), .A3(new_n227), .A4(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT36), .ZN(new_n857));
  OR2_X1    g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n856), .A2(new_n857), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n201), .A2(new_n217), .ZN(new_n860));
  NOR3_X1   g0660(.A1(new_n369), .A2(new_n228), .A3(new_n273), .ZN(new_n861));
  OAI211_X1 g0661(.A(G1), .B(new_n665), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n858), .A2(new_n859), .A3(new_n862), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT100), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n422), .A2(new_n672), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n452), .A2(new_n455), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n653), .A2(new_n672), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n670), .B1(new_n380), .B2(new_n386), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n408), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n670), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n390), .B1(new_n405), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n390), .A2(new_n871), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT101), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n363), .A2(new_n387), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n872), .A2(new_n874), .A3(KEYINPUT37), .A4(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT101), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT37), .B1(new_n869), .B2(new_n877), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n400), .A2(new_n670), .B1(new_n380), .B2(new_n386), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n878), .B1(new_n879), .B2(new_n393), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n870), .A2(new_n881), .A3(KEYINPUT38), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n873), .B1(new_n395), .B2(new_n407), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n876), .A2(new_n880), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n736), .A2(KEYINPUT31), .A3(new_n672), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n888), .B(new_n739), .C1(new_n625), .C2(new_n694), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n868), .A2(new_n887), .A3(new_n823), .A4(new_n889), .ZN(new_n890));
  XOR2_X1   g0690(.A(KEYINPUT104), .B(KEYINPUT40), .Z(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT37), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n879), .B2(new_n393), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n872), .A2(KEYINPUT37), .A3(new_n875), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT102), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n363), .A2(new_n387), .A3(new_n388), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n394), .B1(new_n363), .B2(new_n387), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n389), .B(KEYINPUT102), .C1(new_n393), .C2(new_n394), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n901), .A2(new_n407), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n897), .B1(new_n903), .B2(new_n869), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n882), .B1(new_n904), .B2(KEYINPUT38), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n889), .A2(new_n823), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n905), .A2(new_n906), .A3(KEYINPUT40), .A4(new_n868), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n893), .A2(G330), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n627), .A2(G330), .A3(new_n889), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n910), .B(KEYINPUT105), .Z(new_n911));
  NAND4_X1  g0711(.A1(new_n893), .A2(new_n907), .A3(new_n627), .A4(new_n889), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n657), .A2(new_n663), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n627), .B1(new_n713), .B2(new_n720), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n913), .B(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n452), .A2(new_n672), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT39), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n921), .B(new_n882), .C1(new_n904), .C2(KEYINPUT38), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT38), .B1(new_n870), .B2(new_n881), .ZN(new_n923));
  NOR3_X1   g0723(.A1(new_n884), .A2(new_n885), .A3(new_n883), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT39), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(KEYINPUT103), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT103), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n922), .A2(new_n925), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n920), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n695), .B(new_n823), .C1(new_n634), .C2(new_n644), .ZN(new_n931));
  INV_X1    g0731(.A(new_n818), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n931), .A2(new_n932), .B1(new_n866), .B2(new_n867), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n887), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n661), .A2(new_n670), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n930), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n918), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n260), .B2(new_n666), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n918), .A2(new_n937), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n864), .B1(new_n939), .B2(new_n940), .ZN(G367));
  NOR2_X1   g0741(.A1(new_n714), .A2(new_n695), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n694), .B1(new_n587), .B2(new_n589), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n943), .A2(new_n601), .A3(new_n612), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n944), .A2(KEYINPUT106), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(KEYINPUT106), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n942), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n688), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n694), .B1(new_n949), .B2(new_n601), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n947), .A2(new_n693), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT42), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n553), .A2(new_n566), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n672), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n572), .A2(new_n956), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n956), .A2(new_n571), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT43), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n954), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n951), .A2(new_n953), .A3(new_n961), .A4(new_n960), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n691), .A2(new_n947), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n966), .B(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n704), .B(KEYINPUT41), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n948), .B1(new_n699), .B2(new_n697), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT45), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n948), .B(KEYINPUT45), .C1(new_n699), .C2(new_n697), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n697), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n976), .A2(new_n698), .A3(new_n947), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT44), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n976), .A2(KEYINPUT44), .A3(new_n698), .A4(new_n947), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n975), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n690), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n975), .A2(new_n981), .A3(new_n691), .ZN(new_n984));
  INV_X1    g0784(.A(new_n689), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n693), .B1(new_n985), .B2(new_n692), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(new_n679), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n987), .A2(new_n743), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n983), .A2(new_n984), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n970), .B1(new_n989), .B2(new_n744), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n968), .B1(new_n990), .B2(new_n747), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n765), .A2(new_n273), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n270), .B1(new_n788), .B2(new_n215), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(G137), .C2(new_n784), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n772), .A2(G150), .ZN(new_n995));
  AOI22_X1  g0795(.A1(G143), .A2(new_n769), .B1(new_n774), .B2(G159), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n777), .A2(new_n201), .B1(G68), .B2(new_n806), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n994), .A2(new_n995), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(KEYINPUT109), .B1(new_n789), .B2(G116), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT46), .Z(new_n1000));
  OAI221_X1 g0800(.A(new_n366), .B1(new_n783), .B2(new_n793), .C1(new_n486), .C2(new_n765), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n775), .A2(new_n536), .B1(new_n301), .B2(new_n781), .ZN(new_n1002));
  OR3_X1    g0802(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(KEYINPUT108), .B(G311), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n769), .A2(new_n1004), .B1(new_n777), .B2(G283), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n800), .B2(new_n773), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n998), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT110), .Z(new_n1008));
  AOI21_X1  g0808(.A(new_n810), .B1(new_n1008), .B2(KEYINPUT47), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(KEYINPUT47), .B2(new_n1008), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n960), .A2(new_n751), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n757), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n754), .B1(new_n211), .B2(new_n551), .C1(new_n237), .C2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n748), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT107), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1010), .A2(new_n1011), .A3(new_n1015), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT111), .Z(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n991), .A2(new_n1018), .ZN(G387));
  INV_X1    g0819(.A(new_n987), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n689), .A2(new_n751), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n757), .B1(new_n234), .B2(new_n279), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n761), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1022), .B1(new_n702), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n314), .A2(G50), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT50), .ZN(new_n1026));
  AOI21_X1  g0826(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1026), .A2(new_n702), .A3(new_n1027), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n1024), .A2(new_n1028), .B1(new_n525), .B2(new_n703), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n748), .B1(new_n1029), .B2(new_n755), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n789), .A2(G77), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(KEYINPUT112), .B(G150), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1031), .B1(new_n783), .B2(new_n1033), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n366), .B(new_n1034), .C1(G97), .C2(new_n827), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(G159), .A2(new_n769), .B1(new_n777), .B2(G68), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n772), .A2(G50), .B1(new_n317), .B2(new_n806), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n774), .A2(new_n255), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n270), .B1(new_n784), .B2(G326), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n774), .A2(new_n1004), .B1(new_n777), .B2(G303), .ZN(new_n1041));
  XOR2_X1   g0841(.A(KEYINPUT113), .B(G322), .Z(new_n1042));
  OAI221_X1 g0842(.A(new_n1041), .B1(new_n793), .B2(new_n773), .C1(new_n836), .C2(new_n1042), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT48), .Z(new_n1044));
  OAI22_X1  g0844(.A1(new_n788), .A2(new_n536), .B1(new_n781), .B2(new_n802), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1040), .B1(new_n481), .B2(new_n765), .C1(new_n1046), .C2(KEYINPUT49), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n1046), .A2(KEYINPUT49), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1039), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1030), .B1(new_n1049), .B2(new_n753), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n1020), .A2(new_n747), .B1(new_n1021), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n988), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n704), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1020), .A2(new_n744), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1051), .B1(new_n1053), .B2(new_n1054), .ZN(G393));
  NAND3_X1  g0855(.A1(new_n983), .A2(new_n747), .A3(new_n984), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n947), .A2(new_n751), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n1042), .A2(new_n783), .B1(new_n788), .B2(new_n802), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT114), .Z(new_n1059));
  AOI211_X1 g0859(.A(new_n270), .B(new_n766), .C1(G303), .C2(new_n774), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n777), .A2(G294), .B1(G116), .B2(new_n806), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G311), .A2(new_n772), .B1(new_n769), .B2(G317), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT52), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G150), .A2(new_n769), .B1(new_n772), .B2(G159), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT51), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n777), .A2(new_n315), .B1(G77), .B2(new_n806), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n366), .B1(new_n827), .B2(G87), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n789), .A2(G68), .B1(new_n784), .B2(G143), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n774), .A2(new_n201), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n1062), .A2(new_n1064), .B1(new_n1066), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n753), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n755), .B1(G97), .B2(new_n703), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n241), .A2(new_n757), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n813), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1057), .A2(new_n1073), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1056), .A2(new_n1077), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n975), .A2(new_n981), .A3(new_n691), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n691), .B1(new_n975), .B2(new_n981), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n705), .B1(new_n1081), .B2(new_n988), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1052), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1078), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(G390));
  NAND2_X1  g0885(.A1(new_n931), .A2(new_n932), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n868), .A2(G330), .A3(new_n823), .A4(new_n889), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n741), .A2(G330), .A3(new_n823), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1088), .A2(new_n866), .A3(new_n867), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n889), .A2(G330), .A3(new_n823), .ZN(new_n1091));
  AND3_X1   g0891(.A1(new_n866), .A2(KEYINPUT115), .A3(new_n867), .ZN(new_n1092));
  AOI21_X1  g0892(.A(KEYINPUT115), .B1(new_n866), .B2(new_n867), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1091), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n822), .A2(new_n327), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n719), .A2(new_n685), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n932), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n741), .A2(G330), .A3(new_n823), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1097), .B1(new_n1098), .B2(new_n868), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n1086), .A2(new_n1090), .B1(new_n1094), .B2(new_n1099), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n915), .B(new_n909), .C1(new_n657), .C2(new_n663), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n905), .A2(new_n920), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1104), .B1(new_n1105), .B2(new_n1097), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1086), .A2(new_n868), .ZN(new_n1107));
  AOI21_X1  g0907(.A(KEYINPUT116), .B1(new_n1107), .B2(new_n920), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT116), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1109), .B(new_n919), .C1(new_n1086), .C2(new_n868), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n922), .A2(new_n925), .A3(new_n928), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n928), .B1(new_n922), .B2(new_n925), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1106), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1115), .A2(new_n1087), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1109), .B1(new_n933), .B2(new_n919), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n866), .A2(new_n867), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n818), .B1(new_n711), .B2(new_n823), .ZN(new_n1119));
  OAI211_X1 g0919(.A(KEYINPUT116), .B(new_n920), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n927), .A2(new_n1117), .A3(new_n929), .A4(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1092), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1093), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1122), .A2(new_n1097), .A3(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1124), .A2(new_n920), .A3(new_n905), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1098), .A2(new_n868), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1121), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1103), .B1(new_n1116), .B2(new_n1128), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1102), .B(new_n1127), .C1(new_n1115), .C2(new_n1087), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1129), .A2(new_n704), .A3(new_n1130), .ZN(new_n1131));
  NOR3_X1   g0931(.A1(new_n1112), .A2(new_n1113), .A3(new_n750), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n848), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(G116), .A2(new_n772), .B1(new_n774), .B2(new_n507), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n486), .B2(new_n778), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n784), .A2(G294), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n790), .A2(new_n842), .A3(new_n1136), .A4(new_n366), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n836), .A2(new_n802), .B1(new_n273), .B2(new_n781), .ZN(new_n1138));
  NOR3_X1   g0938(.A1(new_n1135), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1033), .A2(new_n788), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n1142));
  INV_X1    g0942(.A(G128), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n1141), .A2(new_n1142), .B1(new_n836), .B2(new_n1143), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1141), .A2(new_n1142), .B1(new_n772), .B2(G132), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n366), .B1(new_n784), .B2(G125), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1145), .B(new_n1146), .C1(new_n202), .C2(new_n765), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n1144), .B(new_n1147), .C1(G159), .C2(new_n806), .ZN(new_n1148));
  XOR2_X1   g0948(.A(KEYINPUT54), .B(G143), .Z(new_n1149));
  AOI22_X1  g0949(.A1(G137), .A2(new_n774), .B1(new_n777), .B2(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(KEYINPUT117), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1139), .B1(new_n1148), .B2(new_n1152), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n748), .B1(new_n255), .B2(new_n1133), .C1(new_n1153), .C2(new_n810), .ZN(new_n1154));
  OR3_X1    g0954(.A1(new_n1132), .A2(KEYINPUT119), .A3(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(KEYINPUT119), .B1(new_n1132), .B2(new_n1154), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1116), .A2(new_n1128), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1157), .B1(new_n1158), .B2(new_n747), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1131), .A2(new_n1159), .ZN(G378));
  NOR2_X1   g0960(.A1(new_n267), .A2(new_n670), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n333), .B(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1163));
  XOR2_X1   g0963(.A(new_n1162), .B(new_n1163), .Z(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n919), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n936), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1166), .A2(new_n1167), .A3(new_n908), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n908), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1165), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n908), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n930), .B2(new_n936), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1166), .A2(new_n1167), .A3(new_n908), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1172), .A2(new_n1173), .A3(new_n1164), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1170), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1101), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1130), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT57), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n705), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1175), .A2(new_n1177), .A3(KEYINPUT57), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(KEYINPUT122), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT122), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1175), .A2(new_n1177), .A3(new_n1183), .A4(KEYINPUT57), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1180), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n813), .B1(new_n202), .B2(new_n848), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n772), .A2(G128), .B1(new_n789), .B2(new_n1149), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT120), .Z(new_n1188));
  AOI22_X1  g0988(.A1(new_n774), .A2(G132), .B1(G150), .B2(new_n806), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(G125), .A2(new_n769), .B1(new_n777), .B2(G137), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT59), .Z(new_n1192));
  AOI211_X1 g0992(.A(G33), .B(G41), .C1(new_n784), .C2(G124), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1192), .B(new_n1193), .C1(new_n837), .C2(new_n765), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n773), .A2(new_n525), .B1(new_n775), .B2(new_n486), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n765), .A2(new_n215), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(G283), .B2(new_n784), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n777), .A2(new_n317), .B1(G68), .B2(new_n806), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n270), .A2(G41), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1197), .A2(new_n1198), .A3(new_n1031), .A4(new_n1199), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1195), .B(new_n1200), .C1(G116), .C2(new_n769), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(KEYINPUT58), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1199), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1203), .B(new_n263), .C1(G33), .C2(G41), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1201), .A2(KEYINPUT58), .ZN(new_n1205));
  AND4_X1   g1005(.A1(new_n1194), .A2(new_n1202), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1186), .B1(new_n810), .B2(new_n1206), .C1(new_n1165), .C2(new_n750), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT121), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n1175), .B2(new_n747), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1185), .A2(new_n1209), .ZN(G375));
  OAI22_X1  g1010(.A1(new_n802), .A2(new_n773), .B1(new_n778), .B2(new_n301), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(G294), .B2(new_n769), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n775), .A2(new_n481), .B1(new_n551), .B2(new_n781), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n788), .A2(new_n486), .B1(new_n783), .B2(new_n800), .ZN(new_n1214));
  NOR4_X1   g1014(.A1(new_n1213), .A2(new_n1214), .A3(new_n270), .A4(new_n992), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n774), .A2(new_n1149), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n773), .B2(new_n835), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n788), .A2(new_n837), .B1(new_n783), .B2(new_n1143), .ZN(new_n1218));
  NOR4_X1   g1018(.A1(new_n1217), .A2(new_n366), .A3(new_n1196), .A4(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n769), .A2(G132), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n263), .B2(new_n781), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(G150), .B2(new_n777), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1212), .A2(new_n1215), .B1(new_n1219), .B2(new_n1222), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n748), .B1(G68), .B2(new_n1133), .C1(new_n1223), .C2(new_n810), .ZN(new_n1224));
  XOR2_X1   g1024(.A(new_n1224), .B(KEYINPUT123), .Z(new_n1225));
  INV_X1    g1025(.A(new_n1105), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1225), .B1(new_n1226), .B2(new_n749), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1100), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1227), .B1(new_n1228), .B2(new_n747), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1103), .A2(new_n969), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1228), .A2(new_n1176), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1229), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(KEYINPUT124), .ZN(G381));
  INV_X1    g1033(.A(G378), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1185), .A2(new_n1234), .A3(new_n1209), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n991), .A2(new_n1018), .A3(new_n1084), .ZN(new_n1236));
  OR3_X1    g1036(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1237));
  OR4_X1    g1037(.A1(G381), .A2(new_n1235), .A3(new_n1236), .A4(new_n1237), .ZN(G407));
  OAI211_X1 g1038(.A(G407), .B(G213), .C1(G343), .C2(new_n1235), .ZN(G409));
  AND3_X1   g1039(.A1(new_n991), .A2(new_n1018), .A3(new_n1084), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1084), .B1(new_n991), .B2(new_n1018), .ZN(new_n1241));
  OAI21_X1  g1041(.A(KEYINPUT125), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(G387), .A2(G390), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT125), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1243), .A2(new_n1244), .A3(new_n1236), .ZN(new_n1245));
  XOR2_X1   g1045(.A(G393), .B(G396), .Z(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1242), .A2(new_n1245), .A3(new_n1247), .ZN(new_n1248));
  OAI211_X1 g1048(.A(KEYINPUT125), .B(new_n1246), .C1(new_n1240), .C2(new_n1241), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT61), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT60), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n1228), .B2(new_n1176), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1100), .A2(new_n1101), .A3(KEYINPUT60), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1253), .A2(new_n704), .A3(new_n1103), .A4(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1229), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n851), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1255), .A2(G384), .A3(new_n1229), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n671), .A2(G213), .A3(G2897), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1259), .B(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1234), .B1(new_n1185), .B2(new_n1209), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1175), .A2(new_n747), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1131), .A2(new_n1159), .A3(new_n1263), .A4(new_n1207), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1178), .A2(new_n970), .ZN(new_n1265));
  INV_X1    g1065(.A(G213), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n1264), .A2(new_n1265), .B1(new_n1266), .B2(G343), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1261), .B1(new_n1262), .B2(new_n1267), .ZN(new_n1268));
  NOR3_X1   g1068(.A1(new_n1262), .A2(new_n1267), .A3(new_n1259), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT62), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1251), .B(new_n1268), .C1(new_n1269), .C2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(G375), .A2(G378), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1267), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1259), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1272), .A2(new_n1273), .A3(new_n1274), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1275), .A2(KEYINPUT62), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1250), .B1(new_n1271), .B2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT126), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT63), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1275), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1268), .A2(new_n1251), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1269), .A2(KEYINPUT126), .A3(KEYINPUT63), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1248), .A2(new_n1249), .A3(new_n1283), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1280), .A2(new_n1281), .A3(new_n1282), .A4(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1277), .A2(new_n1285), .ZN(G405));
  NAND2_X1  g1086(.A1(new_n1272), .A2(new_n1235), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1259), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1248), .A2(KEYINPUT127), .A3(new_n1249), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1272), .A2(new_n1235), .A3(new_n1274), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1288), .A2(new_n1289), .A3(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT127), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT127), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1250), .A2(new_n1294), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1295), .A2(new_n1288), .A3(new_n1290), .A4(new_n1289), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1293), .A2(new_n1296), .ZN(G402));
endmodule


