//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0 1 1 1 1 0 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 0 1 1 1 0 0 0 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1263, new_n1264, new_n1265, new_n1266, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n202), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n208), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n211), .B(new_n216), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XOR2_X1   g0025(.A(G226), .B(G232), .Z(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT65), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n229), .B(new_n230), .Z(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G87), .B(G97), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT66), .ZN(new_n237));
  XOR2_X1   g0037(.A(G107), .B(G116), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  NOR2_X1   g0043(.A1(new_n206), .A2(G68), .ZN(new_n244));
  NOR2_X1   g0044(.A1(G20), .A2(G33), .ZN(new_n245));
  AOI21_X1  g0045(.A(new_n244), .B1(G50), .B2(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G77), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n206), .A2(G33), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n214), .ZN(new_n251));
  AND2_X1   g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  OR2_X1    g0052(.A1(new_n252), .A2(KEYINPUT11), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n251), .B1(new_n205), .B2(G20), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G68), .ZN(new_n255));
  XOR2_X1   g0055(.A(new_n255), .B(KEYINPUT71), .Z(new_n256));
  NAND2_X1  g0056(.A1(new_n252), .A2(KEYINPUT11), .ZN(new_n257));
  INV_X1    g0057(.A(G13), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G1), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT12), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n259), .B(new_n244), .C1(KEYINPUT72), .C2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(KEYINPUT72), .ZN(new_n262));
  XNOR2_X1  g0062(.A(new_n261), .B(new_n262), .ZN(new_n263));
  NAND4_X1  g0063(.A1(new_n253), .A2(new_n256), .A3(new_n257), .A4(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  AOI21_X1  g0068(.A(G1698), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G226), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n267), .A2(new_n268), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(G232), .A3(G1698), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G97), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n270), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G274), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n278));
  NOR3_X1   g0078(.A1(new_n275), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n214), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n282), .A2(new_n278), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n279), .B1(new_n283), .B2(G238), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n276), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT13), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT13), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n276), .A2(new_n287), .A3(new_n284), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT14), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n289), .A2(new_n290), .A3(G169), .ZN(new_n291));
  INV_X1    g0091(.A(G179), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n291), .B1(new_n292), .B2(new_n289), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n290), .B1(new_n289), .B2(G169), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n264), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G1698), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n271), .A2(G232), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G107), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n271), .A2(G1698), .ZN(new_n299));
  INV_X1    g0099(.A(G238), .ZN(new_n300));
  OAI221_X1 g0100(.A(new_n297), .B1(new_n298), .B2(new_n271), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n275), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n279), .B1(new_n283), .B2(G244), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n304), .A2(G179), .ZN(new_n305));
  INV_X1    g0105(.A(G169), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(G20), .A2(G77), .ZN(new_n308));
  XNOR2_X1  g0108(.A(KEYINPUT15), .B(G87), .ZN(new_n309));
  INV_X1    g0109(.A(new_n245), .ZN(new_n310));
  XNOR2_X1  g0110(.A(KEYINPUT8), .B(G58), .ZN(new_n311));
  OAI221_X1 g0111(.A(new_n308), .B1(new_n309), .B2(new_n248), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n251), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n254), .A2(G77), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n313), .B(new_n314), .C1(G77), .C2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n307), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n295), .B1(new_n305), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n269), .A2(G223), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n271), .A2(G226), .A3(G1698), .ZN(new_n320));
  NAND2_X1  g0120(.A1(G33), .A2(G87), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n275), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n279), .B1(new_n283), .B2(G232), .ZN(new_n324));
  AOI21_X1  g0124(.A(G169), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n324), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n325), .B1(new_n327), .B2(new_n292), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT16), .ZN(new_n329));
  INV_X1    g0129(.A(G68), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT7), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(new_n271), .B2(G20), .ZN(new_n332));
  AND2_X1   g0132(.A1(KEYINPUT3), .A2(G33), .ZN(new_n333));
  NOR2_X1   g0133(.A1(KEYINPUT3), .A2(G33), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n335), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n330), .B1(new_n332), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G58), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n338), .A2(new_n330), .ZN(new_n339));
  OAI21_X1  g0139(.A(G20), .B1(new_n339), .B2(new_n201), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n245), .A2(G159), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n329), .B1(new_n337), .B2(new_n342), .ZN(new_n343));
  NOR3_X1   g0143(.A1(new_n271), .A2(new_n331), .A3(G20), .ZN(new_n344));
  AOI21_X1  g0144(.A(KEYINPUT7), .B1(new_n335), .B2(new_n206), .ZN(new_n345));
  OAI21_X1  g0145(.A(G68), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n342), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(KEYINPUT16), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n343), .A2(new_n348), .A3(new_n251), .ZN(new_n349));
  NAND2_X1  g0149(.A1(KEYINPUT67), .A2(G58), .ZN(new_n350));
  XOR2_X1   g0150(.A(new_n350), .B(KEYINPUT8), .Z(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n352), .A2(new_n315), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n353), .B1(new_n352), .B2(new_n254), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n349), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n328), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT18), .ZN(new_n357));
  INV_X1    g0157(.A(new_n355), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n326), .A2(G200), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n323), .A2(G190), .A3(new_n324), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n358), .A2(new_n361), .A3(KEYINPUT17), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT18), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n328), .A2(new_n355), .A3(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n349), .A2(new_n359), .A3(new_n354), .A4(new_n360), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT17), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n357), .A2(new_n362), .A3(new_n364), .A4(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n368), .A2(KEYINPUT74), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n318), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT70), .ZN(new_n372));
  OR2_X1    g0172(.A1(new_n372), .A2(KEYINPUT10), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(KEYINPUT10), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n351), .A2(new_n248), .ZN(new_n375));
  OAI21_X1  g0175(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n376));
  INV_X1    g0176(.A(G150), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n376), .B1(new_n377), .B2(new_n310), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n251), .B1(new_n375), .B2(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n315), .A2(G50), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n380), .B1(new_n254), .B2(G50), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT68), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT68), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n379), .A2(new_n384), .A3(new_n381), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT9), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g0188(.A(new_n388), .B(KEYINPUT69), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n386), .A2(new_n387), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n269), .A2(G222), .ZN(new_n391));
  INV_X1    g0191(.A(G223), .ZN(new_n392));
  OAI221_X1 g0192(.A(new_n391), .B1(new_n247), .B2(new_n271), .C1(new_n392), .C2(new_n299), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n275), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n279), .B1(new_n283), .B2(G226), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G200), .ZN(new_n397));
  INV_X1    g0197(.A(G190), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n397), .B1(new_n398), .B2(new_n396), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n390), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n373), .B(new_n374), .C1(new_n389), .C2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT69), .ZN(new_n403));
  XNOR2_X1  g0203(.A(new_n388), .B(new_n403), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n404), .A2(new_n400), .A3(new_n372), .A4(KEYINPUT10), .ZN(new_n405));
  INV_X1    g0205(.A(new_n396), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n382), .B1(new_n406), .B2(G169), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n407), .B1(new_n292), .B2(new_n406), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n402), .A2(new_n405), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n368), .A2(KEYINPUT74), .ZN(new_n411));
  INV_X1    g0211(.A(new_n304), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n316), .B1(new_n412), .B2(G190), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n304), .A2(G200), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n286), .A2(new_n288), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n264), .B1(new_n416), .B2(G190), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n289), .A2(G200), .ZN(new_n418));
  AOI21_X1  g0218(.A(KEYINPUT73), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AND4_X1   g0219(.A1(new_n256), .A2(new_n253), .A3(new_n257), .A4(new_n263), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n286), .A2(G190), .A3(new_n288), .ZN(new_n421));
  AND4_X1   g0221(.A1(KEYINPUT73), .A2(new_n420), .A3(new_n418), .A4(new_n421), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n411), .B(new_n415), .C1(new_n419), .C2(new_n422), .ZN(new_n423));
  NOR3_X1   g0223(.A1(new_n371), .A2(new_n410), .A3(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n315), .B1(G1), .B2(new_n266), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n425), .A2(new_n251), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n427), .A2(new_n298), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n315), .A2(G107), .ZN(new_n429));
  XNOR2_X1  g0229(.A(KEYINPUT87), .B(KEYINPUT25), .ZN(new_n430));
  XNOR2_X1  g0230(.A(new_n429), .B(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n206), .B(G87), .C1(new_n333), .C2(new_n334), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT22), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT22), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n271), .A2(new_n436), .A3(new_n206), .A4(G87), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(G33), .A2(G116), .ZN(new_n439));
  OR3_X1    g0239(.A1(new_n439), .A2(KEYINPUT85), .A3(G20), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT23), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n206), .B2(G107), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n298), .A2(KEYINPUT23), .A3(G20), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(KEYINPUT85), .B1(new_n439), .B2(G20), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n440), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n438), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT86), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n438), .A2(KEYINPUT86), .A3(new_n446), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n449), .A2(new_n450), .A3(KEYINPUT24), .ZN(new_n451));
  INV_X1    g0251(.A(new_n251), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT86), .B1(new_n438), .B2(new_n446), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT24), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n433), .B1(new_n451), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(G41), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT5), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n205), .B(G45), .C1(new_n457), .C2(KEYINPUT5), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n282), .B(G264), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  OAI211_X1 g0262(.A(G257), .B(G1698), .C1(new_n333), .C2(new_n334), .ZN(new_n463));
  OAI211_X1 g0263(.A(G250), .B(new_n296), .C1(new_n333), .C2(new_n334), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G294), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n282), .B1(new_n466), .B2(KEYINPUT88), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT88), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n463), .A2(new_n464), .A3(new_n468), .A4(new_n465), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n462), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G45), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(G1), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT78), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n472), .B(new_n473), .C1(KEYINPUT5), .C2(new_n457), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n460), .A2(KEYINPUT78), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n277), .B1(new_n280), .B2(new_n281), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n474), .A2(new_n475), .A3(new_n476), .A4(new_n458), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n470), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(G200), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n470), .A2(G190), .A3(new_n477), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n456), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n478), .A2(G179), .ZN(new_n482));
  AOI21_X1  g0282(.A(G169), .B1(new_n470), .B2(new_n477), .ZN(new_n483));
  NOR3_X1   g0283(.A1(new_n456), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(KEYINPUT89), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n451), .A2(new_n455), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n432), .ZN(new_n487));
  INV_X1    g0287(.A(new_n483), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n487), .B(new_n488), .C1(G179), .C2(new_n478), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT89), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n456), .A2(new_n479), .A3(new_n480), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n485), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n282), .B(G257), .C1(new_n459), .C2(new_n460), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n477), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G33), .A2(G283), .ZN(new_n496));
  OAI211_X1 g0296(.A(G250), .B(G1698), .C1(new_n333), .C2(new_n334), .ZN(new_n497));
  OAI211_X1 g0297(.A(G244), .B(new_n296), .C1(new_n333), .C2(new_n334), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT4), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n496), .B(new_n497), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(KEYINPUT4), .B1(new_n269), .B2(G244), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n275), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n495), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n306), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(G179), .B2(new_n503), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n315), .A2(G97), .ZN(new_n507));
  XNOR2_X1  g0307(.A(new_n507), .B(KEYINPUT77), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n508), .B1(G97), .B2(new_n426), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT75), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n310), .A2(new_n247), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n298), .A2(KEYINPUT6), .A3(G97), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT6), .ZN(new_n515));
  XNOR2_X1  g0315(.A(G97), .B(G107), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n510), .B(new_n512), .C1(new_n517), .C2(new_n206), .ZN(new_n518));
  AND2_X1   g0318(.A1(G97), .A2(G107), .ZN(new_n519));
  NOR2_X1   g0319(.A1(G97), .A2(G107), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n515), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n206), .B1(new_n521), .B2(new_n513), .ZN(new_n522));
  OAI21_X1  g0322(.A(KEYINPUT75), .B1(new_n522), .B2(new_n511), .ZN(new_n523));
  OAI21_X1  g0323(.A(G107), .B1(new_n344), .B2(new_n345), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n518), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n525), .A2(KEYINPUT76), .A3(new_n251), .ZN(new_n526));
  AOI21_X1  g0326(.A(KEYINPUT76), .B1(new_n525), .B2(new_n251), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n509), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n506), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n525), .A2(new_n251), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT76), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n525), .A2(KEYINPUT76), .A3(new_n251), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT79), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G200), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n536), .B1(new_n495), .B2(new_n502), .ZN(new_n537));
  INV_X1    g0337(.A(new_n503), .ZN(new_n538));
  INV_X1    g0338(.A(G200), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n398), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n537), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n534), .A2(new_n509), .A3(new_n541), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n529), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(G87), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n427), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n206), .B(G68), .C1(new_n333), .C2(new_n334), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n206), .A2(G33), .A3(G97), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT19), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g0351(.A(KEYINPUT80), .B(G87), .ZN(new_n552));
  NAND3_X1  g0352(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n552), .A2(new_n520), .B1(new_n206), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n251), .B1(new_n551), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n309), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n556), .A2(new_n315), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  AND3_X1   g0358(.A1(new_n555), .A2(KEYINPUT81), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(KEYINPUT81), .B1(new_n555), .B2(new_n558), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n546), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n300), .A2(new_n296), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n271), .B(new_n562), .C1(G244), .C2(new_n296), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n282), .B1(new_n563), .B2(new_n439), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n282), .B1(G250), .B2(new_n472), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n277), .B2(new_n472), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n568), .A2(new_n398), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n567), .A2(new_n539), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n561), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n568), .A2(G169), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n567), .A2(G179), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT82), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT81), .ZN(new_n577));
  AOI21_X1  g0377(.A(G20), .B1(new_n267), .B2(new_n268), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n578), .A2(G68), .B1(new_n549), .B2(new_n548), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n552), .A2(new_n520), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n553), .A2(new_n206), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n452), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n577), .B1(new_n583), .B2(new_n557), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n555), .A2(KEYINPUT81), .A3(new_n558), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n427), .A2(new_n309), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n576), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  AOI211_X1 g0389(.A(KEYINPUT82), .B(new_n587), .C1(new_n584), .C2(new_n585), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n575), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n572), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g0392(.A(KEYINPUT83), .B(G303), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(G257), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n595), .B1(new_n267), .B2(new_n268), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n335), .A2(new_n594), .B1(new_n596), .B2(new_n296), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n271), .A2(G264), .A3(G1698), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n282), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n282), .B(G270), .C1(new_n459), .C2(new_n460), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n477), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(KEYINPUT84), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n601), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n271), .A2(G257), .A3(new_n296), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n598), .B(new_n604), .C1(new_n271), .C2(new_n593), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n275), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT84), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n603), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(G97), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n496), .B(new_n206), .C1(G33), .C2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(G116), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(G20), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n251), .A3(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT20), .ZN(new_n614));
  XNOR2_X1  g0414(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n315), .A2(G116), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(new_n426), .B2(G116), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n306), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n602), .A2(new_n608), .A3(new_n618), .A4(KEYINPUT21), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n599), .A2(new_n601), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n615), .A2(new_n617), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n620), .A2(G179), .A3(new_n621), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  NOR3_X1   g0423(.A1(new_n599), .A2(KEYINPUT84), .A3(new_n601), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n607), .B1(new_n603), .B2(new_n606), .ZN(new_n625));
  OAI21_X1  g0425(.A(G190), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n621), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n602), .A2(new_n608), .A3(G200), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n602), .A2(new_n608), .A3(new_n618), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT21), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n623), .A2(new_n629), .A3(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n592), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n424), .A2(new_n493), .A3(new_n543), .A4(new_n634), .ZN(new_n635));
  XOR2_X1   g0435(.A(new_n635), .B(KEYINPUT90), .Z(G372));
  NAND2_X1  g0436(.A1(new_n357), .A2(new_n364), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n318), .A2(new_n367), .A3(new_n362), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n417), .A2(new_n418), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n295), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n637), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n402), .A2(new_n405), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n409), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n424), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n586), .A2(new_n588), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n575), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT91), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n561), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n586), .A2(KEYINPUT91), .A3(new_n546), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n570), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT92), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n569), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n570), .ZN(new_n655));
  AOI21_X1  g0455(.A(KEYINPUT91), .B1(new_n586), .B2(new_n546), .ZN(new_n656));
  AOI211_X1 g0456(.A(new_n649), .B(new_n545), .C1(new_n584), .C2(new_n585), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(KEYINPUT92), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n648), .B1(new_n654), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n623), .A2(new_n632), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n481), .B1(new_n662), .B2(new_n489), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n660), .A2(new_n663), .A3(new_n543), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n505), .B1(new_n534), .B2(new_n509), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n572), .A2(new_n591), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n648), .B1(new_n667), .B2(KEYINPUT26), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n653), .B(new_n655), .C1(new_n656), .C2(new_n657), .ZN(new_n669));
  INV_X1    g0469(.A(new_n569), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n650), .A2(new_n651), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n653), .B1(new_n672), .B2(new_n655), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n666), .B(new_n647), .C1(new_n671), .C2(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n668), .B1(new_n674), .B2(KEYINPUT26), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT93), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI211_X1 g0477(.A(KEYINPUT93), .B(new_n668), .C1(new_n674), .C2(KEYINPUT26), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n665), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n644), .B1(new_n645), .B2(new_n679), .ZN(G369));
  NAND2_X1  g0480(.A1(new_n259), .A2(new_n206), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G213), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G343), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n627), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n661), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n633), .B2(new_n688), .ZN(new_n690));
  XOR2_X1   g0490(.A(new_n690), .B(KEYINPUT94), .Z(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G330), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n487), .A2(new_n686), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n493), .A2(new_n693), .B1(new_n484), .B2(new_n686), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n661), .A2(new_n687), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n697), .B1(new_n485), .B2(new_n492), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n698), .B1(new_n484), .B2(new_n687), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n696), .A2(new_n699), .ZN(G399));
  INV_X1    g0500(.A(new_n209), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(G41), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G1), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n552), .A2(new_n611), .A3(new_n520), .ZN(new_n705));
  OAI22_X1  g0505(.A1(new_n704), .A2(new_n705), .B1(new_n212), .B2(new_n703), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT28), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT29), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT96), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT26), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n709), .B1(new_n667), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n674), .B2(new_n710), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n660), .A2(new_n709), .A3(KEYINPUT26), .A4(new_n666), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT97), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n529), .A2(new_n714), .A3(new_n542), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n714), .B1(new_n529), .B2(new_n542), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(new_n660), .A3(new_n663), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n712), .A2(new_n713), .A3(new_n718), .A4(new_n647), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n708), .B1(new_n719), .B2(new_n687), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n679), .A2(new_n686), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n720), .B1(new_n721), .B2(new_n708), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT98), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n493), .A2(new_n634), .A3(new_n543), .A4(new_n687), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n538), .A2(G179), .A3(new_n620), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n470), .A2(KEYINPUT95), .A3(new_n567), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n470), .A2(new_n567), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT95), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n725), .B1(new_n726), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(KEYINPUT30), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n538), .A2(G179), .A3(new_n567), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n733), .A2(new_n478), .A3(new_n602), .A4(new_n608), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(new_n730), .B2(KEYINPUT30), .ZN(new_n735));
  OAI211_X1 g0535(.A(KEYINPUT31), .B(new_n686), .C1(new_n732), .C2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n686), .B1(new_n732), .B2(new_n735), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT31), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n724), .A2(new_n736), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G330), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n722), .A2(new_n723), .A3(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n678), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n659), .A2(new_n670), .A3(new_n669), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n744), .A2(new_n710), .A3(new_n666), .A4(new_n647), .ZN(new_n745));
  AOI21_X1  g0545(.A(KEYINPUT93), .B1(new_n745), .B2(new_n668), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n664), .B1(new_n743), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n747), .A2(new_n708), .A3(new_n687), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n719), .A2(new_n687), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(KEYINPUT29), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n741), .ZN(new_n752));
  OAI21_X1  g0552(.A(KEYINPUT98), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n742), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n707), .B1(new_n754), .B2(G1), .ZN(G364));
  NOR2_X1   g0555(.A1(new_n258), .A2(G20), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n205), .B1(new_n756), .B2(G45), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n702), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n759), .B1(new_n691), .B2(G330), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n760), .B1(G330), .B2(new_n691), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n701), .A2(new_n335), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G355), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(G116), .B2(new_n209), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n701), .A2(new_n271), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(new_n471), .B2(new_n213), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n242), .A2(G45), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n764), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n214), .B1(G20), .B2(new_n306), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n759), .B1(new_n769), .B2(new_n775), .ZN(new_n776));
  NOR4_X1   g0576(.A1(new_n206), .A2(new_n398), .A3(new_n539), .A4(G179), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G303), .ZN(new_n779));
  NOR4_X1   g0579(.A1(new_n206), .A2(new_n539), .A3(G179), .A4(G190), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G283), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n778), .A2(new_n779), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n206), .A2(new_n292), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G190), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n539), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G326), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n785), .A2(G200), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n783), .B(new_n789), .C1(G322), .C2(new_n790), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n292), .A2(new_n539), .A3(KEYINPUT99), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(KEYINPUT99), .B1(new_n292), .B2(new_n539), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n206), .B1(new_n796), .B2(G190), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G294), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n206), .A2(G190), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n795), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G329), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n784), .A2(new_n398), .A3(new_n539), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n805), .A2(G311), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n801), .A2(new_n292), .A3(new_n539), .ZN(new_n807));
  XNOR2_X1  g0607(.A(KEYINPUT33), .B(G317), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n271), .B(new_n806), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n791), .A2(new_n799), .A3(new_n803), .A4(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n802), .ZN(new_n811));
  XNOR2_X1  g0611(.A(KEYINPUT100), .B(G159), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT32), .Z(new_n814));
  NAND2_X1  g0614(.A1(new_n798), .A2(G97), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n271), .B1(new_n804), .B2(new_n247), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(G68), .B2(new_n807), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n781), .A2(new_n298), .ZN(new_n818));
  INV_X1    g0618(.A(new_n552), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n818), .B1(new_n819), .B2(new_n777), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n790), .A2(G58), .B1(new_n786), .B2(G50), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n815), .A2(new_n817), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n810), .B1(new_n814), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n776), .B1(new_n823), .B2(new_n773), .ZN(new_n824));
  INV_X1    g0624(.A(new_n772), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n824), .B1(new_n691), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n761), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(G396));
  INV_X1    g0628(.A(KEYINPUT104), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n317), .B2(new_n305), .ZN(new_n830));
  INV_X1    g0630(.A(new_n305), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n831), .A2(KEYINPUT104), .A3(new_n316), .A4(new_n307), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n316), .A2(new_n686), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n830), .A2(new_n832), .A3(new_n415), .A4(new_n833), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n831), .A2(new_n316), .A3(new_n307), .A4(new_n686), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n679), .B2(new_n686), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n830), .A2(new_n832), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n415), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n747), .A2(new_n687), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n837), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n752), .ZN(new_n844));
  INV_X1    g0644(.A(new_n759), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n837), .A2(new_n741), .A3(new_n842), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT105), .ZN(new_n848));
  INV_X1    g0648(.A(G294), .ZN(new_n849));
  INV_X1    g0649(.A(new_n790), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n849), .A2(new_n850), .B1(new_n787), .B2(new_n779), .ZN(new_n851));
  INV_X1    g0651(.A(new_n807), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n852), .A2(new_n782), .B1(new_n611), .B2(new_n804), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n781), .A2(new_n544), .ZN(new_n854));
  NOR3_X1   g0654(.A1(new_n851), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n271), .B1(new_n777), .B2(G107), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT101), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n802), .A2(G311), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n855), .A2(new_n815), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n781), .A2(new_n330), .ZN(new_n860));
  INV_X1    g0660(.A(G50), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n271), .B1(new_n778), .B2(new_n861), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n860), .B(new_n862), .C1(new_n802), .C2(G132), .ZN(new_n863));
  AOI22_X1  g0663(.A1(G150), .A2(new_n807), .B1(new_n786), .B2(G137), .ZN(new_n864));
  XOR2_X1   g0664(.A(new_n864), .B(KEYINPUT102), .Z(new_n865));
  NAND2_X1  g0665(.A1(new_n790), .A2(G143), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n865), .B(new_n866), .C1(new_n804), .C2(new_n812), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT103), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT34), .ZN(new_n869));
  OAI221_X1 g0669(.A(new_n863), .B1(new_n338), .B2(new_n797), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n868), .A2(new_n869), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n859), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n773), .A2(new_n770), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n872), .A2(new_n773), .B1(new_n247), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n836), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n874), .B1(new_n771), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n759), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n847), .A2(new_n848), .A3(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n848), .B1(new_n847), .B2(new_n877), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(G384));
  INV_X1    g0682(.A(new_n517), .ZN(new_n883));
  OR2_X1    g0683(.A1(new_n883), .A2(KEYINPUT35), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(KEYINPUT35), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n884), .A2(G116), .A3(new_n215), .A4(new_n885), .ZN(new_n886));
  XOR2_X1   g0686(.A(new_n886), .B(KEYINPUT36), .Z(new_n887));
  OR3_X1    g0687(.A1(new_n212), .A2(new_n247), .A3(new_n339), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n861), .A2(G68), .ZN(new_n889));
  AOI211_X1 g0689(.A(new_n205), .B(G13), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT108), .B1(new_n751), .B2(new_n424), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT108), .ZN(new_n893));
  AOI211_X1 g0693(.A(new_n893), .B(new_n645), .C1(new_n748), .C2(new_n750), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n644), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n420), .A2(new_n687), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n419), .A2(new_n422), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n293), .A2(new_n294), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n639), .A2(new_n896), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n295), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n839), .A2(new_n686), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n903), .B1(new_n842), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT38), .ZN(new_n907));
  INV_X1    g0707(.A(new_n684), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n355), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n368), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT106), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT37), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n909), .A2(new_n365), .ZN(new_n914));
  INV_X1    g0714(.A(new_n356), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n912), .B(new_n913), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n328), .A2(new_n355), .B1(KEYINPUT106), .B2(KEYINPUT37), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n912), .A2(new_n913), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n917), .A2(new_n365), .A3(new_n909), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n907), .B1(new_n911), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n368), .A2(new_n910), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n922), .A2(KEYINPUT38), .A3(new_n916), .A4(new_n919), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n906), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n362), .A2(new_n367), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(KEYINPUT107), .ZN(new_n927));
  INV_X1    g0727(.A(new_n637), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT107), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n362), .A2(new_n929), .A3(new_n367), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n920), .B1(new_n931), .B2(new_n910), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n923), .B1(new_n932), .B2(KEYINPUT38), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT39), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n921), .A2(new_n923), .A3(KEYINPUT39), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n295), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n687), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n937), .A2(new_n939), .B1(new_n928), .B2(new_n908), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n925), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n895), .B(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n836), .B1(new_n899), .B2(new_n901), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n740), .A2(new_n944), .A3(new_n924), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT40), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n933), .A2(new_n740), .A3(KEYINPUT40), .A4(new_n944), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT109), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n424), .A2(new_n740), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n951), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n952), .A2(G330), .A3(new_n953), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n943), .A2(new_n954), .B1(new_n205), .B2(new_n756), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(KEYINPUT110), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n943), .A2(new_n954), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n955), .A2(KEYINPUT110), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n891), .B1(new_n958), .B2(new_n959), .ZN(G367));
  NOR2_X1   g0760(.A1(new_n672), .A2(new_n687), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n647), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n660), .B2(new_n961), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n963), .A2(KEYINPUT111), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(KEYINPUT111), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n772), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n765), .A2(new_n234), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n775), .B1(new_n701), .B2(new_n556), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n845), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n773), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n271), .B1(new_n804), .B2(new_n861), .C1(new_n852), .C2(new_n812), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(G137), .B2(new_n802), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n798), .A2(G68), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n781), .A2(new_n247), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(G150), .B2(new_n790), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n786), .A2(G143), .B1(G58), .B2(new_n777), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n973), .A2(new_n974), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n335), .B1(new_n782), .B2(new_n804), .C1(new_n852), .C2(new_n849), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(G317), .B2(new_n802), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n777), .A2(G116), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT46), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n798), .A2(G107), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n850), .A2(new_n593), .B1(new_n609), .B2(new_n781), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(G311), .B2(new_n786), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n980), .A2(new_n982), .A3(new_n983), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n978), .A2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT47), .Z(new_n988));
  OAI211_X1 g0788(.A(new_n967), .B(new_n970), .C1(new_n971), .C2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n528), .A2(new_n686), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n717), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n529), .A2(new_n687), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n698), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(KEYINPUT42), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n717), .A2(new_n990), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n529), .B2(new_n687), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT42), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n996), .A2(new_n997), .A3(new_n698), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n529), .B1(new_n995), .B2(new_n489), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n687), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n994), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT43), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n966), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n964), .A2(KEYINPUT43), .A3(new_n965), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1001), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n993), .A2(KEYINPUT42), .B1(new_n999), .B2(new_n687), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1006), .A2(new_n1002), .A3(new_n966), .A4(new_n998), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT112), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n695), .A2(new_n996), .ZN(new_n1010));
  AND3_X1   g0810(.A1(new_n1009), .A2(KEYINPUT113), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(KEYINPUT113), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1012));
  AND2_X1   g0812(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n1011), .A2(new_n1012), .B1(new_n1008), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT113), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1013), .A2(new_n1008), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1009), .A2(KEYINPUT113), .A3(new_n1010), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1014), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n996), .A2(new_n699), .ZN(new_n1022));
  XOR2_X1   g0822(.A(KEYINPUT114), .B(KEYINPUT44), .Z(new_n1023));
  XNOR2_X1  g0823(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n996), .A2(new_n699), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT45), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1025), .A2(new_n696), .A3(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n695), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  AND2_X1   g0831(.A1(new_n692), .A2(KEYINPUT115), .ZN(new_n1032));
  MUX2_X1   g0832(.A(new_n493), .B(new_n694), .S(new_n697), .Z(new_n1033));
  OR2_X1    g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n692), .A2(KEYINPUT115), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1033), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n754), .B1(new_n1031), .B2(new_n1037), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n702), .B(KEYINPUT41), .Z(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n758), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n989), .B1(new_n1021), .B2(new_n1041), .ZN(G387));
  AOI21_X1  g0842(.A(new_n1037), .B1(new_n753), .B2(new_n742), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1037), .A2(new_n742), .A3(new_n753), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1044), .A2(new_n702), .A3(new_n1045), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n762), .A2(new_n705), .B1(new_n298), .B2(new_n701), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT116), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n471), .B1(new_n330), .B2(new_n247), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n311), .A2(G50), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT50), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AND2_X1   g0852(.A1(new_n705), .A2(KEYINPUT117), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n705), .A2(KEYINPUT117), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1052), .B1(new_n1051), .B2(new_n1050), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1055), .A2(KEYINPUT118), .A3(new_n765), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n231), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1056), .B1(new_n1057), .B2(new_n471), .ZN(new_n1058));
  AOI21_X1  g0858(.A(KEYINPUT118), .B1(new_n1055), .B2(new_n765), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1048), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n845), .B1(new_n1060), .B2(new_n774), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n335), .B1(new_n805), .B2(G68), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(new_n609), .B2(new_n781), .C1(new_n811), .C2(new_n377), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n797), .A2(new_n309), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n351), .A2(new_n852), .B1(new_n850), .B2(new_n861), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n786), .A2(G159), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n247), .B2(new_n778), .ZN(new_n1067));
  NOR4_X1   g0867(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .A4(new_n1067), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G317), .A2(new_n790), .B1(new_n805), .B2(new_n594), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1069), .A2(KEYINPUT119), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(KEYINPUT119), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(G311), .A2(new_n807), .B1(new_n786), .B2(G322), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT48), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n798), .A2(G283), .B1(G294), .B2(new_n777), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT49), .Z(new_n1079));
  OR2_X1    g0879(.A1(new_n1079), .A2(KEYINPUT120), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n335), .B1(new_n611), .B2(new_n781), .C1(new_n811), .C2(new_n788), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n1079), .B2(KEYINPUT120), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1068), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1061), .B1(new_n1083), .B2(new_n971), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n694), .B2(new_n772), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1037), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1085), .B1(new_n1086), .B2(new_n758), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1046), .A2(new_n1087), .ZN(G393));
  INV_X1    g0888(.A(KEYINPUT121), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1044), .A2(new_n1089), .A3(new_n1031), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1031), .ZN(new_n1091));
  OAI21_X1  g0891(.A(KEYINPUT121), .B1(new_n1043), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n703), .B1(new_n1043), .B2(new_n1091), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1091), .A2(new_n758), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n239), .A2(new_n766), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n774), .B1(new_n609), .B2(new_n209), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n759), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n271), .B1(new_n311), .B2(new_n804), .C1(new_n852), .C2(new_n861), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n854), .B(new_n1100), .C1(G68), .C2(new_n777), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n790), .A2(G159), .B1(new_n786), .B2(G150), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT51), .Z(new_n1103));
  NAND2_X1  g0903(.A1(new_n798), .A2(G77), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n802), .A2(G143), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1101), .A2(new_n1103), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n335), .B1(new_n849), .B2(new_n804), .C1(new_n852), .C2(new_n593), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n818), .B(new_n1107), .C1(G283), .C2(new_n777), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n802), .A2(G322), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1108), .B(new_n1109), .C1(new_n611), .C2(new_n797), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n790), .A2(G311), .B1(new_n786), .B2(G317), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT52), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1106), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1099), .B1(new_n1113), .B2(new_n773), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n996), .B2(new_n825), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1096), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1095), .A2(new_n1117), .ZN(G390));
  NOR2_X1   g0918(.A1(new_n645), .A2(new_n741), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n644), .B(new_n1120), .C1(new_n892), .C2(new_n894), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n741), .A2(new_n836), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n902), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n903), .B1(new_n741), .B2(new_n836), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n842), .A2(new_n905), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n719), .A2(new_n687), .A3(new_n841), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n905), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n1132), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1133));
  OR2_X1    g0933(.A1(new_n1129), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1124), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n937), .ZN(new_n1136));
  NOR3_X1   g0936(.A1(new_n679), .A2(new_n686), .A3(new_n840), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n902), .B1(new_n1137), .B2(new_n904), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1136), .B1(new_n1138), .B2(new_n939), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n933), .A2(new_n939), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n1131), .B2(new_n902), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1135), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n939), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n937), .B1(new_n906), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1141), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1144), .A2(new_n1124), .A3(new_n1145), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1122), .A2(new_n1134), .A3(new_n1142), .A4(new_n1146), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1144), .A2(new_n1124), .A3(new_n1145), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1124), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1129), .A2(new_n1133), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n1148), .A2(new_n1149), .B1(new_n1150), .B2(new_n1121), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1147), .A2(new_n1151), .A3(new_n702), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n758), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n845), .B1(new_n351), .B2(new_n873), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n777), .A2(G150), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT53), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT54), .B(G143), .ZN(new_n1158));
  INV_X1    g0958(.A(G137), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n271), .B1(new_n804), .B2(new_n1158), .C1(new_n852), .C2(new_n1159), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1157), .B(new_n1160), .C1(G125), .C2(new_n802), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n786), .A2(G128), .ZN(new_n1162));
  INV_X1    g0962(.A(G132), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1162), .B1(new_n861), .B2(new_n781), .C1(new_n850), .C2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G159), .B2(new_n798), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n335), .B1(new_n609), .B2(new_n804), .C1(new_n852), .C2(new_n298), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n811), .A2(new_n849), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n611), .A2(new_n850), .B1(new_n787), .B2(new_n782), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n778), .A2(new_n544), .B1(new_n781), .B2(new_n330), .ZN(new_n1169));
  NOR4_X1   g0969(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n1161), .A2(new_n1165), .B1(new_n1170), .B2(new_n1104), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1155), .B1(new_n971), .B2(new_n1171), .C1(new_n1136), .C2(new_n771), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1152), .A2(new_n1154), .A3(new_n1172), .ZN(G378));
  XOR2_X1   g0973(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1174));
  NAND2_X1  g0974(.A1(new_n410), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1174), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n402), .A2(new_n405), .A3(new_n409), .A4(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n386), .A2(new_n908), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT123), .Z(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1178), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1175), .A2(new_n1180), .A3(new_n1177), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n947), .A2(G330), .A3(new_n948), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1184), .A2(new_n947), .A3(G330), .A4(new_n948), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  AND3_X1   g0989(.A1(new_n1127), .A2(new_n924), .A3(new_n902), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1189), .B1(new_n1190), .B2(new_n940), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n925), .A2(new_n941), .A3(new_n1188), .A4(new_n1187), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1191), .A2(KEYINPUT124), .A3(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT124), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n942), .A2(new_n1194), .A3(new_n1189), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1185), .A2(new_n770), .ZN(new_n1197));
  NOR3_X1   g0997(.A1(new_n773), .A2(G50), .A3(new_n770), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n852), .A2(new_n1163), .B1(new_n1159), .B2(new_n804), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1158), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1199), .B1(new_n777), .B2(new_n1200), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n790), .A2(G128), .B1(new_n786), .B2(G125), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(new_n377), .C2(new_n797), .ZN(new_n1203));
  OR2_X1    g1003(.A1(new_n1203), .A2(KEYINPUT59), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(KEYINPUT59), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n266), .B(new_n457), .C1(new_n781), .C2(new_n812), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n802), .B2(G124), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1204), .A2(new_n1205), .A3(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n271), .A2(G41), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1209), .B1(new_n309), .B2(new_n804), .C1(new_n852), .C2(new_n609), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G283), .B2(new_n802), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n786), .A2(G116), .B1(G77), .B2(new_n777), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n781), .A2(new_n338), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G107), .B2(new_n790), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1211), .A2(new_n974), .A3(new_n1212), .A4(new_n1214), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1209), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1218), .B(new_n861), .C1(G33), .C2(G41), .ZN(new_n1219));
  OR2_X1    g1019(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1208), .A2(new_n1217), .A3(new_n1219), .A4(new_n1220), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n845), .B(new_n1198), .C1(new_n1221), .C2(new_n773), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1196), .A2(new_n758), .B1(new_n1197), .B2(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1150), .A2(new_n1121), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1121), .B1(new_n1153), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT57), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n702), .B1(new_n1225), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1142), .A2(new_n1146), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1122), .B1(new_n1230), .B2(new_n1150), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT57), .B1(new_n1231), .B2(new_n1196), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1223), .B1(new_n1229), .B2(new_n1232), .ZN(G375));
  NAND2_X1  g1033(.A1(new_n1122), .A2(new_n1134), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1150), .A2(new_n1121), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1234), .A2(new_n1040), .A3(new_n1235), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n1163), .A2(new_n787), .B1(new_n850), .B2(new_n1159), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n1213), .B(new_n1237), .C1(G159), .C2(new_n777), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n271), .B1(new_n804), .B2(new_n377), .C1(new_n852), .C2(new_n1158), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(G128), .B2(new_n802), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1238), .B(new_n1240), .C1(new_n861), .C2(new_n797), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n782), .A2(new_n850), .B1(new_n787), .B2(new_n849), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n975), .B(new_n1242), .C1(G97), .C2(new_n777), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n335), .B1(new_n804), .B2(new_n298), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G116), .B2(new_n807), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1243), .B(new_n1245), .C1(new_n779), .C2(new_n811), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1241), .B1(new_n1246), .B2(new_n1064), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n773), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n845), .B1(new_n330), .B2(new_n873), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n903), .B2(new_n770), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n1134), .B2(new_n758), .ZN(new_n1252));
  AND2_X1   g1052(.A1(new_n1236), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(G381));
  NAND3_X1  g1054(.A1(new_n1046), .A2(new_n827), .A3(new_n1087), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(G390), .A2(new_n1255), .A3(G384), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(G378), .A2(G387), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n1256), .A2(new_n1253), .A3(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(G375), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1258), .A2(KEYINPUT125), .A3(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT125), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1261));
  OR2_X1    g1061(.A1(new_n1260), .A2(new_n1261), .ZN(G407));
  OAI21_X1  g1062(.A(new_n1172), .B1(new_n1230), .B2(new_n757), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n703), .B1(new_n1234), .B2(new_n1230), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1263), .B1(new_n1264), .B2(new_n1147), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n685), .ZN(new_n1266));
  OAI221_X1 g1066(.A(G213), .B1(G375), .B2(new_n1266), .C1(new_n1260), .C2(new_n1261), .ZN(G409));
  NAND2_X1  g1067(.A1(G393), .A2(G396), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1255), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1095), .A2(G387), .A3(new_n1117), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(G387), .B1(new_n1095), .B2(new_n1117), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1269), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  OR2_X1    g1073(.A1(new_n1021), .A2(new_n1041), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1094), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1275), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1274), .B(new_n989), .C1(new_n1276), .C2(new_n1116), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1277), .A2(new_n1255), .A3(new_n1268), .A4(new_n1270), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1273), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(G213), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1280), .A2(G343), .ZN(new_n1281));
  OAI211_X1 g1081(.A(G378), .B(new_n1223), .C1(new_n1229), .C2(new_n1232), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1283));
  NOR3_X1   g1083(.A1(new_n1225), .A2(new_n1039), .A3(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n757), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1197), .A2(new_n1222), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  OR2_X1    g1087(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1265), .B1(new_n1284), .B2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1281), .B1(new_n1282), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT126), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT60), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1291), .B1(new_n1235), .B2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n703), .B1(new_n1122), .B2(new_n1134), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1150), .A2(new_n1121), .A3(KEYINPUT126), .A4(KEYINPUT60), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1235), .A2(new_n1292), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1293), .A2(new_n1294), .A3(new_n1295), .A4(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1252), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(G384), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1297), .A2(new_n881), .A3(new_n1252), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1290), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT63), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1279), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1281), .A2(G2897), .ZN(new_n1305));
  AND3_X1   g1105(.A1(new_n1297), .A2(new_n881), .A3(new_n1252), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n881), .B1(new_n1297), .B2(new_n1252), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1305), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1305), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1299), .A2(new_n1300), .A3(new_n1309), .ZN(new_n1310));
  AND2_X1   g1110(.A1(new_n1308), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1290), .ZN(new_n1312));
  AOI21_X1  g1112(.A(KEYINPUT61), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1290), .A2(KEYINPUT63), .A3(new_n1301), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1304), .A2(new_n1313), .A3(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT61), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1308), .A2(new_n1310), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1316), .B1(new_n1317), .B2(new_n1290), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT62), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1282), .A2(new_n1289), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1281), .ZN(new_n1321));
  AND4_X1   g1121(.A1(new_n1319), .A2(new_n1320), .A3(new_n1321), .A4(new_n1301), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1319), .B1(new_n1290), .B2(new_n1301), .ZN(new_n1323));
  NOR3_X1   g1123(.A1(new_n1318), .A2(new_n1322), .A3(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1279), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1315), .B1(new_n1324), .B2(new_n1325), .ZN(G405));
  INV_X1    g1126(.A(KEYINPUT127), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1282), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1226), .B1(new_n1225), .B2(new_n1283), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n703), .B1(new_n1231), .B2(new_n1227), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(G378), .B1(new_n1331), .B2(new_n1223), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1327), .B1(new_n1328), .B2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1301), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(G375), .A2(new_n1265), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1335), .A2(KEYINPUT127), .A3(new_n1282), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1333), .A2(new_n1334), .A3(new_n1336), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1335), .A2(new_n1301), .A3(KEYINPUT127), .A4(new_n1282), .ZN(new_n1338));
  AND3_X1   g1138(.A1(new_n1337), .A2(new_n1325), .A3(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1325), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1339), .A2(new_n1340), .ZN(G402));
endmodule


