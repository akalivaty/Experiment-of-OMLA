//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 0 0 0 1 1 1 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 1 0 1 1 1 1 1 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1232, new_n1233, new_n1234, new_n1235, new_n1237,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G13), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT0), .Z(new_n214));
  AOI22_X1  g0014(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G97), .A2(G257), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G68), .A2(G238), .ZN(new_n217));
  NAND3_X1  g0017(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n219));
  INV_X1    g0019(.A(G116), .ZN(new_n220));
  INV_X1    g0020(.A(G270), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AOI211_X1 g0022(.A(new_n218), .B(new_n222), .C1(G58), .C2(G232), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n223), .A2(new_n209), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT1), .Z(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n208), .ZN(new_n227));
  OAI21_X1  g0027(.A(G50), .B1(G58), .B2(G68), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n214), .B(new_n225), .C1(new_n227), .C2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT2), .ZN(new_n234));
  INV_X1    g0034(.A(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G264), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n221), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G97), .B(G107), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G87), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(new_n220), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  XNOR2_X1  g0047(.A(KEYINPUT3), .B(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n248), .A2(G257), .A3(new_n249), .ZN(new_n250));
  AND2_X1   g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G303), .ZN(new_n254));
  OAI211_X1 g0054(.A(G264), .B(G1698), .C1(new_n251), .C2(new_n252), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n250), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  OAI211_X1 g0058(.A(G1), .B(G13), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT5), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n207), .B(G45), .C1(new_n262), .C2(G41), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n258), .A2(KEYINPUT5), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(new_n260), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G270), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  INV_X1    g0068(.A(G274), .ZN(new_n269));
  NOR3_X1   g0069(.A1(new_n268), .A2(new_n269), .A3(G1), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n262), .A2(G41), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT79), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n272), .B1(new_n262), .B2(G41), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n258), .A2(KEYINPUT79), .A3(KEYINPUT5), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n270), .A2(new_n271), .A3(new_n273), .A4(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n261), .A2(new_n267), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G200), .ZN(new_n277));
  NOR3_X1   g0077(.A1(new_n210), .A2(new_n208), .A3(G1), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n226), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n207), .A2(G33), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n279), .A2(G116), .A3(new_n282), .A4(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n278), .A2(new_n220), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n280), .A2(new_n226), .B1(G20), .B2(new_n220), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G283), .ZN(new_n287));
  INV_X1    g0087(.A(G97), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n287), .B(new_n208), .C1(G33), .C2(new_n288), .ZN(new_n289));
  AND3_X1   g0089(.A1(new_n286), .A2(KEYINPUT20), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(KEYINPUT20), .B1(new_n286), .B2(new_n289), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n284), .B(new_n285), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G190), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n277), .B(new_n293), .C1(new_n294), .C2(new_n276), .ZN(new_n295));
  INV_X1    g0095(.A(G179), .ZN(new_n296));
  NOR3_X1   g0096(.A1(new_n276), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT21), .ZN(new_n299));
  INV_X1    g0099(.A(G169), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n256), .A2(new_n260), .B1(new_n266), .B2(G270), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n300), .B1(new_n301), .B2(new_n275), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n299), .B1(new_n302), .B2(new_n292), .ZN(new_n303));
  AND4_X1   g0103(.A1(new_n299), .A2(new_n276), .A3(new_n292), .A4(G169), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n295), .B(new_n298), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT86), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n276), .A2(new_n292), .A3(G169), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT21), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n302), .A2(new_n299), .A3(new_n292), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n297), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n311), .A2(KEYINPUT86), .A3(new_n295), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n278), .A2(new_n202), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n281), .B1(new_n207), .B2(G20), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G50), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT8), .B(G58), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n208), .A2(G33), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(G20), .A2(G33), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G150), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI211_X1 g0123(.A(new_n319), .B(new_n323), .C1(new_n204), .C2(G20), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n314), .B(new_n316), .C1(new_n324), .C2(new_n282), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT9), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n328), .A2(new_n269), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n259), .A2(new_n328), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n330), .B1(new_n331), .B2(new_n235), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n332), .B(KEYINPUT65), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n253), .A2(new_n249), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G223), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n248), .A2(new_n249), .ZN(new_n337));
  INV_X1    g0137(.A(G222), .ZN(new_n338));
  INV_X1    g0138(.A(G77), .ZN(new_n339));
  OAI22_X1  g0139(.A1(new_n337), .A2(new_n338), .B1(new_n339), .B2(new_n248), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n260), .B1(new_n336), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n333), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G200), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n323), .B1(new_n204), .B2(G20), .ZN(new_n344));
  INV_X1    g0144(.A(new_n319), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n281), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n347), .A2(KEYINPUT9), .A3(new_n314), .A4(new_n316), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n333), .A2(G190), .A3(new_n341), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n327), .A2(new_n343), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT10), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT71), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n350), .A2(KEYINPUT71), .A3(KEYINPUT10), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n327), .A2(new_n348), .A3(KEYINPUT70), .ZN(new_n355));
  AND3_X1   g0155(.A1(new_n355), .A2(new_n343), .A3(new_n349), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n327), .A2(new_n348), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT70), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT10), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n353), .A2(new_n354), .B1(new_n356), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n342), .A2(G179), .ZN(new_n361));
  XNOR2_X1  g0161(.A(new_n361), .B(KEYINPUT66), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n342), .A2(new_n300), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n362), .A2(new_n363), .A3(new_n325), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  OAI211_X1 g0165(.A(G232), .B(G1698), .C1(new_n251), .C2(new_n252), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT72), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT72), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n248), .A2(new_n368), .A3(G232), .A4(G1698), .ZN(new_n369));
  NAND2_X1  g0169(.A1(G33), .A2(G97), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n248), .A2(G226), .A3(new_n249), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n367), .A2(new_n369), .A3(new_n370), .A4(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n260), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT73), .ZN(new_n374));
  INV_X1    g0174(.A(new_n331), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G238), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT73), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n372), .A2(new_n377), .A3(new_n260), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n374), .A2(new_n376), .A3(new_n378), .A4(new_n330), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT13), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n329), .B1(new_n373), .B2(KEYINPUT73), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT13), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n381), .A2(new_n382), .A3(new_n376), .A4(new_n378), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n384), .A2(new_n294), .ZN(new_n385));
  INV_X1    g0185(.A(G68), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(G20), .ZN(new_n387));
  OAI221_X1 g0187(.A(new_n387), .B1(new_n318), .B2(new_n339), .C1(new_n321), .C2(new_n202), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n388), .A2(KEYINPUT11), .A3(new_n281), .ZN(new_n389));
  INV_X1    g0189(.A(new_n315), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n389), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n278), .A2(new_n386), .ZN(new_n392));
  XOR2_X1   g0192(.A(new_n392), .B(KEYINPUT12), .Z(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT11), .B1(new_n388), .B2(new_n281), .ZN(new_n394));
  NOR3_X1   g0194(.A1(new_n391), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G200), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n397), .B1(new_n380), .B2(new_n383), .ZN(new_n398));
  NOR3_X1   g0198(.A1(new_n385), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  NOR3_X1   g0199(.A1(new_n360), .A2(new_n365), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n334), .A2(G238), .ZN(new_n401));
  XNOR2_X1  g0201(.A(KEYINPUT67), .B(G107), .ZN(new_n402));
  OAI221_X1 g0202(.A(new_n401), .B1(new_n232), .B2(new_n337), .C1(new_n248), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n260), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n375), .A2(G244), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(new_n330), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT68), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT68), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n404), .A2(new_n408), .A3(new_n330), .A4(new_n405), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n296), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n279), .A2(G77), .ZN(new_n412));
  OAI22_X1  g0212(.A1(new_n317), .A2(new_n321), .B1(new_n208), .B2(new_n339), .ZN(new_n413));
  XNOR2_X1  g0213(.A(new_n413), .B(KEYINPUT69), .ZN(new_n414));
  XOR2_X1   g0214(.A(KEYINPUT15), .B(G87), .Z(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n414), .B1(new_n416), .B2(new_n318), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n412), .B1(new_n417), .B2(new_n281), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n339), .B2(new_n390), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n411), .B(new_n419), .C1(G169), .C2(new_n410), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n384), .A2(G169), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT14), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n380), .A2(G179), .A3(new_n383), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT14), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n384), .A2(new_n425), .A3(G169), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n423), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n421), .B1(new_n427), .B2(new_n396), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n419), .B1(new_n410), .B2(G190), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n407), .A2(G200), .A3(new_n409), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n317), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n432), .A2(new_n278), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n433), .B1(new_n390), .B2(new_n432), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n248), .A2(G226), .A3(G1698), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n248), .A2(G223), .A3(new_n249), .ZN(new_n437));
  NAND2_X1  g0237(.A1(G33), .A2(G87), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n329), .B1(new_n439), .B2(new_n260), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT76), .B1(new_n331), .B2(new_n232), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT76), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n259), .A2(new_n442), .A3(G232), .A4(new_n328), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n440), .A2(G190), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT7), .B1(new_n253), .B2(new_n208), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT3), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n257), .ZN(new_n448));
  NAND2_X1  g0248(.A1(KEYINPUT3), .A2(G33), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n448), .A2(KEYINPUT7), .A3(new_n208), .A4(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(G68), .B1(new_n446), .B2(new_n451), .ZN(new_n452));
  AND2_X1   g0252(.A1(G58), .A2(G68), .ZN(new_n453));
  OAI21_X1  g0253(.A(G20), .B1(new_n453), .B2(new_n201), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n320), .A2(G159), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n452), .A2(KEYINPUT16), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT74), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n448), .A2(new_n208), .A3(new_n449), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT7), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n450), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n456), .B1(new_n464), .B2(G68), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n465), .A2(KEYINPUT74), .A3(KEYINPUT16), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n460), .A2(new_n281), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n463), .A2(KEYINPUT75), .A3(new_n450), .ZN(new_n468));
  OR2_X1    g0268(.A1(new_n450), .A2(KEYINPUT75), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n468), .A2(G68), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT16), .B1(new_n470), .B2(new_n457), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n435), .B(new_n445), .C1(new_n467), .C2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT77), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n439), .A2(new_n260), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n475), .A2(new_n444), .A3(new_n330), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G200), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n473), .A2(new_n474), .A3(KEYINPUT17), .A4(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT17), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n470), .A2(new_n457), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT16), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n482), .A2(new_n281), .A3(new_n460), .A4(new_n466), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n483), .A2(new_n477), .A3(new_n435), .A4(new_n445), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n479), .B1(new_n484), .B2(KEYINPUT77), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n478), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n435), .B1(new_n467), .B2(new_n471), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n476), .A2(new_n296), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n300), .B1(new_n440), .B2(new_n444), .ZN(new_n489));
  OR2_X1    g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n487), .A2(KEYINPUT18), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(KEYINPUT18), .B1(new_n487), .B2(new_n490), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n486), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n400), .A2(new_n428), .A3(new_n431), .A4(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n278), .A2(new_n288), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n279), .A2(new_n282), .A3(new_n283), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n497), .B1(new_n498), .B2(new_n288), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n288), .A2(G107), .ZN(new_n500));
  MUX2_X1   g0300(.A(new_n244), .B(new_n500), .S(KEYINPUT6), .Z(new_n501));
  AOI22_X1  g0301(.A1(new_n501), .A2(G20), .B1(G77), .B2(new_n320), .ZN(new_n502));
  INV_X1    g0302(.A(new_n402), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n468), .A2(new_n503), .A3(new_n469), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n499), .B1(new_n505), .B2(new_n281), .ZN(new_n506));
  OAI211_X1 g0306(.A(G244), .B(new_n249), .C1(new_n251), .C2(new_n252), .ZN(new_n507));
  XNOR2_X1  g0307(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OR2_X1    g0309(.A1(KEYINPUT78), .A2(KEYINPUT4), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n248), .A2(G244), .A3(new_n249), .A4(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n248), .A2(G250), .A3(G1698), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n509), .A2(new_n511), .A3(new_n287), .A4(new_n512), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n513), .A2(new_n260), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n259), .B(G257), .C1(new_n263), .C2(new_n264), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n275), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT80), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT80), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n515), .A2(new_n275), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(G200), .B1(new_n514), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n516), .B1(new_n513), .B2(new_n260), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G190), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n506), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT81), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n513), .A2(new_n260), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n527), .A2(new_n296), .A3(new_n517), .A4(new_n519), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n282), .B1(new_n502), .B2(new_n504), .ZN(new_n529));
  OAI221_X1 g0329(.A(new_n528), .B1(G169), .B2(new_n522), .C1(new_n529), .C2(new_n499), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n506), .A2(new_n521), .A3(KEYINPUT81), .A4(new_n523), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n526), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n208), .B(G87), .C1(new_n251), .C2(new_n252), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT22), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT22), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n248), .A2(new_n535), .A3(new_n208), .A4(G87), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n402), .A2(G20), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT23), .ZN(new_n539));
  INV_X1    g0339(.A(G107), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n539), .A2(new_n540), .A3(G20), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT87), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n539), .A2(new_n540), .A3(KEYINPUT87), .A4(G20), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n538), .A2(KEYINPUT23), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n208), .A2(G33), .A3(G116), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n537), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT24), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n537), .A2(new_n545), .A3(KEYINPUT24), .A4(new_n546), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n549), .A2(new_n281), .A3(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n279), .A2(G107), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT88), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT25), .ZN(new_n554));
  OAI22_X1  g0354(.A1(new_n540), .A2(new_n498), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  XNOR2_X1  g0355(.A(KEYINPUT88), .B(KEYINPUT25), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n555), .B1(new_n552), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n551), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(G257), .B(G1698), .C1(new_n251), .C2(new_n252), .ZN(new_n559));
  OAI211_X1 g0359(.A(G250), .B(new_n249), .C1(new_n251), .C2(new_n252), .ZN(new_n560));
  NAND2_X1  g0360(.A1(G33), .A2(G294), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT89), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT89), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n559), .A2(new_n560), .A3(new_n564), .A4(new_n561), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n563), .A2(new_n260), .A3(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n259), .B(G264), .C1(new_n263), .C2(new_n264), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n567), .A2(new_n275), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT90), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n566), .A2(KEYINPUT90), .A3(new_n568), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(new_n294), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n569), .A2(new_n397), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n558), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n532), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT85), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n248), .A2(G244), .A3(G1698), .ZN(new_n578));
  NAND2_X1  g0378(.A1(G33), .A2(G116), .ZN(new_n579));
  OAI211_X1 g0379(.A(G238), .B(new_n249), .C1(new_n251), .C2(new_n252), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n260), .ZN(new_n582));
  INV_X1    g0382(.A(new_n270), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT82), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n268), .B2(G1), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n207), .A2(KEYINPUT82), .A3(G45), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n259), .A2(new_n585), .A3(G250), .A4(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n582), .A2(new_n583), .A3(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n577), .B1(new_n588), .B2(new_n294), .ZN(new_n589));
  INV_X1    g0389(.A(new_n587), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n590), .B1(new_n581), .B2(new_n260), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n591), .A2(KEYINPUT85), .A3(G190), .A4(new_n583), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n588), .A2(G200), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n279), .A2(new_n415), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT84), .ZN(new_n596));
  AND2_X1   g0396(.A1(KEYINPUT83), .A2(KEYINPUT19), .ZN(new_n597));
  NOR2_X1   g0397(.A1(KEYINPUT83), .A2(KEYINPUT19), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n370), .ZN(new_n600));
  AOI21_X1  g0400(.A(G20), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(G87), .ZN(new_n602));
  AND2_X1   g0402(.A1(KEYINPUT67), .A2(G107), .ZN(new_n603));
  NOR2_X1   g0403(.A1(KEYINPUT67), .A2(G107), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n602), .B(new_n288), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n596), .B1(new_n601), .B2(new_n606), .ZN(new_n607));
  XNOR2_X1  g0407(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n208), .B1(new_n608), .B2(new_n370), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n609), .A2(KEYINPUT84), .A3(new_n605), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n248), .A2(new_n208), .A3(G68), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n608), .B1(new_n288), .B2(new_n318), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n607), .A2(new_n610), .A3(new_n611), .A4(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n595), .B1(new_n613), .B2(new_n281), .ZN(new_n614));
  INV_X1    g0414(.A(new_n498), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G87), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n593), .A2(new_n594), .A3(new_n614), .A4(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n415), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n588), .A2(new_n300), .ZN(new_n620));
  AOI211_X1 g0420(.A(new_n270), .B(new_n590), .C1(new_n260), .C2(new_n581), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n296), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n619), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n617), .A2(new_n623), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n551), .A2(new_n557), .ZN(new_n625));
  INV_X1    g0425(.A(new_n572), .ZN(new_n626));
  AOI21_X1  g0426(.A(KEYINPUT90), .B1(new_n566), .B2(new_n568), .ZN(new_n627));
  OAI21_X1  g0427(.A(G169), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n569), .A2(new_n296), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n625), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n624), .A2(new_n631), .ZN(new_n632));
  AND4_X1   g0432(.A1(new_n313), .A2(new_n496), .A3(new_n576), .A4(new_n632), .ZN(G372));
  INV_X1    g0433(.A(KEYINPUT94), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n491), .B2(new_n492), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT18), .ZN(new_n636));
  AOI21_X1  g0436(.A(KEYINPUT74), .B1(new_n465), .B2(KEYINPUT16), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n386), .B1(new_n463), .B2(new_n450), .ZN(new_n638));
  NOR4_X1   g0438(.A1(new_n638), .A2(new_n459), .A3(new_n481), .A4(new_n456), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n637), .A2(new_n639), .A3(new_n282), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n434), .B1(new_n640), .B2(new_n482), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n488), .A2(new_n489), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n636), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n487), .A2(new_n490), .A3(KEYINPUT18), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(KEYINPUT94), .A3(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n635), .A2(new_n645), .ZN(new_n646));
  OR3_X1    g0446(.A1(new_n385), .A2(new_n396), .A3(new_n398), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n425), .B1(new_n384), .B2(G169), .ZN(new_n648));
  AOI211_X1 g0448(.A(KEYINPUT14), .B(new_n300), .C1(new_n380), .C2(new_n383), .ZN(new_n649));
  INV_X1    g0449(.A(new_n424), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n651), .A2(new_n395), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n647), .B1(new_n652), .B2(new_n421), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n646), .B1(new_n653), .B2(new_n486), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n356), .A2(new_n359), .ZN(new_n655));
  INV_X1    g0455(.A(new_n354), .ZN(new_n656));
  AOI21_X1  g0456(.A(KEYINPUT71), .B1(new_n350), .B2(KEYINPUT10), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n365), .B1(new_n654), .B2(new_n658), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n626), .A2(new_n627), .A3(G190), .ZN(new_n660));
  INV_X1    g0460(.A(new_n574), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n625), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n662), .A2(new_n530), .A3(new_n526), .A4(new_n531), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n614), .A2(new_n594), .A3(new_n616), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT91), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n614), .A2(KEYINPUT91), .A3(new_n594), .A4(new_n616), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(new_n593), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n623), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT92), .B1(new_n663), .B2(new_n669), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n619), .A2(new_n620), .A3(new_n622), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n667), .A2(new_n593), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n671), .B1(new_n672), .B2(new_n666), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n526), .A2(new_n530), .A3(new_n531), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT92), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n673), .A2(new_n674), .A3(new_n675), .A4(new_n662), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n311), .A2(KEYINPUT93), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n300), .B1(new_n571), .B2(new_n572), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n558), .B1(new_n678), .B2(new_n629), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n311), .A2(KEYINPUT93), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n677), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n670), .A2(new_n676), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(KEYINPUT26), .B1(new_n624), .B2(new_n530), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT26), .ZN(new_n684));
  INV_X1    g0484(.A(new_n530), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n668), .A2(new_n684), .A3(new_n685), .A4(new_n623), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n683), .A2(new_n686), .A3(new_n623), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n682), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n496), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n659), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT95), .ZN(G369));
  INV_X1    g0491(.A(G330), .ZN(new_n692));
  XOR2_X1   g0492(.A(KEYINPUT96), .B(KEYINPUT27), .Z(new_n693));
  NOR3_X1   g0493(.A1(new_n210), .A2(G1), .A3(G20), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G213), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G343), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(new_n293), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n701), .B1(new_n307), .B2(new_n312), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n677), .A2(new_n680), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n701), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n692), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n625), .A2(new_n700), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n679), .B1(new_n707), .B2(new_n575), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n631), .A2(new_n700), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n711), .A2(KEYINPUT97), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(KEYINPUT97), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n311), .A2(new_n699), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n710), .A2(new_n715), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n716), .A2(new_n709), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n714), .A2(new_n717), .ZN(G399));
  NOR2_X1   g0518(.A1(new_n211), .A2(G41), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G1), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n606), .A2(new_n220), .ZN(new_n722));
  OAI22_X1  g0522(.A1(new_n721), .A2(new_n722), .B1(new_n228), .B2(new_n720), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT28), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n699), .B1(new_n682), .B2(new_n687), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(KEYINPUT29), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n576), .A2(new_n313), .A3(new_n632), .A4(new_n700), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT31), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n301), .A2(new_n583), .A3(new_n591), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n629), .A2(new_n730), .A3(new_n522), .A4(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n621), .A2(new_n301), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n522), .A2(G179), .A3(new_n566), .A4(new_n568), .ZN(new_n734));
  OAI21_X1  g0534(.A(KEYINPUT30), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n621), .A2(G179), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n527), .A2(new_n517), .A3(new_n519), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n737), .A2(new_n276), .A3(new_n569), .A4(new_n738), .ZN(new_n739));
  AND3_X1   g0539(.A1(new_n736), .A2(KEYINPUT98), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(KEYINPUT98), .B1(new_n736), .B2(new_n739), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n740), .A2(new_n741), .A3(new_n700), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n729), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT31), .ZN(new_n745));
  AOI211_X1 g0545(.A(new_n745), .B(new_n700), .C1(new_n736), .C2(new_n739), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n692), .B1(new_n744), .B2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT29), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n679), .A2(new_n311), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n673), .A2(new_n674), .A3(new_n662), .A4(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(KEYINPUT26), .B1(new_n669), .B2(new_n530), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n617), .A2(new_n685), .A3(new_n684), .A4(new_n623), .ZN(new_n753));
  AND2_X1   g0553(.A1(new_n753), .A2(new_n623), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n751), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n749), .B1(new_n755), .B2(new_n700), .ZN(new_n756));
  NOR3_X1   g0556(.A1(new_n727), .A2(new_n748), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n724), .B1(new_n757), .B2(G1), .ZN(G364));
  NOR2_X1   g0558(.A1(new_n210), .A2(G20), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n207), .B1(new_n759), .B2(G45), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n719), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n706), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n703), .A2(new_n705), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n763), .B1(G330), .B2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n762), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n208), .A2(new_n296), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n768), .A2(new_n294), .A3(G200), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n248), .B1(new_n769), .B2(G322), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n294), .A2(G179), .A3(G200), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n208), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n294), .A2(new_n397), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n767), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n773), .A2(G294), .B1(new_n776), .B2(G326), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n770), .A2(new_n777), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n768), .A2(new_n397), .A3(G190), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n779), .A2(KEYINPUT101), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(KEYINPUT101), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(KEYINPUT33), .B(G317), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n778), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n768), .A2(G190), .A3(G200), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G311), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n774), .A2(G20), .A3(new_n296), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n788), .A2(KEYINPUT100), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(KEYINPUT100), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G303), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n294), .A2(G20), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT99), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(new_n296), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n397), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(G200), .ZN(new_n798));
  AOI22_X1  g0598(.A1(G283), .A2(new_n797), .B1(new_n798), .B2(G329), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n785), .A2(new_n787), .A3(new_n793), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n798), .A2(G159), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT32), .Z(new_n802));
  INV_X1    g0602(.A(new_n797), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n803), .A2(new_n540), .B1(new_n791), .B2(new_n602), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n773), .A2(G97), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(new_n202), .B2(new_n775), .ZN(new_n806));
  INV_X1    g0606(.A(new_n769), .ZN(new_n807));
  INV_X1    g0607(.A(G58), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n248), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n804), .A2(new_n806), .A3(new_n809), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n802), .B(new_n810), .C1(new_n386), .C2(new_n782), .ZN(new_n811));
  INV_X1    g0611(.A(new_n786), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n339), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n800), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n226), .B1(G20), .B2(new_n300), .ZN(new_n815));
  NOR2_X1   g0615(.A1(G13), .A2(G33), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(G20), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(new_n815), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n243), .A2(G45), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n211), .A2(new_n248), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n820), .B(new_n821), .C1(G45), .C2(new_n228), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n211), .A2(new_n253), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(G355), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n822), .B(new_n824), .C1(G116), .C2(new_n212), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n814), .A2(new_n815), .B1(new_n819), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n818), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n826), .B1(new_n764), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n765), .B1(new_n766), .B2(new_n828), .ZN(G396));
  NOR2_X1   g0629(.A1(new_n420), .A2(new_n699), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n419), .A2(new_n699), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n431), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n420), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n726), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n830), .B1(new_n420), .B2(new_n833), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n688), .A2(new_n700), .A3(new_n837), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n839), .A2(new_n748), .ZN(new_n840));
  OR2_X1    g0640(.A1(new_n840), .A2(KEYINPUT103), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n839), .A2(KEYINPUT103), .A3(new_n748), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n839), .A2(new_n748), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n841), .A2(new_n766), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n786), .A2(G159), .B1(new_n776), .B2(G137), .ZN(new_n845));
  INV_X1    g0645(.A(G143), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n845), .B1(new_n846), .B2(new_n807), .C1(new_n782), .C2(new_n322), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT34), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n797), .A2(G68), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n202), .B2(new_n791), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n253), .B(new_n850), .C1(G132), .C2(new_n798), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n848), .B(new_n851), .C1(new_n808), .C2(new_n772), .ZN(new_n852));
  INV_X1    g0652(.A(G303), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n805), .B1(new_n853), .B2(new_n775), .C1(new_n812), .C2(new_n220), .ZN(new_n854));
  INV_X1    g0654(.A(new_n798), .ZN(new_n855));
  INV_X1    g0655(.A(G311), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n602), .A2(new_n803), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n854), .B(new_n857), .C1(G283), .C2(new_n783), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n253), .B1(new_n791), .B2(new_n540), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n859), .B(KEYINPUT102), .Z(new_n860));
  INV_X1    g0660(.A(G294), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n858), .B(new_n860), .C1(new_n861), .C2(new_n807), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n852), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n815), .A2(new_n816), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n863), .A2(new_n815), .B1(new_n339), .B2(new_n864), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n762), .B(new_n865), .C1(new_n837), .C2(new_n817), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n844), .A2(new_n866), .ZN(G384));
  AOI21_X1  g0667(.A(new_n742), .B1(new_n728), .B2(KEYINPUT31), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n742), .A2(KEYINPUT31), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n837), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n396), .A2(new_n699), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n647), .B(new_n871), .C1(new_n651), .C2(new_n395), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n396), .B(new_n699), .C1(new_n427), .C2(new_n399), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n481), .B1(new_n638), .B2(new_n456), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n460), .A2(new_n466), .A3(new_n281), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n435), .ZN(new_n879));
  INV_X1    g0679(.A(new_n697), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n486), .B2(new_n493), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n490), .A2(new_n879), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n884), .A2(new_n484), .A3(new_n881), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT104), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n885), .A2(new_n886), .A3(KEYINPUT37), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n885), .A2(KEYINPUT37), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n487), .B1(new_n490), .B2(new_n880), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT37), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n889), .A2(new_n890), .A3(new_n484), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n888), .A2(KEYINPUT104), .A3(new_n891), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n883), .A2(KEYINPUT38), .A3(new_n887), .A4(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n891), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n890), .B1(new_n889), .B2(new_n484), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n635), .A2(new_n645), .A3(new_n485), .A4(new_n478), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n641), .A2(new_n697), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n893), .B1(new_n899), .B2(KEYINPUT38), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n876), .A2(KEYINPUT40), .A3(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT40), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n883), .A2(new_n887), .A3(new_n892), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT38), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n906), .A2(new_n893), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n874), .B(new_n837), .C1(new_n868), .C2(new_n869), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n903), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT105), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n906), .A2(new_n893), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n876), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n913), .A2(KEYINPUT105), .A3(new_n903), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n902), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n868), .A2(new_n869), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n495), .A2(new_n916), .ZN(new_n917));
  XOR2_X1   g0717(.A(new_n915), .B(new_n917), .Z(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(G330), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n652), .A2(new_n700), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT39), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n893), .B(new_n922), .C1(new_n899), .C2(KEYINPUT38), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n922), .B1(new_n906), .B2(new_n893), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n921), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n646), .A2(new_n880), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n838), .A2(new_n831), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(new_n912), .A3(new_n874), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n926), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n756), .B1(new_n725), .B2(new_n749), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n932), .A2(new_n495), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n659), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n931), .B(new_n934), .Z(new_n935));
  XNOR2_X1  g0735(.A(new_n919), .B(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n207), .B2(new_n759), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n220), .B1(new_n501), .B2(KEYINPUT35), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n938), .B(new_n227), .C1(KEYINPUT35), .C2(new_n501), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT36), .ZN(new_n940));
  OAI21_X1  g0740(.A(G77), .B1(new_n808), .B2(new_n386), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n941), .A2(new_n228), .B1(G50), .B2(new_n386), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n942), .A2(G1), .A3(new_n210), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n937), .A2(new_n940), .A3(new_n943), .ZN(G367));
  NAND2_X1  g0744(.A1(new_n614), .A2(new_n616), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n699), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n673), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n623), .B2(new_n946), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT43), .Z(new_n949));
  OAI21_X1  g0749(.A(new_n674), .B1(new_n506), .B2(new_n700), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n950), .B(new_n717), .C1(KEYINPUT42), .C2(new_n709), .ZN(new_n951));
  OAI21_X1  g0751(.A(KEYINPUT42), .B1(new_n716), .B2(new_n950), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n530), .B2(new_n699), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n949), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT106), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n957));
  OR3_X1    g0757(.A1(new_n951), .A2(new_n957), .A3(new_n953), .ZN(new_n958));
  OAI211_X1 g0758(.A(KEYINPUT106), .B(new_n949), .C1(new_n951), .C2(new_n953), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n956), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT107), .ZN(new_n961));
  INV_X1    g0761(.A(new_n714), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n950), .B1(new_n530), .B2(new_n700), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n960), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n961), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n960), .A2(new_n961), .A3(new_n964), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n719), .B(KEYINPUT41), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n710), .B(new_n715), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(new_n706), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n757), .A2(new_n972), .ZN(new_n973));
  AND3_X1   g0773(.A1(new_n712), .A2(KEYINPUT108), .A3(new_n713), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n717), .A2(new_n963), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n975), .A2(KEYINPUT44), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT44), .ZN(new_n977));
  NOR3_X1   g0777(.A1(new_n717), .A2(new_n977), .A3(new_n963), .ZN(new_n978));
  AND4_X1   g0778(.A1(KEYINPUT45), .A2(new_n716), .A3(new_n709), .A4(new_n963), .ZN(new_n979));
  AOI21_X1  g0779(.A(KEYINPUT45), .B1(new_n717), .B2(new_n963), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n976), .A2(new_n978), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n973), .B1(new_n974), .B2(new_n981), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n981), .A2(new_n974), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n970), .B1(new_n984), .B2(new_n757), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n967), .B(new_n968), .C1(new_n985), .C2(new_n761), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n783), .A2(G159), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n792), .A2(G58), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n798), .A2(G137), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n775), .A2(new_n846), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n772), .A2(new_n386), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n990), .B(new_n991), .C1(G150), .C2(new_n769), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n987), .A2(new_n988), .A3(new_n989), .A4(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n253), .B1(new_n797), .B2(G77), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT109), .Z(new_n995));
  AOI211_X1 g0795(.A(new_n993), .B(new_n995), .C1(G50), .C2(new_n786), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n803), .A2(new_n288), .ZN(new_n997));
  INV_X1    g0797(.A(G317), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n855), .A2(new_n998), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n772), .A2(new_n402), .B1(new_n775), .B2(new_n856), .ZN(new_n1000));
  INV_X1    g0800(.A(G283), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n253), .B1(new_n812), .B2(new_n1001), .ZN(new_n1002));
  NOR4_X1   g0802(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .A4(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n853), .B2(new_n807), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(G294), .B2(new_n783), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n792), .A2(G116), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT46), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n996), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT47), .Z(new_n1009));
  AOI21_X1  g0809(.A(new_n766), .B1(new_n1009), .B2(new_n815), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n821), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n819), .B1(new_n212), .B2(new_n416), .C1(new_n239), .C2(new_n1011), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1010), .B(new_n1012), .C1(new_n827), .C2(new_n948), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n986), .A2(new_n1013), .ZN(G387));
  OR2_X1    g0814(.A1(new_n757), .A2(new_n972), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1015), .A2(new_n719), .A3(new_n973), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n972), .A2(new_n761), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n786), .A2(G303), .B1(new_n776), .B2(G322), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n998), .B2(new_n807), .C1(new_n782), .C2(new_n856), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT48), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n1001), .B2(new_n772), .C1(new_n861), .C2(new_n791), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT49), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n798), .A2(G326), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n248), .B1(new_n797), .B2(G116), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n791), .A2(new_n339), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(KEYINPUT110), .B(G150), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1028), .B(new_n997), .C1(new_n798), .C2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(G159), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n416), .A2(new_n772), .B1(new_n1031), .B2(new_n775), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n248), .B1(new_n812), .B2(new_n386), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1032), .B(new_n1033), .C1(new_n783), .C2(new_n432), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1030), .B(new_n1034), .C1(new_n202), .C2(new_n807), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1027), .A2(new_n1035), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n236), .A2(new_n268), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1037), .A2(new_n821), .B1(new_n722), .B2(new_n823), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n317), .A2(G50), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT50), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n386), .B2(new_n339), .ZN(new_n1041));
  NOR3_X1   g0841(.A1(new_n1041), .A2(G45), .A3(new_n722), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n1038), .A2(new_n1042), .B1(G107), .B2(new_n212), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n1036), .A2(new_n815), .B1(new_n819), .B2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1044), .B(new_n762), .C1(new_n710), .C2(new_n827), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1016), .A2(new_n1017), .A3(new_n1045), .ZN(G393));
  OR2_X1    g0846(.A1(new_n981), .A2(new_n714), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n981), .A2(new_n714), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1047), .A2(new_n973), .A3(new_n1048), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n984), .A2(new_n1049), .A3(new_n719), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n761), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n769), .A2(G311), .B1(new_n776), .B2(G317), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT52), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n253), .B1(new_n812), .B2(new_n861), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n803), .A2(new_n540), .B1(new_n220), .B2(new_n772), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1055), .B(new_n1056), .C1(G322), .C2(new_n798), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n792), .A2(G283), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1054), .B(new_n1059), .C1(G303), .C2(new_n783), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n792), .A2(G68), .B1(new_n798), .B2(G143), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT112), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n769), .A2(G159), .B1(new_n776), .B2(G150), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT51), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n248), .B1(new_n339), .B2(new_n772), .C1(new_n812), .C2(new_n317), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n782), .A2(new_n202), .B1(new_n803), .B2(new_n602), .ZN(new_n1066));
  NOR4_X1   g0866(.A1(new_n1062), .A2(new_n1064), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n815), .B1(new_n1060), .B2(new_n1067), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n819), .B1(new_n288), .B2(new_n212), .C1(new_n246), .C2(new_n1011), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n762), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT111), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1068), .B(new_n1071), .C1(new_n963), .C2(new_n827), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1050), .A2(new_n1052), .A3(new_n1072), .ZN(G390));
  NAND2_X1  g0873(.A1(new_n900), .A2(new_n920), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n755), .A2(new_n700), .A3(new_n834), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n1075), .A2(new_n831), .B1(new_n872), .B2(new_n873), .ZN(new_n1076));
  OAI21_X1  g0876(.A(KEYINPUT113), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1075), .A2(new_n831), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n874), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT113), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1079), .A2(new_n1080), .A3(new_n920), .A4(new_n900), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1077), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n925), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n875), .B1(new_n838), .B2(new_n831), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1083), .B(new_n923), .C1(new_n1084), .C2(new_n921), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n837), .B(G330), .C1(new_n868), .C2(new_n746), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1086), .A2(new_n875), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1082), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT114), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n908), .B2(new_n692), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n742), .A2(KEYINPUT31), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n835), .B1(new_n744), .B2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1093), .A2(KEYINPUT114), .A3(G330), .A4(new_n874), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1091), .A2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1088), .B1(new_n1089), .B2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n831), .B(new_n1075), .C1(new_n1086), .C2(new_n875), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n874), .B1(new_n1093), .B2(G330), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1086), .A2(new_n875), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1091), .A2(new_n1094), .A3(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1099), .B1(new_n929), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT115), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n917), .B2(G330), .ZN(new_n1104));
  NOR4_X1   g0904(.A1(new_n495), .A2(new_n916), .A3(KEYINPUT115), .A4(new_n692), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n933), .B(new_n659), .C1(new_n1104), .C2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1102), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1096), .A2(new_n1107), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n1082), .A2(new_n1087), .A3(new_n1085), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1095), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1101), .A2(new_n929), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1099), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1106), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1111), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1108), .A2(new_n1117), .A3(new_n719), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1083), .A2(new_n816), .A3(new_n923), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n773), .A2(G77), .B1(new_n776), .B2(G283), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1120), .B(new_n253), .C1(new_n288), .C2(new_n812), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n783), .B2(new_n503), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n792), .A2(G87), .B1(new_n798), .B2(G294), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n769), .A2(G116), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1122), .A2(new_n849), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(G125), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n248), .B1(new_n855), .B2(new_n1126), .C1(new_n202), .C2(new_n803), .ZN(new_n1127));
  XOR2_X1   g0927(.A(new_n1127), .B(KEYINPUT116), .Z(new_n1128));
  AOI22_X1  g0928(.A1(new_n769), .A2(G132), .B1(new_n776), .B2(G128), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT117), .ZN(new_n1130));
  XOR2_X1   g0930(.A(KEYINPUT54), .B(G143), .Z(new_n1131));
  NAND2_X1  g0931(.A1(new_n786), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n792), .A2(new_n1029), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1132), .B1(new_n1133), .B2(KEYINPUT53), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1133), .A2(KEYINPUT53), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1134), .B(new_n1135), .C1(G137), .C2(new_n783), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1128), .A2(new_n1130), .A3(new_n1136), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n772), .A2(new_n1031), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1125), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1139), .A2(new_n815), .B1(new_n317), .B2(new_n864), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1119), .A2(new_n762), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(KEYINPUT118), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1141), .A2(KEYINPUT118), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n1096), .B2(new_n761), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1118), .A2(new_n1142), .A3(new_n1144), .ZN(G378));
  INV_X1    g0945(.A(KEYINPUT57), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n325), .A2(new_n880), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n360), .A2(new_n365), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1147), .B1(new_n658), .B2(new_n364), .ZN(new_n1150));
  OAI21_X1  g0950(.A(KEYINPUT55), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1148), .B1(new_n360), .B2(new_n365), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n658), .A2(new_n364), .A3(new_n1147), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT55), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1151), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT56), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1151), .A2(KEYINPUT56), .A3(new_n1155), .ZN(new_n1159));
  AND2_X1   g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n931), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1162), .A2(new_n926), .A3(new_n928), .A4(new_n930), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n909), .A2(new_n910), .ZN(new_n1165));
  AOI21_X1  g0965(.A(KEYINPUT105), .B1(new_n913), .B2(new_n903), .ZN(new_n1166));
  OAI211_X1 g0966(.A(G330), .B(new_n901), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(G330), .A2(new_n915), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1106), .B1(new_n1096), .B2(new_n1107), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1146), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1115), .B1(new_n1111), .B2(new_n1116), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n915), .A2(new_n1161), .A3(G330), .A4(new_n1163), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1173), .A2(new_n1176), .A3(KEYINPUT57), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1172), .A2(new_n719), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1160), .A2(new_n816), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n864), .A2(new_n202), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n803), .A2(new_n808), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1028), .B(new_n1181), .C1(G283), .C2(new_n798), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n248), .B1(new_n769), .B2(G107), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1183), .B(new_n258), .C1(new_n416), .C2(new_n812), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n991), .B(new_n1184), .C1(new_n783), .C2(G97), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1182), .B(new_n1185), .C1(new_n220), .C2(new_n775), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT58), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n783), .A2(G132), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n786), .A2(G137), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n792), .A2(new_n1131), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n769), .A2(G128), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n1126), .B2(new_n775), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G150), .B2(new_n773), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .A4(new_n1193), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n1194), .B(KEYINPUT59), .Z(new_n1195));
  AOI21_X1  g0995(.A(G41), .B1(new_n797), .B2(G159), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(KEYINPUT119), .A2(G124), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n855), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(KEYINPUT119), .A2(G124), .ZN(new_n1199));
  AOI21_X1  g0999(.A(G33), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1195), .A2(new_n1196), .A3(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n202), .B1(new_n251), .B2(G41), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1187), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n766), .B1(new_n1203), .B2(new_n815), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1179), .A2(new_n1180), .A3(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n1176), .B2(new_n761), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1178), .A2(new_n1207), .ZN(G375));
  AOI21_X1  g1008(.A(new_n253), .B1(new_n769), .B2(G137), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n773), .A2(G50), .B1(new_n776), .B2(G132), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1211), .B(new_n1181), .C1(new_n783), .C2(new_n1131), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n792), .A2(G159), .B1(new_n798), .B2(G128), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT121), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1212), .B(new_n1214), .C1(new_n322), .C2(new_n812), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n807), .A2(new_n1001), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n416), .A2(new_n772), .B1(new_n861), .B2(new_n775), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n253), .B1(new_n812), .B2(new_n402), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1217), .B(new_n1218), .C1(new_n783), .C2(G116), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n792), .A2(G97), .B1(new_n797), .B2(G77), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1219), .B(new_n1220), .C1(new_n853), .C2(new_n855), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1215), .B1(new_n1216), .B2(new_n1221), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1222), .A2(new_n815), .B1(new_n386), .B2(new_n864), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n762), .B(new_n1223), .C1(new_n874), .C2(new_n817), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n760), .B(KEYINPUT120), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1224), .B1(new_n1102), .B2(new_n1226), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1227), .B(KEYINPUT122), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1102), .A2(new_n1106), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1116), .A2(new_n1229), .A3(new_n969), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1228), .A2(new_n1230), .ZN(G381));
  AND3_X1   g1031(.A1(new_n1118), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1232));
  AND3_X1   g1032(.A1(new_n1178), .A2(new_n1232), .A3(new_n1207), .ZN(new_n1233));
  NOR3_X1   g1033(.A1(G381), .A2(G396), .A3(G393), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(G387), .A2(G384), .A3(G390), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .ZN(G407));
  NAND3_X1  g1036(.A1(new_n1178), .A2(new_n1232), .A3(new_n1207), .ZN(new_n1237));
  OAI211_X1 g1037(.A(G407), .B(G213), .C1(G343), .C2(new_n1237), .ZN(G409));
  INV_X1    g1038(.A(KEYINPUT124), .ZN(new_n1239));
  XOR2_X1   g1039(.A(G393), .B(G396), .Z(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n986), .A2(new_n1013), .A3(G390), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(G390), .B1(new_n986), .B2(new_n1013), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1241), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(G390), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(G387), .A2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1247), .A2(new_n1240), .A3(new_n1242), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1245), .A2(KEYINPUT123), .A3(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(KEYINPUT123), .B1(new_n1245), .B2(new_n1248), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT62), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1232), .B1(new_n1178), .B2(new_n1207), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n698), .A2(G213), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1225), .B1(new_n1173), .B2(new_n969), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1205), .B1(new_n1255), .B2(new_n1170), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1254), .B1(new_n1256), .B2(G378), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1253), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT60), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n720), .B1(new_n1229), .B2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1102), .A2(KEYINPUT60), .A3(new_n1106), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1260), .A2(new_n1116), .A3(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1228), .A2(G384), .A3(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(G384), .B1(new_n1228), .B2(new_n1262), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1252), .B1(new_n1258), .B2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1228), .A2(new_n1262), .ZN(new_n1268));
  INV_X1    g1068(.A(G384), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1263), .ZN(new_n1271));
  NOR4_X1   g1071(.A1(new_n1253), .A2(new_n1257), .A3(new_n1271), .A4(KEYINPUT62), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1267), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n698), .A2(G213), .A3(G2897), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1270), .A2(new_n1263), .A3(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1274), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1275), .B(new_n1277), .C1(new_n1253), .C2(new_n1257), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT61), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1251), .B1(new_n1273), .B2(new_n1280), .ZN(new_n1281));
  AOI22_X1  g1081(.A1(new_n1278), .A2(KEYINPUT63), .B1(new_n1258), .B2(new_n1266), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1173), .A2(new_n1176), .A3(KEYINPUT57), .ZN(new_n1283));
  AOI21_X1  g1083(.A(KEYINPUT57), .B1(new_n1173), .B2(new_n1176), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1283), .A2(new_n1284), .A3(new_n720), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1207), .ZN(new_n1286));
  OAI21_X1  g1086(.A(G378), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1226), .B1(new_n1171), .B2(new_n970), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1206), .B1(new_n1288), .B2(new_n1176), .ZN(new_n1289));
  AOI22_X1  g1089(.A1(new_n1289), .A2(new_n1232), .B1(G213), .B2(new_n698), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1287), .A2(KEYINPUT63), .A3(new_n1290), .A4(new_n1266), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1291), .A2(new_n1248), .A3(new_n1245), .ZN(new_n1292));
  NOR3_X1   g1092(.A1(new_n1282), .A2(new_n1292), .A3(KEYINPUT61), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1239), .B1(new_n1281), .B2(new_n1293), .ZN(new_n1294));
  OR3_X1    g1094(.A1(new_n1282), .A2(new_n1292), .A3(KEYINPUT61), .ZN(new_n1295));
  OR2_X1    g1095(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1287), .A2(new_n1290), .A3(new_n1266), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(KEYINPUT62), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1258), .A2(new_n1252), .A3(new_n1266), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1298), .A2(new_n1299), .A3(new_n1279), .A4(new_n1278), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1296), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1295), .A2(new_n1301), .A3(KEYINPUT124), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1294), .A2(new_n1302), .ZN(G405));
  OAI21_X1  g1103(.A(new_n1271), .B1(new_n1233), .B2(new_n1253), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(KEYINPUT126), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT126), .ZN(new_n1306));
  OAI211_X1 g1106(.A(new_n1306), .B(new_n1271), .C1(new_n1233), .C2(new_n1253), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1305), .A2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1287), .A2(new_n1237), .A3(new_n1266), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT125), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1287), .A2(KEYINPUT125), .A3(new_n1237), .A4(new_n1266), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT127), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1308), .A2(new_n1313), .A3(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1314), .B1(new_n1308), .B2(new_n1313), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1296), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1308), .A2(new_n1313), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(KEYINPUT127), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1308), .A2(new_n1313), .A3(new_n1314), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1319), .A2(new_n1251), .A3(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1317), .A2(new_n1321), .ZN(G402));
endmodule


