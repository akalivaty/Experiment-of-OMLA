//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 0 1 0 1 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n543,
    new_n544, new_n546, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n564, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n461), .A2(G137), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n469), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n462), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n465), .A2(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n467), .A2(new_n469), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G136), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n474), .A2(new_n462), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n476), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  NAND4_X1  g057(.A1(new_n467), .A2(new_n469), .A3(G126), .A4(G2105), .ZN(new_n483));
  OR2_X1    g058(.A1(G102), .A2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G114), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n484), .A2(new_n486), .A3(G2104), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT67), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n483), .A2(KEYINPUT67), .A3(new_n487), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n467), .A2(new_n469), .A3(G138), .A4(new_n462), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT68), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n461), .A2(G138), .A3(new_n462), .A4(new_n494), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n490), .A2(new_n491), .B1(new_n496), .B2(new_n497), .ZN(G164));
  XNOR2_X1  g073(.A(KEYINPUT5), .B(G543), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n499), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT6), .B(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G50), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  OAI22_X1  g084(.A1(new_n506), .A2(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n504), .A2(new_n505), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n502), .A2(new_n512), .ZN(G166));
  NAND3_X1  g088(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n514));
  XNOR2_X1  g089(.A(new_n514), .B(KEYINPUT7), .ZN(new_n515));
  INV_X1    g090(.A(G89), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n516), .B2(new_n510), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT69), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n517), .B(new_n518), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n503), .A2(G543), .ZN(new_n520));
  AND2_X1   g095(.A1(G63), .A2(G651), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n520), .A2(G51), .B1(new_n499), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(G168));
  NAND2_X1  g099(.A1(G77), .A2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n507), .A2(new_n506), .ZN(new_n526));
  INV_X1    g101(.A(G64), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT70), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n501), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n530), .B1(new_n529), .B2(new_n528), .ZN(new_n531));
  INV_X1    g106(.A(new_n510), .ZN(new_n532));
  AOI22_X1  g107(.A1(G52), .A2(new_n520), .B1(new_n532), .B2(G90), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(G301));
  INV_X1    g109(.A(G301), .ZN(G171));
  AOI22_X1  g110(.A1(new_n499), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n501), .ZN(new_n537));
  INV_X1    g112(.A(G43), .ZN(new_n538));
  INV_X1    g113(.A(G81), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n504), .A2(new_n538), .B1(new_n510), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  AND3_X1   g117(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G36), .ZN(new_n544));
  XOR2_X1   g119(.A(new_n544), .B(KEYINPUT71), .Z(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT72), .ZN(G188));
  INV_X1    g124(.A(KEYINPUT73), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n510), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n499), .A2(new_n503), .A3(KEYINPUT73), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n551), .A2(G91), .A3(new_n552), .ZN(new_n553));
  OAI211_X1 g128(.A(G53), .B(G543), .C1(new_n508), .C2(new_n509), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(KEYINPUT9), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT9), .ZN(new_n556));
  NAND4_X1  g131(.A1(new_n503), .A2(new_n556), .A3(G53), .A4(G543), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n526), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G651), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n553), .A2(new_n558), .A3(new_n562), .ZN(G299));
  INV_X1    g138(.A(KEYINPUT74), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n523), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n519), .A2(KEYINPUT74), .A3(new_n522), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(G286));
  OR2_X1    g143(.A1(new_n502), .A2(new_n512), .ZN(G303));
  INV_X1    g144(.A(G74), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n501), .B1(new_n526), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n571), .B1(G49), .B2(new_n520), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n551), .A2(G87), .A3(new_n552), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(G288));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n526), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n577), .A2(G651), .B1(new_n520), .B2(G48), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n551), .A2(G86), .A3(new_n552), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(G305));
  AOI22_X1  g155(.A1(new_n499), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n501), .ZN(new_n582));
  INV_X1    g157(.A(G47), .ZN(new_n583));
  INV_X1    g158(.A(G85), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n504), .A2(new_n583), .B1(new_n510), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n551), .A2(G92), .A3(new_n552), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT10), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n551), .A2(KEYINPUT10), .A3(G92), .A4(new_n552), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n526), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G651), .B1(new_n520), .B2(G54), .ZN(new_n597));
  AND2_X1   g172(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n588), .B1(new_n598), .B2(G868), .ZN(G284));
  OAI21_X1  g174(.A(new_n588), .B1(new_n598), .B2(G868), .ZN(G321));
  NOR2_X1   g175(.A1(G299), .A2(G868), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n601), .B1(new_n567), .B2(G868), .ZN(G297));
  AOI21_X1  g177(.A(new_n601), .B1(new_n567), .B2(G868), .ZN(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n598), .B1(new_n604), .B2(G860), .ZN(G148));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(new_n537), .B2(new_n540), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n593), .A2(new_n597), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n607), .B1(new_n609), .B2(new_n606), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g186(.A(KEYINPUT75), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G2100), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n475), .A2(G2104), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT12), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT13), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n612), .A2(G2100), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n613), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n475), .A2(G135), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n477), .A2(G123), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT76), .ZN(new_n621));
  NOR3_X1   g196(.A1(new_n621), .A2(new_n462), .A3(G111), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n462), .B2(G111), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n623), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n619), .B(new_n620), .C1(new_n622), .C2(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(G2096), .Z(new_n626));
  OAI211_X1 g201(.A(new_n618), .B(new_n626), .C1(new_n616), .C2(new_n613), .ZN(G156));
  XOR2_X1   g202(.A(G2451), .B(G2454), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT16), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT77), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2427), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2443), .B(G2446), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n639), .A2(new_n641), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n631), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n646), .A2(new_n630), .A3(new_n642), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n645), .A2(new_n647), .A3(G14), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(G401));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2072), .B(G2078), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT79), .ZN(new_n655));
  INV_X1    g230(.A(new_n650), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n651), .B(KEYINPUT17), .Z(new_n657));
  OAI21_X1  g232(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(new_n656), .A3(new_n653), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n653), .A2(new_n650), .A3(new_n651), .ZN(new_n660));
  XOR2_X1   g235(.A(KEYINPUT78), .B(KEYINPUT18), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n658), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2096), .B(G2100), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(G227));
  XOR2_X1   g240(.A(G1971), .B(G1976), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  XOR2_X1   g242(.A(G1956), .B(G2474), .Z(new_n668));
  XOR2_X1   g243(.A(G1961), .B(G1966), .Z(new_n669));
  AND2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n668), .A2(new_n669), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  MUX2_X1   g250(.A(new_n675), .B(new_n674), .S(new_n667), .Z(new_n676));
  OR3_X1    g251(.A1(new_n673), .A2(new_n676), .A3(G1981), .ZN(new_n677));
  OAI21_X1  g252(.A(G1981), .B1(new_n673), .B2(new_n676), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT80), .B(KEYINPUT81), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  INV_X1    g259(.A(G1986), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n682), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n677), .A2(new_n678), .A3(new_n687), .ZN(new_n688));
  AND3_X1   g263(.A1(new_n683), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n686), .B1(new_n683), .B2(new_n688), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(G229));
  XNOR2_X1  g266(.A(KEYINPUT30), .B(G28), .ZN(new_n692));
  INV_X1    g267(.A(G29), .ZN(new_n693));
  OR2_X1    g268(.A1(KEYINPUT31), .A2(G11), .ZN(new_n694));
  NAND2_X1  g269(.A1(KEYINPUT31), .A2(G11), .ZN(new_n695));
  AOI22_X1  g270(.A1(new_n692), .A2(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(new_n625), .B2(new_n693), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT82), .B(G16), .Z(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n699), .A2(G19), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n541), .B2(new_n699), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(G1341), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT90), .B(G2067), .Z(new_n703));
  NAND2_X1  g278(.A1(new_n693), .A2(G26), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT28), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n475), .A2(G140), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n477), .A2(G128), .ZN(new_n707));
  OR2_X1    g282(.A1(G104), .A2(G2105), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n708), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n706), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n705), .B1(new_n711), .B2(new_n693), .ZN(new_n712));
  AOI211_X1 g287(.A(new_n697), .B(new_n702), .C1(new_n703), .C2(new_n712), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n712), .A2(new_n703), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT24), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n693), .B1(new_n715), .B2(G34), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n715), .B2(G34), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G160), .B2(G29), .ZN(new_n718));
  INV_X1    g293(.A(G2084), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(G16), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G21), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G168), .B2(new_n721), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(G5), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G171), .B2(new_n721), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n723), .A2(G1966), .B1(G1961), .B2(new_n725), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n713), .A2(new_n714), .A3(new_n720), .A4(new_n726), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n693), .A2(G33), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT91), .B(KEYINPUT25), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n729), .A2(new_n730), .ZN(new_n732));
  INV_X1    g307(.A(G139), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n461), .A2(new_n462), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n731), .B(new_n732), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT92), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(new_n462), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n728), .B1(new_n739), .B2(G29), .ZN(new_n740));
  INV_X1    g315(.A(G2072), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT96), .B(G1956), .Z(new_n742));
  NAND2_X1  g317(.A1(new_n698), .A2(G20), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT23), .Z(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G16), .B2(G299), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n740), .A2(new_n741), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n693), .A2(G32), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n477), .A2(G129), .ZN(new_n748));
  NAND3_X1  g323(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT26), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n752));
  INV_X1    g327(.A(G141), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n734), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n747), .B1(new_n755), .B2(new_n693), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT93), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT27), .B(G1996), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(G2090), .ZN(new_n760));
  NOR2_X1   g335(.A1(G29), .A2(G35), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G162), .B2(G29), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n746), .B(new_n759), .C1(new_n760), .C2(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n727), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n764), .A2(new_n760), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT95), .ZN(new_n768));
  NOR2_X1   g343(.A1(G4), .A2(G16), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT87), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n598), .B2(G16), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT89), .B(G1348), .Z(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT88), .Z(new_n773));
  XNOR2_X1  g348(.A(new_n771), .B(new_n773), .ZN(new_n774));
  OAI22_X1  g349(.A1(new_n757), .A2(new_n758), .B1(new_n740), .B2(new_n741), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n693), .A2(G27), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G164), .B2(new_n693), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(G2078), .Z(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n723), .B2(G1966), .ZN(new_n779));
  OAI22_X1  g354(.A1(new_n725), .A2(G1961), .B1(new_n742), .B2(new_n745), .ZN(new_n780));
  NOR3_X1   g355(.A1(new_n775), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n766), .A2(new_n768), .A3(new_n774), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n721), .A2(G23), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n572), .A2(new_n573), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(new_n721), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT33), .B(G1976), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT85), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n785), .B(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n699), .A2(G22), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G166), .B2(new_n699), .ZN(new_n790));
  INV_X1    g365(.A(G1971), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n721), .A2(G6), .ZN(new_n794));
  INV_X1    g369(.A(G305), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(new_n721), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT32), .B(G1981), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(KEYINPUT86), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT86), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n793), .A2(new_n801), .A3(new_n798), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT84), .B(KEYINPUT34), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n804), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n800), .A2(new_n802), .A3(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n699), .A2(G24), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n586), .B(KEYINPUT83), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(new_n699), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1986), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n693), .A2(G25), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n475), .A2(G131), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n477), .A2(G119), .ZN(new_n814));
  OR2_X1    g389(.A1(G95), .A2(G2105), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n815), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n816));
  AND3_X1   g391(.A1(new_n813), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n812), .B1(new_n817), .B2(new_n693), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT35), .B(G1991), .Z(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n818), .B(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n811), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n805), .A2(new_n807), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(KEYINPUT36), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT36), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n805), .A2(new_n825), .A3(new_n807), .A4(new_n822), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n782), .B1(new_n824), .B2(new_n826), .ZN(G311));
  INV_X1    g402(.A(KEYINPUT97), .ZN(new_n828));
  XNOR2_X1  g403(.A(G311), .B(new_n828), .ZN(G150));
  AOI22_X1  g404(.A1(new_n499), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n830), .A2(new_n501), .ZN(new_n831));
  INV_X1    g406(.A(G55), .ZN(new_n832));
  INV_X1    g407(.A(G93), .ZN(new_n833));
  OAI22_X1  g408(.A1(new_n504), .A2(new_n832), .B1(new_n510), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(G860), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT37), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n598), .A2(G559), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT38), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n541), .B(new_n835), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(KEYINPUT39), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT98), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n842), .A2(KEYINPUT39), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n845), .A2(G860), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n838), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT99), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(G145));
  XNOR2_X1  g424(.A(new_n481), .B(G160), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(new_n625), .Z(new_n851));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n475), .A2(G142), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n477), .A2(G130), .ZN(new_n854));
  OR2_X1    g429(.A1(G106), .A2(G2105), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n855), .B(G2104), .C1(G118), .C2(new_n462), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n615), .A2(new_n853), .A3(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT12), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n614), .B(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n857), .A2(new_n853), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n858), .A2(new_n862), .A3(new_n817), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n817), .B1(new_n858), .B2(new_n862), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n852), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n858), .A2(new_n862), .ZN(new_n867));
  INV_X1    g442(.A(new_n817), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n869), .A2(KEYINPUT100), .A3(new_n863), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n755), .B(new_n710), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n496), .A2(new_n497), .ZN(new_n873));
  INV_X1    g448(.A(new_n488), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n739), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n739), .A2(new_n876), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n872), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n879), .ZN(new_n881));
  INV_X1    g456(.A(new_n872), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n881), .A2(new_n882), .A3(new_n877), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n871), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT100), .B1(new_n869), .B2(new_n863), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n885), .B1(new_n880), .B2(new_n883), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n851), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n871), .A2(new_n880), .A3(new_n883), .ZN(new_n888));
  INV_X1    g463(.A(new_n851), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n880), .A2(new_n883), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n888), .B(new_n889), .C1(new_n890), .C2(new_n885), .ZN(new_n891));
  INV_X1    g466(.A(G37), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n887), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g469(.A1(new_n795), .A2(G288), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n784), .A2(G305), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n898));
  XNOR2_X1  g473(.A(G166), .B(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(G290), .ZN(new_n900));
  XNOR2_X1  g475(.A(G166), .B(KEYINPUT103), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n586), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n897), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n897), .A2(new_n902), .A3(new_n900), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n904), .A2(new_n905), .A3(KEYINPUT104), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT104), .ZN(new_n907));
  INV_X1    g482(.A(new_n905), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n907), .B1(new_n908), .B2(new_n903), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n910), .A2(KEYINPUT42), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT105), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n908), .A2(new_n903), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n912), .B1(new_n913), .B2(KEYINPUT42), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n911), .A2(KEYINPUT105), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT101), .ZN(new_n917));
  OR2_X1    g492(.A1(G299), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n598), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(G299), .A2(new_n917), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n598), .A2(new_n920), .A3(new_n918), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XOR2_X1   g499(.A(KEYINPUT102), .B(KEYINPUT41), .Z(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  XOR2_X1   g502(.A(new_n841), .B(new_n609), .Z(new_n928));
  INV_X1    g503(.A(KEYINPUT41), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n922), .A2(new_n929), .A3(new_n923), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n924), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n931), .B1(new_n928), .B2(new_n932), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n915), .A2(new_n916), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n933), .B1(new_n915), .B2(new_n916), .ZN(new_n935));
  OAI21_X1  g510(.A(G868), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n836), .A2(new_n606), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(G295));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n937), .ZN(G331));
  INV_X1    g514(.A(new_n841), .ZN(new_n940));
  AOI21_X1  g515(.A(G301), .B1(new_n565), .B2(new_n566), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n523), .A2(G301), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n940), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n566), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT74), .B1(new_n519), .B2(new_n522), .ZN(new_n946));
  OAI21_X1  g521(.A(G171), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n947), .A2(new_n841), .A3(new_n942), .ZN(new_n948));
  AOI22_X1  g523(.A1(new_n927), .A2(new_n930), .B1(new_n944), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n944), .A2(new_n948), .A3(KEYINPUT106), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT106), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n947), .A2(new_n951), .A3(new_n841), .A4(new_n942), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n949), .B1(new_n953), .B2(new_n932), .ZN(new_n954));
  AOI21_X1  g529(.A(G37), .B1(new_n954), .B2(new_n910), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n932), .A2(new_n944), .A3(new_n948), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n924), .A2(new_n929), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(new_n924), .B2(new_n925), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n956), .B1(new_n953), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n906), .A2(new_n909), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n955), .A2(KEYINPUT43), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n924), .B1(new_n950), .B2(new_n952), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n960), .B1(new_n963), .B2(new_n949), .ZN(new_n964));
  AOI21_X1  g539(.A(KEYINPUT43), .B1(new_n955), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT44), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n953), .A2(new_n932), .ZN(new_n967));
  INV_X1    g542(.A(new_n949), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(new_n910), .A3(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n969), .A2(new_n892), .A3(new_n964), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n955), .A2(new_n972), .A3(new_n961), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n966), .B1(new_n975), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g551(.A(G2067), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n710), .B(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(G1996), .B1(new_n751), .B2(new_n754), .ZN(new_n979));
  INV_X1    g554(.A(G1996), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n978), .A2(new_n979), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(G1384), .B1(new_n873), .B2(new_n874), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n983), .A2(KEYINPUT45), .ZN(new_n984));
  INV_X1    g559(.A(G40), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n465), .A2(new_n472), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n982), .A2(new_n988), .ZN(new_n989));
  XOR2_X1   g564(.A(new_n989), .B(KEYINPUT107), .Z(new_n990));
  NOR2_X1   g565(.A1(new_n817), .A2(new_n819), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n868), .A2(new_n820), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n988), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n987), .A2(G1986), .A3(G290), .ZN(new_n995));
  XOR2_X1   g570(.A(new_n995), .B(KEYINPUT48), .Z(new_n996));
  NAND2_X1  g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n988), .A2(KEYINPUT46), .A3(new_n980), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT46), .B1(new_n988), .B2(new_n980), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n987), .B1(new_n755), .B2(new_n978), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  XOR2_X1   g576(.A(new_n1001), .B(KEYINPUT47), .Z(new_n1002));
  NAND2_X1  g577(.A1(new_n990), .A2(new_n992), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n711), .A2(new_n977), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n987), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT126), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n997), .B(new_n1002), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1007), .B1(new_n1006), .B2(new_n1005), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(G164), .B2(G1384), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n470), .A2(new_n471), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(G2105), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1012), .A2(G40), .A3(new_n464), .A4(new_n463), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1013), .B1(new_n983), .B2(KEYINPUT45), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1010), .A2(new_n1014), .A3(new_n980), .ZN(new_n1015));
  XNOR2_X1  g590(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1016), .B(G1341), .ZN(new_n1017));
  INV_X1    g592(.A(G1384), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n875), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1017), .B1(new_n1019), .B2(new_n1013), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1015), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n541), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT59), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT50), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1013), .B1(new_n983), .B2(new_n1025), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n483), .A2(KEYINPUT67), .A3(new_n487), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT67), .B1(new_n483), .B2(new_n487), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n873), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1025), .B1(new_n1029), .B2(new_n1018), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1026), .B1(new_n1030), .B2(KEYINPUT109), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT109), .ZN(new_n1032));
  AOI211_X1 g607(.A(new_n1032), .B(new_n1025), .C1(new_n1029), .C2(new_n1018), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n772), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n593), .A2(KEYINPUT60), .A3(new_n597), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT121), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT121), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n593), .A2(new_n1037), .A3(KEYINPUT60), .A4(new_n597), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n983), .A2(new_n977), .A3(new_n986), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT60), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n608), .A2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1034), .A2(new_n1039), .A3(new_n1040), .A4(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1021), .A2(KEYINPUT59), .A3(new_n541), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1024), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT120), .ZN(new_n1046));
  INV_X1    g621(.A(G1956), .ZN(new_n1047));
  AND3_X1   g622(.A1(new_n1029), .A2(new_n1025), .A3(new_n1018), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n986), .B1(new_n983), .B2(new_n1025), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1047), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n1051));
  OR2_X1    g626(.A1(new_n1051), .A2(KEYINPUT57), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n553), .A2(new_n558), .A3(new_n562), .A4(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(KEYINPUT57), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n1053), .B(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g630(.A(KEYINPUT56), .B(G2072), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1010), .A2(new_n1014), .A3(new_n1056), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1050), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1055), .B1(new_n1050), .B2(new_n1057), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1046), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT61), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1034), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1062), .A2(new_n1038), .A3(new_n1036), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT61), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1046), .B(new_n1064), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1045), .A2(new_n1061), .A3(new_n1063), .A4(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1034), .A2(new_n1040), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1059), .B1(new_n1067), .B2(new_n598), .ZN(new_n1068));
  OR2_X1    g643(.A1(new_n1068), .A2(new_n1058), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n523), .A2(G8), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1029), .A2(KEYINPUT45), .A3(new_n1018), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1013), .B1(new_n1019), .B2(new_n1009), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1029), .A2(KEYINPUT116), .A3(KEYINPUT45), .A4(new_n1018), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G1966), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n1032), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1030), .A2(KEYINPUT109), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1081), .A2(new_n1082), .A3(new_n719), .A4(new_n1026), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1071), .B1(new_n1079), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT51), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT122), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1086), .B1(new_n1071), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1079), .A2(new_n1083), .ZN(new_n1089));
  OAI211_X1 g664(.A(G8), .B(new_n1088), .C1(new_n1089), .C2(new_n523), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1071), .ZN(new_n1092));
  AOI211_X1 g667(.A(new_n1092), .B(new_n1088), .C1(new_n1089), .C2(G8), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1085), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(G1961), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT53), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1097), .B1(new_n1098), .B2(G2078), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1097), .A2(G2078), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1075), .B(new_n1100), .C1(new_n1009), .C2(new_n1019), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1096), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .A4(new_n1100), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1096), .A2(new_n1099), .A3(G301), .A4(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1107));
  OAI221_X1 g682(.A(KEYINPUT54), .B1(G301), .B2(new_n1102), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(G1976), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT52), .B1(G288), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G8), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1111), .B1(new_n983), .B2(new_n986), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n572), .A2(new_n573), .A3(G1976), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1110), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT112), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT112), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1110), .A2(new_n1112), .A3(new_n1116), .A4(new_n1113), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT111), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1112), .A2(KEYINPUT111), .A3(new_n1113), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1121), .A2(KEYINPUT52), .A3(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT113), .B(G1981), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n578), .A2(new_n579), .A3(new_n1124), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n499), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1126));
  INV_X1    g701(.A(G48), .ZN(new_n1127));
  OAI22_X1  g702(.A1(new_n1126), .A2(new_n501), .B1(new_n1127), .B2(new_n504), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n532), .A2(G86), .ZN(new_n1129));
  OAI21_X1  g704(.A(G1981), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1125), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT49), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1125), .A2(new_n1130), .A3(KEYINPUT49), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1133), .A2(new_n1112), .A3(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1118), .A2(new_n1123), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  XOR2_X1   g712(.A(KEYINPUT110), .B(G2090), .Z(new_n1138));
  NAND4_X1  g713(.A1(new_n1081), .A2(new_n1082), .A3(new_n1026), .A4(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1098), .A2(new_n791), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1111), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1142));
  OAI211_X1 g717(.A(KEYINPUT55), .B(G8), .C1(new_n502), .C2(new_n512), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1141), .A2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1148), .A2(new_n1138), .B1(new_n1098), .B2(new_n791), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1145), .B1(new_n1149), .B2(new_n1111), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1137), .A2(new_n1147), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1096), .A2(new_n1099), .A3(new_n1103), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(G171), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1096), .A2(new_n1099), .A3(G301), .A4(new_n1101), .ZN(new_n1154));
  AOI21_X1  g729(.A(KEYINPUT54), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1151), .A2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1070), .A2(new_n1094), .A3(new_n1108), .A4(new_n1156), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1137), .B(KEYINPUT117), .C1(new_n1146), .C2(new_n1141), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1089), .A2(G8), .A3(new_n567), .ZN(new_n1159));
  AOI211_X1 g734(.A(new_n1111), .B(new_n1145), .C1(new_n1139), .C2(new_n1140), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT63), .ZN(new_n1161));
  NOR3_X1   g736(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT117), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1141), .A2(new_n1146), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1163), .B1(new_n1164), .B2(new_n1136), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1158), .A2(new_n1162), .A3(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1161), .B1(new_n1151), .B2(new_n1159), .ZN(new_n1167));
  XOR2_X1   g742(.A(new_n1112), .B(KEYINPUT114), .Z(new_n1168));
  NOR2_X1   g743(.A1(G288), .A2(G1976), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1135), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1125), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1168), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1172), .B1(new_n1147), .B2(new_n1136), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT115), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  OAI211_X1 g750(.A(new_n1172), .B(KEYINPUT115), .C1(new_n1147), .C2(new_n1136), .ZN(new_n1176));
  AOI22_X1  g751(.A1(new_n1166), .A2(new_n1167), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  AND3_X1   g752(.A1(new_n1157), .A2(new_n1177), .A3(KEYINPUT124), .ZN(new_n1178));
  AOI21_X1  g753(.A(KEYINPUT124), .B1(new_n1157), .B2(new_n1177), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1088), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1181));
  AOI22_X1  g756(.A1(new_n1181), .A2(new_n719), .B1(new_n1078), .B2(new_n1077), .ZN(new_n1182));
  OAI211_X1 g757(.A(new_n1071), .B(new_n1180), .C1(new_n1182), .C2(new_n1111), .ZN(new_n1183));
  AOI211_X1 g758(.A(KEYINPUT62), .B(new_n1084), .C1(new_n1183), .C2(new_n1090), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1153), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1185), .A2(new_n1147), .A3(new_n1150), .A4(new_n1137), .ZN(new_n1186));
  OAI21_X1  g761(.A(KEYINPUT125), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT62), .ZN(new_n1188));
  OAI211_X1 g763(.A(new_n1188), .B(new_n1085), .C1(new_n1091), .C2(new_n1093), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1186), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT125), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1094), .A2(KEYINPUT62), .ZN(new_n1193));
  AND3_X1   g768(.A1(new_n1187), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  NOR3_X1   g769(.A1(new_n1178), .A2(new_n1179), .A3(new_n1194), .ZN(new_n1195));
  XNOR2_X1  g770(.A(new_n586), .B(G1986), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n994), .B1(new_n987), .B2(new_n1196), .ZN(new_n1197));
  XOR2_X1   g772(.A(new_n1197), .B(KEYINPUT108), .Z(new_n1198));
  OAI21_X1  g773(.A(new_n1008), .B1(new_n1195), .B2(new_n1198), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g774(.A(G229), .ZN(new_n1201));
  NOR2_X1   g775(.A1(G227), .A2(new_n459), .ZN(new_n1202));
  AND2_X1   g776(.A1(new_n648), .A2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g777(.A1(new_n893), .A2(new_n1201), .A3(new_n1203), .ZN(new_n1204));
  AOI211_X1 g778(.A(KEYINPUT127), .B(new_n1204), .C1(new_n971), .C2(new_n973), .ZN(new_n1205));
  INV_X1    g779(.A(KEYINPUT127), .ZN(new_n1206));
  INV_X1    g780(.A(new_n1204), .ZN(new_n1207));
  AOI21_X1  g781(.A(new_n1206), .B1(new_n974), .B2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g782(.A1(new_n1205), .A2(new_n1208), .ZN(G308));
  AND3_X1   g783(.A1(new_n955), .A2(new_n972), .A3(new_n961), .ZN(new_n1210));
  AOI21_X1  g784(.A(new_n972), .B1(new_n955), .B2(new_n964), .ZN(new_n1211));
  OAI21_X1  g785(.A(new_n1207), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g786(.A1(new_n1212), .A2(KEYINPUT127), .ZN(new_n1213));
  NAND3_X1  g787(.A1(new_n974), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1214));
  NAND2_X1  g788(.A1(new_n1213), .A2(new_n1214), .ZN(G225));
endmodule


