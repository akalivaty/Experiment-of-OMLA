//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 0 0 0 1 0 0 0 0 1 0 1 1 1 1 0 0 0 1 0 1 1 1 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n569, new_n570, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT64), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n454), .A2(new_n458), .B1(new_n459), .B2(new_n455), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  XNOR2_X1  g040(.A(new_n465), .B(KEYINPUT68), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n462), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT69), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n469), .A2(new_n471), .A3(KEYINPUT3), .ZN(new_n472));
  OR2_X1    g047(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n472), .A2(G137), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n469), .A2(new_n471), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n467), .B1(new_n477), .B2(new_n462), .ZN(G160));
  AND3_X1   g053(.A1(new_n472), .A2(KEYINPUT70), .A3(new_n473), .ZN(new_n479));
  AOI21_X1  g054(.A(KEYINPUT70), .B1(new_n472), .B2(new_n473), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n462), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n462), .A2(G112), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  OAI22_X1  g059(.A1(new_n481), .A2(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g060(.A(G2105), .B1(new_n479), .B2(new_n480), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT71), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g063(.A(KEYINPUT71), .B(G2105), .C1(new_n479), .C2(new_n480), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n485), .B1(new_n490), .B2(G124), .ZN(G162));
  AND2_X1   g066(.A1(G126), .A2(G2105), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n472), .A2(new_n473), .A3(new_n492), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G114), .C2(new_n462), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n462), .A2(G138), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n472), .A2(new_n473), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT72), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n498), .A2(new_n501), .A3(KEYINPUT4), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n463), .A2(new_n504), .A3(new_n497), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n496), .B1(new_n503), .B2(new_n505), .ZN(G164));
  XNOR2_X1  g081(.A(KEYINPUT5), .B(G543), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n507), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n510), .A2(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  AND2_X1   g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT73), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT73), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n507), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g098(.A1(G63), .A2(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n521), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT6), .B(G651), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT74), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n512), .A2(KEYINPUT74), .A3(new_n513), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n528), .A2(G543), .A3(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G51), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n525), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT75), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g109(.A(new_n525), .B(KEYINPUT75), .C1(new_n530), .C2(new_n531), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n507), .A2(new_n526), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT76), .B(KEYINPUT7), .ZN(new_n538));
  AND3_X1   g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n538), .A2(new_n539), .ZN(new_n541));
  AOI22_X1  g116(.A1(G89), .A2(new_n537), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n534), .A2(new_n535), .A3(new_n542), .ZN(G286));
  INV_X1    g118(.A(G286), .ZN(G168));
  NAND3_X1  g119(.A1(new_n521), .A2(new_n523), .A3(G64), .ZN(new_n545));
  NAND2_X1  g120(.A1(G77), .A2(G543), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT77), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n545), .A2(KEYINPUT77), .A3(new_n546), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n549), .A2(G651), .A3(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n530), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n552), .A2(G52), .B1(G90), .B2(new_n537), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n551), .A2(new_n553), .ZN(G301));
  INV_X1    g129(.A(G301), .ZN(G171));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n521), .A2(new_n523), .ZN(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G651), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n537), .A2(G81), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n528), .A2(G43), .A3(G543), .A4(new_n529), .ZN(new_n562));
  AND3_X1   g137(.A1(new_n561), .A2(KEYINPUT78), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g138(.A(KEYINPUT78), .B1(new_n561), .B2(new_n562), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n560), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(G188));
  NAND4_X1  g146(.A1(new_n528), .A2(G53), .A3(G543), .A4(new_n529), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT9), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G65), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n520), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n537), .A2(G91), .B1(new_n576), .B2(G651), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n573), .A2(new_n577), .ZN(G299));
  NAND2_X1  g153(.A1(new_n537), .A2(G87), .ZN(new_n579));
  INV_X1    g154(.A(G49), .ZN(new_n580));
  AOI21_X1  g155(.A(G74), .B1(new_n521), .B2(new_n523), .ZN(new_n581));
  OAI221_X1 g156(.A(new_n579), .B1(new_n530), .B2(new_n580), .C1(new_n581), .C2(new_n509), .ZN(G288));
  NAND2_X1  g157(.A1(G48), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G86), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n520), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(new_n526), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(new_n587));
  OAI21_X1  g162(.A(G61), .B1(new_n518), .B2(new_n519), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n509), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT79), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI211_X1 g167(.A(KEYINPUT79), .B(new_n509), .C1(new_n588), .C2(new_n589), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n587), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G305));
  INV_X1    g171(.A(G47), .ZN(new_n597));
  INV_X1    g172(.A(G85), .ZN(new_n598));
  OAI22_X1  g173(.A1(new_n530), .A2(new_n597), .B1(new_n598), .B2(new_n536), .ZN(new_n599));
  INV_X1    g174(.A(G60), .ZN(new_n600));
  INV_X1    g175(.A(G72), .ZN(new_n601));
  INV_X1    g176(.A(G543), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n557), .A2(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(KEYINPUT80), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT80), .ZN(new_n605));
  OAI221_X1 g180(.A(new_n605), .B1(new_n601), .B2(new_n602), .C1(new_n557), .C2(new_n600), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n604), .A2(G651), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n599), .B1(new_n607), .B2(KEYINPUT81), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT81), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n604), .A2(new_n609), .A3(new_n606), .A4(G651), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n608), .A2(new_n610), .ZN(G290));
  NAND3_X1  g186(.A1(new_n537), .A2(KEYINPUT10), .A3(G92), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT10), .ZN(new_n613));
  INV_X1    g188(.A(G92), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n536), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(G79), .A2(G543), .ZN(new_n616));
  INV_X1    g191(.A(G66), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n520), .B2(new_n617), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n612), .A2(new_n615), .B1(G651), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n552), .A2(G54), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(G868), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G171), .B2(new_n622), .ZN(G284));
  OAI21_X1  g199(.A(new_n623), .B1(G171), .B2(new_n622), .ZN(G321));
  NAND2_X1  g200(.A1(G299), .A2(new_n622), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G168), .B2(new_n622), .ZN(G280));
  XOR2_X1   g202(.A(G280), .B(KEYINPUT82), .Z(G297));
  INV_X1    g203(.A(new_n621), .ZN(new_n629));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(G860), .ZN(G148));
  OR3_X1    g206(.A1(new_n621), .A2(KEYINPUT83), .A3(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(KEYINPUT83), .B1(new_n621), .B2(G559), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  MUX2_X1   g209(.A(new_n565), .B(new_n634), .S(G868), .Z(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g211(.A(G135), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n462), .A2(G111), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n639));
  OAI22_X1  g214(.A1(new_n481), .A2(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n640), .B1(new_n490), .B2(G123), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n641), .A2(KEYINPUT86), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(KEYINPUT86), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n644), .A2(G2096), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(G2096), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n475), .A2(new_n463), .A3(new_n462), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT12), .Z(new_n648));
  XOR2_X1   g223(.A(KEYINPUT84), .B(KEYINPUT13), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT85), .B(G2100), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n645), .A2(new_n646), .A3(new_n652), .ZN(G156));
  INV_X1    g228(.A(KEYINPUT14), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2427), .B(G2438), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2430), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT15), .B(G2435), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n654), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n658), .B1(new_n657), .B2(new_n656), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2451), .B(G2454), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1341), .B(G1348), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n659), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2443), .B(G2446), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  AND3_X1   g242(.A1(new_n666), .A2(G14), .A3(new_n667), .ZN(G401));
  XOR2_X1   g243(.A(G2072), .B(G2078), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT17), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n672), .B2(new_n669), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n673), .B1(KEYINPUT87), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n676), .B1(KEYINPUT87), .B2(new_n675), .ZN(new_n677));
  INV_X1    g252(.A(new_n669), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n678), .A2(new_n674), .A3(new_n671), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT18), .Z(new_n680));
  NAND3_X1  g255(.A1(new_n670), .A2(new_n674), .A3(new_n672), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n677), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G2096), .B(G2100), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(G227));
  XOR2_X1   g259(.A(G1971), .B(G1976), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT19), .ZN(new_n686));
  XOR2_X1   g261(.A(G1956), .B(G2474), .Z(new_n687));
  XOR2_X1   g262(.A(G1961), .B(G1966), .Z(new_n688));
  AND2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT20), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n687), .A2(new_n688), .ZN(new_n692));
  NOR3_X1   g267(.A1(new_n686), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(new_n686), .B2(new_n692), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT88), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n695), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1991), .B(G1996), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(G229));
  NAND3_X1  g279(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT26), .Z(new_n706));
  NAND3_X1  g281(.A1(new_n475), .A2(G105), .A3(new_n462), .ZN(new_n707));
  INV_X1    g282(.A(G141), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n706), .B(new_n707), .C1(new_n481), .C2(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n490), .B2(G129), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT96), .Z(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G29), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G29), .B2(G32), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT27), .B(G1996), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT97), .Z(new_n716));
  NOR2_X1   g291(.A1(G4), .A2(G16), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n629), .B2(G16), .ZN(new_n718));
  INV_X1    g293(.A(G1348), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(G29), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT24), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(G34), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n722), .B2(G34), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G160), .B2(G29), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n720), .B1(G2084), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n721), .A2(G27), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G164), .B2(new_n721), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n726), .B1(G2078), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n721), .A2(G26), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT28), .ZN(new_n731));
  INV_X1    g306(.A(G140), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n462), .A2(G116), .ZN(new_n733));
  OAI21_X1  g308(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n734));
  OAI22_X1  g309(.A1(new_n481), .A2(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(new_n490), .B2(G128), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n731), .B1(new_n736), .B2(new_n721), .ZN(new_n737));
  INV_X1    g312(.A(G2067), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n566), .A2(G16), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G16), .B2(G19), .ZN(new_n741));
  INV_X1    g316(.A(G1341), .ZN(new_n742));
  INV_X1    g317(.A(G16), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G21), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G168), .B2(new_n743), .ZN(new_n745));
  OAI22_X1  g320(.A1(new_n741), .A2(new_n742), .B1(G1966), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G1966), .B2(new_n745), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n728), .A2(G2078), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n741), .B2(new_n742), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n729), .A2(new_n739), .A3(new_n747), .A4(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n713), .A2(new_n714), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n743), .A2(G5), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G171), .B2(new_n743), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G1961), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n721), .A2(G33), .ZN(new_n755));
  INV_X1    g330(.A(new_n481), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G139), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n463), .A2(G127), .ZN(new_n758));
  INV_X1    g333(.A(G115), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n759), .B2(new_n468), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT25), .ZN(new_n761));
  NAND2_X1  g336(.A1(G103), .A2(G2104), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(new_n762), .B2(G2105), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n462), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n760), .A2(G2105), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n757), .A2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n755), .B1(new_n767), .B2(new_n721), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n768), .A2(G2072), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(G2072), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT30), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n771), .A2(G28), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n721), .B1(new_n771), .B2(G28), .ZN(new_n773));
  AND2_X1   g348(.A1(KEYINPUT31), .A2(G11), .ZN(new_n774));
  NOR2_X1   g349(.A1(KEYINPUT31), .A2(G11), .ZN(new_n775));
  OAI22_X1  g350(.A1(new_n772), .A2(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n725), .B2(G2084), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n770), .A2(new_n777), .ZN(new_n778));
  NOR3_X1   g353(.A1(new_n754), .A2(new_n769), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n721), .A2(G35), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G162), .B2(new_n721), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT29), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n782), .A2(G2090), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n642), .A2(G29), .A3(new_n643), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n779), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n750), .A2(new_n751), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n782), .A2(G2090), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT98), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n743), .A2(G20), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT23), .Z(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G299), .B2(G16), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT99), .ZN(new_n793));
  INV_X1    g368(.A(G1956), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n789), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n796), .A2(KEYINPUT100), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT100), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n789), .A2(new_n798), .A3(new_n795), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n716), .A2(new_n786), .A3(new_n797), .A4(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT95), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n743), .A2(G22), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G303), .B2(G16), .ZN(new_n803));
  INV_X1    g378(.A(G1971), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(G288), .A2(G16), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT33), .B(G1976), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT93), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n743), .A2(G23), .ZN(new_n809));
  AND3_X1   g384(.A1(new_n806), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n808), .B1(new_n806), .B2(new_n809), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n805), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n743), .A2(G6), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n595), .B2(new_n743), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n814), .A2(KEYINPUT92), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n814), .A2(KEYINPUT92), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT32), .B(G1981), .ZN(new_n817));
  OR3_X1    g392(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n815), .B2(new_n816), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n812), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n820), .A2(KEYINPUT94), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(KEYINPUT94), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT34), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n801), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n821), .A2(KEYINPUT95), .A3(KEYINPUT34), .A4(new_n822), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AND2_X1   g402(.A1(new_n721), .A2(G25), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n488), .A2(new_n489), .ZN(new_n829));
  INV_X1    g404(.A(G119), .ZN(new_n830));
  OAI21_X1  g405(.A(KEYINPUT89), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n832));
  INV_X1    g407(.A(G107), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(G2105), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(G131), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n835), .B1(new_n481), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n830), .B1(new_n488), .B2(new_n489), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT89), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n831), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n828), .B1(new_n841), .B2(G29), .ZN(new_n842));
  XOR2_X1   g417(.A(KEYINPUT35), .B(G1991), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT91), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT90), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n743), .A2(G24), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(G290), .B2(G16), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(G1986), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n842), .A2(new_n845), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI211_X1 g426(.A(new_n846), .B(new_n851), .C1(new_n823), .C2(new_n824), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n827), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(KEYINPUT36), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT36), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n827), .A2(new_n852), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n800), .B1(new_n854), .B2(new_n856), .ZN(G311));
  AND4_X1   g432(.A1(new_n797), .A2(new_n716), .A3(new_n786), .A4(new_n799), .ZN(new_n858));
  INV_X1    g433(.A(new_n856), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n855), .B1(new_n827), .B2(new_n852), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(G150));
  NAND2_X1  g436(.A1(new_n629), .A2(G559), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT38), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n521), .A2(new_n523), .A3(G67), .ZN(new_n864));
  NAND2_X1  g439(.A1(G80), .A2(G543), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n509), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(G55), .ZN(new_n867));
  XNOR2_X1  g442(.A(KEYINPUT101), .B(G93), .ZN(new_n868));
  OAI22_X1  g443(.A1(new_n530), .A2(new_n867), .B1(new_n536), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n565), .A2(new_n871), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n870), .B(new_n560), .C1(new_n564), .C2(new_n563), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n863), .B(new_n874), .Z(new_n875));
  AND2_X1   g450(.A1(new_n875), .A2(KEYINPUT39), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(KEYINPUT39), .ZN(new_n877));
  NOR3_X1   g452(.A1(new_n876), .A2(new_n877), .A3(G860), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n871), .A2(G860), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT102), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n880), .B(KEYINPUT37), .Z(new_n881));
  OR2_X1    g456(.A1(new_n878), .A2(new_n881), .ZN(G145));
  XNOR2_X1  g457(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  XOR2_X1   g459(.A(G162), .B(G160), .Z(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n644), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT105), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n490), .A2(new_n839), .A3(G119), .ZN(new_n889));
  INV_X1    g464(.A(new_n837), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n838), .A2(new_n839), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n888), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n831), .A2(new_n840), .A3(KEYINPUT105), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n498), .A2(new_n501), .A3(KEYINPUT4), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n501), .B1(new_n498), .B2(KEYINPUT4), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n505), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n493), .A2(KEYINPUT103), .A3(new_n495), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT103), .B1(new_n493), .B2(new_n495), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n736), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(G128), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n903), .B1(new_n488), .B2(new_n489), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n897), .B(new_n900), .C1(new_n904), .C2(new_n735), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n893), .A2(new_n894), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n906), .B1(new_n893), .B2(new_n894), .ZN(new_n908));
  INV_X1    g483(.A(new_n648), .ZN(new_n909));
  INV_X1    g484(.A(G130), .ZN(new_n910));
  OAI21_X1  g485(.A(KEYINPUT104), .B1(new_n829), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n912));
  INV_X1    g487(.A(G118), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n912), .B1(new_n913), .B2(G2105), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G142), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n915), .B1(new_n481), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n910), .B1(new_n488), .B2(new_n489), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT104), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n909), .B1(new_n911), .B2(new_n920), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n911), .A2(new_n920), .A3(new_n909), .ZN(new_n922));
  OAI22_X1  g497(.A1(new_n907), .A2(new_n908), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n710), .A2(new_n766), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(new_n711), .B2(new_n766), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n902), .A2(new_n905), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n891), .A2(new_n888), .A3(new_n892), .ZN(new_n927));
  AOI21_X1  g502(.A(KEYINPUT105), .B1(new_n831), .B2(new_n840), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n922), .A2(new_n921), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n893), .A2(new_n894), .A3(new_n906), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n923), .A2(new_n925), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n925), .B1(new_n923), .B2(new_n932), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n887), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n925), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n930), .B1(new_n929), .B2(new_n931), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT106), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n923), .A2(new_n925), .A3(new_n932), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n939), .A2(new_n940), .A3(new_n941), .A4(new_n886), .ZN(new_n942));
  INV_X1    g517(.A(G37), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n935), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n939), .A2(new_n886), .A3(new_n941), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n945), .A2(KEYINPUT106), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n884), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n939), .A2(new_n941), .ZN(new_n948));
  AOI21_X1  g523(.A(G37), .B1(new_n948), .B2(new_n887), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n945), .A2(KEYINPUT106), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n949), .A2(new_n950), .A3(new_n942), .A4(new_n883), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n947), .A2(new_n951), .ZN(G395));
  XNOR2_X1  g527(.A(G288), .B(G303), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n608), .A2(G305), .A3(new_n610), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(G305), .B1(new_n608), .B2(new_n610), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n957), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n959), .A2(new_n953), .A3(new_n955), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n961), .A2(KEYINPUT111), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT42), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n962), .B(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n634), .B(new_n874), .ZN(new_n965));
  XOR2_X1   g540(.A(KEYINPUT109), .B(KEYINPUT41), .Z(new_n966));
  NAND2_X1  g541(.A1(G299), .A2(new_n621), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n573), .A2(new_n619), .A3(new_n577), .A4(new_n620), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT41), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OR3_X1    g548(.A1(new_n965), .A2(KEYINPUT110), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n970), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(KEYINPUT108), .B1(new_n967), .B2(new_n968), .ZN(new_n977));
  OR2_X1    g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n965), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT110), .B1(new_n965), .B2(new_n973), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n974), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT112), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT112), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n974), .B(new_n983), .C1(new_n979), .C2(new_n980), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n964), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n964), .A2(new_n984), .ZN(new_n986));
  OAI21_X1  g561(.A(G868), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n987), .B1(G868), .B2(new_n870), .ZN(G295));
  OAI21_X1  g563(.A(new_n987), .B1(G868), .B2(new_n870), .ZN(G331));
  AND3_X1   g564(.A1(new_n545), .A2(KEYINPUT77), .A3(new_n546), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT77), .B1(new_n545), .B2(new_n546), .ZN(new_n991));
  NOR3_X1   g566(.A1(new_n990), .A2(new_n991), .A3(new_n509), .ZN(new_n992));
  INV_X1    g567(.A(new_n553), .ZN(new_n993));
  OAI21_X1  g568(.A(G286), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n535), .A2(new_n542), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n551), .A2(new_n995), .A3(new_n534), .A4(new_n553), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n997), .A2(new_n874), .ZN(new_n998));
  AOI22_X1  g573(.A1(new_n994), .A2(new_n996), .B1(new_n872), .B2(new_n873), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n970), .A2(new_n972), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1001), .B1(new_n970), .B2(new_n966), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(KEYINPUT114), .B1(new_n998), .B2(new_n999), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n997), .A2(new_n874), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1004), .A2(new_n978), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1003), .B1(new_n1008), .B2(KEYINPUT115), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n994), .A2(new_n996), .A3(new_n872), .A4(new_n873), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1006), .B1(new_n1005), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n976), .A2(new_n977), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n999), .A2(KEYINPUT114), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT115), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1009), .A2(new_n1016), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n958), .A2(new_n960), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT43), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n998), .A2(new_n999), .A3(new_n970), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n961), .B(new_n1022), .C1(new_n1023), .C2(new_n973), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n943), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1019), .A2(new_n1020), .A3(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n973), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1018), .B1(new_n1028), .B2(new_n1021), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT43), .B1(new_n1030), .B2(new_n1025), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1027), .A2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT113), .B(KEYINPUT44), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1029), .A2(new_n1024), .A3(new_n1020), .A4(new_n943), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n1035), .A2(KEYINPUT44), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n961), .B1(new_n1009), .B2(new_n1016), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT43), .B1(new_n1038), .B2(new_n1025), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n1036), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1037), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1034), .B1(new_n1040), .B2(new_n1041), .ZN(G397));
  INV_X1    g617(.A(G1384), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT45), .B1(new_n901), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G40), .ZN(new_n1045));
  AOI211_X1 g620(.A(new_n1045), .B(new_n467), .C1(new_n477), .C2(new_n462), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n841), .A2(new_n844), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n841), .A2(new_n844), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1048), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n736), .B(new_n738), .ZN(new_n1052));
  INV_X1    g627(.A(G1996), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n710), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1048), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1048), .A2(KEYINPUT117), .A3(new_n1053), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1057), .B1(new_n1047), .B2(G1996), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n711), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1060), .A2(KEYINPUT118), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1060), .A2(KEYINPUT118), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1051), .B(new_n1055), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g638(.A(G290), .B(G1986), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1063), .B1(new_n1048), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(G160), .A2(G40), .ZN(new_n1066));
  AOI21_X1  g641(.A(G1384), .B1(new_n897), .B2(new_n900), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT50), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n505), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1070), .B1(new_n500), .B2(new_n502), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1043), .B1(new_n1071), .B2(new_n496), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT50), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1069), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1961), .ZN(new_n1075));
  INV_X1    g650(.A(G2078), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT53), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1044), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT45), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1079), .A2(G1384), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1066), .B1(new_n901), .B2(new_n1080), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1074), .A2(new_n1075), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1072), .A2(new_n1079), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1083), .A2(new_n1081), .A3(new_n1076), .ZN(new_n1084));
  XNOR2_X1  g659(.A(KEYINPUT125), .B(KEYINPUT53), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1084), .A2(KEYINPUT126), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT126), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1087));
  OAI211_X1 g662(.A(G301), .B(new_n1082), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1044), .ZN(new_n1089));
  INV_X1    g664(.A(new_n496), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n897), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1066), .B1(new_n1091), .B2(new_n1080), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1077), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1089), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n899), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n493), .A2(KEYINPUT103), .A3(new_n495), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1068), .B(new_n1043), .C1(new_n1071), .C2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n1046), .ZN(new_n1099));
  AOI21_X1  g674(.A(G1384), .B1(new_n897), .B2(new_n1090), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1100), .A2(new_n1068), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1075), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1094), .A2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1080), .B1(new_n1071), .B2(new_n1097), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1104), .B(new_n1046), .C1(new_n1100), .C2(KEYINPUT45), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1085), .B1(new_n1105), .B2(G2078), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT126), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1084), .A2(KEYINPUT126), .A3(new_n1085), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1103), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1088), .B1(new_n1110), .B2(G301), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT54), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n1114));
  INV_X1    g689(.A(G1966), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1080), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1046), .B1(G164), .B2(new_n1116), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1114), .B(new_n1115), .C1(new_n1117), .C2(new_n1044), .ZN(new_n1118));
  INV_X1    g693(.A(G2084), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1069), .A2(new_n1119), .A3(new_n1073), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1092), .B1(KEYINPUT45), .B2(new_n1067), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1114), .B1(new_n1122), .B2(new_n1115), .ZN(new_n1123));
  OAI21_X1  g698(.A(G8), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(G286), .A2(G8), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT51), .B1(new_n1125), .B2(KEYINPUT124), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1124), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1115), .B1(new_n1117), .B2(new_n1044), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT119), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1130), .A2(new_n1120), .A3(new_n1118), .ZN(new_n1131));
  OAI211_X1 g706(.A(G8), .B(new_n1126), .C1(new_n1131), .C2(G286), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1131), .A2(G8), .A3(G286), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1128), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1094), .A2(new_n1102), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1135), .B(G301), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(new_n1102), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1138), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1136), .B(KEYINPUT54), .C1(new_n1139), .C2(G301), .ZN(new_n1140));
  NAND2_X1  g715(.A1(G303), .A2(G8), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n1141), .B(KEYINPUT55), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n1099), .A2(new_n1101), .A3(G2090), .ZN(new_n1144));
  AOI21_X1  g719(.A(G1971), .B1(new_n1083), .B2(new_n1081), .ZN(new_n1145));
  OAI211_X1 g720(.A(G8), .B(new_n1143), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n901), .A2(new_n1043), .A3(new_n1046), .ZN(new_n1147));
  INV_X1    g722(.A(G288), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(G1976), .ZN(new_n1149));
  INV_X1    g724(.A(G1976), .ZN(new_n1150));
  AOI21_X1  g725(.A(KEYINPUT52), .B1(G288), .B2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1147), .A2(G8), .A3(new_n1149), .A4(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(G1981), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n590), .A2(new_n591), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1153), .B(new_n586), .C1(new_n1154), .C2(new_n593), .ZN(new_n1155));
  OAI21_X1  g730(.A(G1981), .B1(new_n587), .B2(new_n590), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT49), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1155), .A2(new_n1156), .A3(KEYINPUT49), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1147), .A2(new_n1159), .A3(G8), .A4(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1152), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT52), .ZN(new_n1163));
  INV_X1    g738(.A(G8), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1164), .B1(new_n1067), .B2(new_n1046), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1163), .B1(new_n1165), .B2(new_n1149), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1162), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1066), .B1(new_n1100), .B2(new_n1068), .ZN(new_n1168));
  INV_X1    g743(.A(G2090), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1168), .B(new_n1169), .C1(new_n1068), .C2(new_n1067), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1105), .A2(new_n804), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1164), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n1146), .B(new_n1167), .C1(new_n1143), .C2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1173), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1113), .A2(new_n1134), .A3(new_n1140), .A4(new_n1174), .ZN(new_n1175));
  XOR2_X1   g750(.A(KEYINPUT58), .B(G1341), .Z(new_n1176));
  NAND2_X1  g751(.A1(new_n1147), .A2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1177), .B1(new_n1105), .B2(G1996), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(new_n566), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT59), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n1179), .B(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g756(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n1182));
  INV_X1    g757(.A(G2072), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1182), .B(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(KEYINPUT122), .B1(new_n1105), .B2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1046), .B1(new_n1072), .B2(KEYINPUT50), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n794), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT122), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1083), .A2(new_n1081), .A3(new_n1190), .A4(new_n1184), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1186), .A2(new_n1189), .A3(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g767(.A(G299), .B(KEYINPUT57), .ZN(new_n1193));
  AND2_X1   g768(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1181), .B1(new_n1196), .B2(KEYINPUT61), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT123), .ZN(new_n1198));
  AOI21_X1  g773(.A(G1348), .B1(new_n1069), .B2(new_n1073), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1147), .A2(G2067), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1198), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n719), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1200), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1202), .A2(new_n1203), .A3(KEYINPUT123), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1201), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n621), .B1(new_n1205), .B2(KEYINPUT60), .ZN(new_n1206));
  INV_X1    g781(.A(KEYINPUT60), .ZN(new_n1207));
  AOI211_X1 g782(.A(new_n1207), .B(new_n629), .C1(new_n1201), .C2(new_n1204), .ZN(new_n1208));
  OAI22_X1  g783(.A1(new_n1206), .A2(new_n1208), .B1(KEYINPUT60), .B2(new_n1205), .ZN(new_n1209));
  INV_X1    g784(.A(KEYINPUT61), .ZN(new_n1210));
  OAI21_X1  g785(.A(new_n1210), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1197), .A2(new_n1209), .A3(new_n1211), .ZN(new_n1212));
  NOR3_X1   g787(.A1(new_n1195), .A2(new_n1205), .A3(new_n621), .ZN(new_n1213));
  NOR2_X1   g788(.A1(new_n1213), .A2(new_n1194), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1175), .B1(new_n1212), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1134), .A2(KEYINPUT62), .ZN(new_n1216));
  INV_X1    g791(.A(KEYINPUT62), .ZN(new_n1217));
  NAND4_X1  g792(.A1(new_n1128), .A2(new_n1132), .A3(new_n1217), .A4(new_n1133), .ZN(new_n1218));
  NOR3_X1   g793(.A1(new_n1173), .A2(G301), .A3(new_n1110), .ZN(new_n1219));
  NAND3_X1  g794(.A1(new_n1216), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  NAND3_X1  g795(.A1(new_n1069), .A2(new_n1169), .A3(new_n1073), .ZN(new_n1221));
  AOI21_X1  g796(.A(new_n1164), .B1(new_n1171), .B2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g797(.A1(new_n1167), .A2(new_n1222), .A3(new_n1143), .ZN(new_n1223));
  AND3_X1   g798(.A1(new_n1161), .A2(new_n1150), .A3(new_n1148), .ZN(new_n1224));
  INV_X1    g799(.A(new_n1155), .ZN(new_n1225));
  OAI21_X1  g800(.A(new_n1165), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1223), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1146), .A2(KEYINPUT63), .ZN(new_n1228));
  OAI211_X1 g803(.A(G8), .B(G168), .C1(new_n1121), .C2(new_n1123), .ZN(new_n1229));
  NOR2_X1   g804(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g805(.A(G8), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n1231), .A2(new_n1142), .ZN(new_n1232));
  AOI21_X1  g807(.A(KEYINPUT120), .B1(new_n1232), .B2(new_n1167), .ZN(new_n1233));
  OAI211_X1 g808(.A(new_n1167), .B(KEYINPUT120), .C1(new_n1222), .C2(new_n1143), .ZN(new_n1234));
  INV_X1    g809(.A(new_n1234), .ZN(new_n1235));
  OAI21_X1  g810(.A(new_n1230), .B1(new_n1233), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g811(.A(KEYINPUT63), .ZN(new_n1237));
  OAI21_X1  g812(.A(new_n1237), .B1(new_n1173), .B2(new_n1229), .ZN(new_n1238));
  AOI21_X1  g813(.A(new_n1227), .B1(new_n1236), .B2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g814(.A1(new_n1220), .A2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g815(.A(new_n1065), .B1(new_n1215), .B2(new_n1240), .ZN(new_n1241));
  AND3_X1   g816(.A1(new_n1056), .A2(KEYINPUT46), .A3(new_n1058), .ZN(new_n1242));
  AOI21_X1  g817(.A(KEYINPUT46), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1243));
  OR2_X1    g818(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g819(.A(KEYINPUT47), .ZN(new_n1245));
  INV_X1    g820(.A(new_n710), .ZN(new_n1246));
  OAI21_X1  g821(.A(new_n1048), .B1(new_n1052), .B2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g822(.A1(new_n1244), .A2(new_n1245), .A3(new_n1247), .ZN(new_n1248));
  INV_X1    g823(.A(new_n1248), .ZN(new_n1249));
  AOI21_X1  g824(.A(new_n1245), .B1(new_n1244), .B2(new_n1247), .ZN(new_n1250));
  NOR3_X1   g825(.A1(G290), .A2(new_n1047), .A3(G1986), .ZN(new_n1251));
  XNOR2_X1  g826(.A(new_n1251), .B(KEYINPUT48), .ZN(new_n1252));
  OAI22_X1  g827(.A1(new_n1249), .A2(new_n1250), .B1(new_n1063), .B2(new_n1252), .ZN(new_n1253));
  OAI211_X1 g828(.A(new_n1050), .B(new_n1055), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1254));
  NAND2_X1  g829(.A1(new_n736), .A2(new_n738), .ZN(new_n1255));
  AOI21_X1  g830(.A(new_n1047), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  NOR2_X1   g831(.A1(new_n1253), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g832(.A1(new_n1241), .A2(new_n1257), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g833(.A(G319), .ZN(new_n1260));
  NOR3_X1   g834(.A1(G401), .A2(G227), .A3(new_n1260), .ZN(new_n1261));
  NAND3_X1  g835(.A1(new_n702), .A2(new_n703), .A3(new_n1261), .ZN(new_n1262));
  AOI21_X1  g836(.A(new_n1262), .B1(new_n1027), .B2(new_n1031), .ZN(new_n1263));
  NAND3_X1  g837(.A1(new_n949), .A2(new_n950), .A3(new_n942), .ZN(new_n1264));
  NAND2_X1  g838(.A1(new_n1263), .A2(new_n1264), .ZN(G225));
  INV_X1    g839(.A(G225), .ZN(G308));
endmodule


