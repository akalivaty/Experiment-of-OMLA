

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727;

  NOR2_X1 U366 ( .A1(n684), .A2(G902), .ZN(n456) );
  XNOR2_X1 U367 ( .A(n363), .B(n475), .ZN(n695) );
  AND2_X4 U368 ( .A1(n611), .A2(n610), .ZN(n690) );
  XNOR2_X2 U369 ( .A(n578), .B(KEYINPUT1), .ZN(n633) );
  INV_X2 U370 ( .A(n364), .ZN(n474) );
  XNOR2_X2 U371 ( .A(G119), .B(G110), .ZN(n364) );
  INV_X1 U372 ( .A(n633), .ZN(n559) );
  NOR2_X1 U373 ( .A1(n678), .A2(n680), .ZN(n628) );
  INV_X1 U374 ( .A(KEYINPUT22), .ZN(n374) );
  INV_X4 U375 ( .A(G953), .ZN(n715) );
  XNOR2_X1 U376 ( .A(G143), .B(G128), .ZN(n402) );
  XNOR2_X1 U377 ( .A(n522), .B(n521), .ZN(n723) );
  NOR2_X1 U378 ( .A1(n451), .A2(n507), .ZN(n662) );
  NAND2_X1 U379 ( .A1(n388), .A2(n387), .ZN(n522) );
  NOR2_X1 U380 ( .A1(n410), .A2(n344), .ZN(n408) );
  AND2_X1 U381 ( .A1(n520), .A2(n547), .ZN(n387) );
  NAND2_X1 U382 ( .A1(n572), .A2(n391), .ZN(n390) );
  XNOR2_X1 U383 ( .A(n356), .B(KEYINPUT67), .ZN(n632) );
  BUF_X1 U384 ( .A(n636), .Z(n451) );
  XNOR2_X1 U385 ( .A(n506), .B(n367), .ZN(n533) );
  XNOR2_X1 U386 ( .A(n400), .B(G146), .ZN(n469) );
  XNOR2_X1 U387 ( .A(n402), .B(n401), .ZN(n471) );
  INV_X1 U388 ( .A(KEYINPUT4), .ZN(n400) );
  XNOR2_X1 U389 ( .A(n448), .B(n426), .ZN(n636) );
  XNOR2_X1 U390 ( .A(n695), .B(n477), .ZN(n612) );
  XNOR2_X1 U391 ( .A(n473), .B(n472), .ZN(n477) );
  XNOR2_X1 U392 ( .A(n399), .B(n396), .ZN(n473) );
  OR2_X1 U393 ( .A1(G902), .A2(G237), .ZN(n483) );
  NOR2_X1 U394 ( .A1(G953), .A2(G237), .ZN(n489) );
  XNOR2_X1 U395 ( .A(n457), .B(G113), .ZN(n476) );
  XNOR2_X1 U396 ( .A(G101), .B(KEYINPUT3), .ZN(n457) );
  XNOR2_X1 U397 ( .A(n471), .B(G134), .ZN(n502) );
  OR2_X1 U398 ( .A1(n661), .A2(G902), .ZN(n413) );
  NOR2_X1 U399 ( .A1(n533), .A2(n532), .ZN(n572) );
  XNOR2_X1 U400 ( .A(n493), .B(n372), .ZN(n687) );
  XNOR2_X1 U401 ( .A(n495), .B(n373), .ZN(n372) );
  INV_X1 U402 ( .A(G113), .ZN(n373) );
  XNOR2_X1 U403 ( .A(n502), .B(n453), .ZN(n707) );
  XNOR2_X1 U404 ( .A(n469), .B(n452), .ZN(n453) );
  XOR2_X1 U405 ( .A(G137), .B(G131), .Z(n452) );
  NAND2_X1 U406 ( .A1(n690), .A2(G472), .ZN(n395) );
  XNOR2_X1 U407 ( .A(KEYINPUT20), .B(n449), .ZN(n460) );
  XNOR2_X1 U408 ( .A(n381), .B(n516), .ZN(n380) );
  INV_X1 U409 ( .A(KEYINPUT16), .ZN(n358) );
  XOR2_X1 U410 ( .A(G122), .B(G104), .Z(n494) );
  XOR2_X1 U411 ( .A(G116), .B(G107), .Z(n501) );
  NOR2_X1 U412 ( .A1(n636), .A2(n635), .ZN(n356) );
  XNOR2_X1 U413 ( .A(n414), .B(n707), .ZN(n661) );
  XNOR2_X1 U414 ( .A(n459), .B(n348), .ZN(n414) );
  XNOR2_X1 U415 ( .A(n361), .B(n476), .ZN(n459) );
  NOR2_X1 U416 ( .A1(n407), .A2(n571), .ZN(n406) );
  XNOR2_X1 U417 ( .A(n360), .B(n359), .ZN(n557) );
  INV_X1 U418 ( .A(KEYINPUT104), .ZN(n359) );
  NOR2_X1 U419 ( .A1(n550), .A2(n549), .ZN(n360) );
  INV_X1 U420 ( .A(KEYINPUT85), .ZN(n479) );
  INV_X1 U421 ( .A(G478), .ZN(n367) );
  XNOR2_X1 U422 ( .A(n497), .B(n496), .ZN(n532) );
  NAND2_X1 U423 ( .A1(n608), .A2(n607), .ZN(n611) );
  XNOR2_X1 U424 ( .A(n707), .B(n346), .ZN(n684) );
  XNOR2_X1 U425 ( .A(n368), .B(n345), .ZN(n428) );
  XNOR2_X1 U426 ( .A(n614), .B(n613), .ZN(n615) );
  NOR2_X1 U427 ( .A1(n725), .A2(n726), .ZN(n583) );
  XNOR2_X1 U428 ( .A(KEYINPUT92), .B(n462), .ZN(n635) );
  XNOR2_X1 U429 ( .A(n458), .B(G116), .ZN(n361) );
  XOR2_X1 U430 ( .A(KEYINPUT5), .B(G119), .Z(n458) );
  INV_X1 U431 ( .A(KEYINPUT98), .ZN(n377) );
  XNOR2_X1 U432 ( .A(KEYINPUT11), .B(KEYINPUT94), .ZN(n487) );
  INV_X1 U433 ( .A(n478), .ZN(n605) );
  XNOR2_X1 U434 ( .A(n469), .B(n470), .ZN(n399) );
  XNOR2_X1 U435 ( .A(n468), .B(n397), .ZN(n396) );
  XNOR2_X1 U436 ( .A(G125), .B(KEYINPUT84), .ZN(n468) );
  XNOR2_X1 U437 ( .A(n398), .B(KEYINPUT18), .ZN(n397) );
  INV_X1 U438 ( .A(KEYINPUT17), .ZN(n398) );
  INV_X1 U439 ( .A(KEYINPUT65), .ZN(n401) );
  XOR2_X1 U440 ( .A(KEYINPUT15), .B(G902), .Z(n478) );
  XNOR2_X1 U441 ( .A(n450), .B(n447), .ZN(n426) );
  INV_X1 U442 ( .A(n635), .ZN(n391) );
  XNOR2_X1 U443 ( .A(n476), .B(n357), .ZN(n363) );
  XNOR2_X1 U444 ( .A(n474), .B(n358), .ZN(n357) );
  XOR2_X1 U445 ( .A(KEYINPUT23), .B(KEYINPUT88), .Z(n440) );
  XNOR2_X1 U446 ( .A(G128), .B(G137), .ZN(n439) );
  XNOR2_X1 U447 ( .A(n706), .B(G146), .ZN(n492) );
  XNOR2_X1 U448 ( .A(n355), .B(n474), .ZN(n436) );
  XNOR2_X1 U449 ( .A(n431), .B(KEYINPUT89), .ZN(n355) );
  XNOR2_X1 U450 ( .A(KEYINPUT24), .B(KEYINPUT90), .ZN(n431) );
  XOR2_X1 U451 ( .A(KEYINPUT7), .B(G122), .Z(n504) );
  NOR2_X1 U452 ( .A1(n609), .A2(n701), .ZN(n620) );
  XNOR2_X1 U453 ( .A(n454), .B(n369), .ZN(n368) );
  XNOR2_X1 U454 ( .A(G107), .B(G104), .ZN(n454) );
  XNOR2_X1 U455 ( .A(n574), .B(n573), .ZN(n655) );
  XNOR2_X1 U456 ( .A(n383), .B(n511), .ZN(n643) );
  INV_X1 U457 ( .A(KEYINPUT93), .ZN(n511) );
  NAND2_X1 U458 ( .A1(n527), .A2(n384), .ZN(n383) );
  NOR2_X1 U459 ( .A1(n633), .A2(n514), .ZN(n384) );
  XNOR2_X1 U460 ( .A(n563), .B(n412), .ZN(n411) );
  INV_X1 U461 ( .A(KEYINPUT30), .ZN(n412) );
  BUF_X1 U462 ( .A(n633), .Z(n365) );
  XNOR2_X1 U463 ( .A(n687), .B(n686), .ZN(n688) );
  XNOR2_X1 U464 ( .A(n561), .B(KEYINPUT109), .ZN(n720) );
  NOR2_X1 U465 ( .A1(n508), .A2(n533), .ZN(n678) );
  NAND2_X1 U466 ( .A1(n394), .A2(n423), .ZN(n393) );
  XNOR2_X1 U467 ( .A(n395), .B(n350), .ZN(n394) );
  XNOR2_X1 U468 ( .A(n386), .B(n385), .ZN(n685) );
  NAND2_X1 U469 ( .A1(n424), .A2(n423), .ZN(n422) );
  XNOR2_X1 U470 ( .A(n425), .B(n615), .ZN(n424) );
  XNOR2_X1 U471 ( .A(n660), .B(KEYINPUT117), .ZN(n404) );
  INV_X1 U472 ( .A(n547), .ZN(n418) );
  INV_X1 U473 ( .A(n628), .ZN(n382) );
  AND2_X1 U474 ( .A1(n409), .A2(KEYINPUT39), .ZN(n344) );
  XOR2_X1 U475 ( .A(G110), .B(G101), .Z(n345) );
  XOR2_X1 U476 ( .A(n428), .B(n455), .Z(n346) );
  XOR2_X1 U477 ( .A(KEYINPUT38), .B(n568), .Z(n571) );
  OR2_X1 U478 ( .A1(n677), .A2(n664), .ZN(n347) );
  AND2_X1 U479 ( .A1(n489), .A2(G210), .ZN(n348) );
  INV_X1 U480 ( .A(G140), .ZN(n369) );
  XNOR2_X1 U481 ( .A(KEYINPUT33), .B(KEYINPUT69), .ZN(n349) );
  XOR2_X1 U482 ( .A(n661), .B(KEYINPUT62), .Z(n350) );
  NOR2_X1 U483 ( .A1(G952), .A2(n715), .ZN(n694) );
  INV_X1 U484 ( .A(n694), .ZN(n423) );
  XNOR2_X1 U485 ( .A(KEYINPUT63), .B(KEYINPUT110), .ZN(n351) );
  XOR2_X1 U486 ( .A(KEYINPUT66), .B(KEYINPUT60), .Z(n352) );
  XOR2_X1 U487 ( .A(KEYINPUT118), .B(KEYINPUT53), .Z(n353) );
  XOR2_X1 U488 ( .A(KEYINPUT80), .B(KEYINPUT56), .Z(n354) );
  NOR2_X1 U489 ( .A1(n601), .A2(n724), .ZN(n603) );
  NOR2_X1 U490 ( .A1(n632), .A2(n578), .ZN(n566) );
  NAND2_X1 U491 ( .A1(n690), .A2(G210), .ZN(n425) );
  XNOR2_X1 U492 ( .A(n362), .B(n539), .ZN(n415) );
  NAND2_X1 U493 ( .A1(n416), .A2(n722), .ZN(n362) );
  XNOR2_X1 U494 ( .A(n366), .B(n505), .ZN(n617) );
  XNOR2_X1 U495 ( .A(n503), .B(n504), .ZN(n366) );
  NAND2_X1 U496 ( .A1(n380), .A2(n379), .ZN(n378) );
  XNOR2_X2 U497 ( .A(n456), .B(G469), .ZN(n578) );
  XNOR2_X2 U498 ( .A(n370), .B(n540), .ZN(n701) );
  NAND2_X1 U499 ( .A1(n415), .A2(n430), .ZN(n370) );
  XNOR2_X1 U500 ( .A(n371), .B(n352), .ZN(G60) );
  NAND2_X1 U501 ( .A1(n420), .A2(n423), .ZN(n371) );
  XNOR2_X1 U502 ( .A(n490), .B(n427), .ZN(n491) );
  XNOR2_X1 U503 ( .A(n421), .B(n688), .ZN(n420) );
  NAND2_X1 U504 ( .A1(n404), .A2(n715), .ZN(n403) );
  XNOR2_X1 U505 ( .A(n403), .B(n353), .ZN(G75) );
  XNOR2_X2 U506 ( .A(n375), .B(n374), .ZN(n524) );
  NOR2_X2 U507 ( .A1(n529), .A2(n390), .ZN(n375) );
  XNOR2_X1 U508 ( .A(n378), .B(n377), .ZN(n518) );
  XNOR2_X1 U509 ( .A(n616), .B(n376), .ZN(n618) );
  INV_X1 U510 ( .A(n617), .ZN(n376) );
  INV_X1 U511 ( .A(n662), .ZN(n379) );
  NAND2_X1 U512 ( .A1(n347), .A2(n382), .ZN(n381) );
  XNOR2_X1 U513 ( .A(n684), .B(n683), .ZN(n385) );
  NAND2_X1 U514 ( .A1(n690), .A2(G469), .ZN(n386) );
  NOR2_X1 U515 ( .A1(n524), .A2(n418), .ZN(n389) );
  INV_X1 U516 ( .A(n524), .ZN(n388) );
  NAND2_X1 U517 ( .A1(n389), .A2(n365), .ZN(n507) );
  XNOR2_X2 U518 ( .A(n392), .B(KEYINPUT0), .ZN(n529) );
  NAND2_X1 U519 ( .A1(n485), .A2(n486), .ZN(n392) );
  XNOR2_X1 U520 ( .A(n393), .B(n351), .ZN(G57) );
  NAND2_X1 U521 ( .A1(n411), .A2(n567), .ZN(n590) );
  NAND2_X1 U522 ( .A1(n408), .A2(n405), .ZN(n602) );
  NAND2_X1 U523 ( .A1(n411), .A2(n406), .ZN(n405) );
  NAND2_X1 U524 ( .A1(n567), .A2(n569), .ZN(n407) );
  NAND2_X1 U525 ( .A1(n624), .A2(n567), .ZN(n409) );
  NOR2_X1 U526 ( .A1(n411), .A2(n569), .ZN(n410) );
  XNOR2_X2 U527 ( .A(n413), .B(G472), .ZN(n639) );
  XNOR2_X1 U528 ( .A(n526), .B(KEYINPUT81), .ZN(n416) );
  XNOR2_X1 U529 ( .A(n537), .B(KEYINPUT35), .ZN(n722) );
  NOR2_X1 U530 ( .A1(n654), .A2(n529), .ZN(n531) );
  XNOR2_X2 U531 ( .A(n417), .B(n349), .ZN(n654) );
  NAND2_X1 U532 ( .A1(n419), .A2(n418), .ZN(n417) );
  XNOR2_X1 U533 ( .A(n528), .B(KEYINPUT101), .ZN(n419) );
  NAND2_X1 U534 ( .A1(n690), .A2(G475), .ZN(n421) );
  XNOR2_X1 U535 ( .A(n422), .B(n354), .ZN(G51) );
  XNOR2_X1 U536 ( .A(n556), .B(n484), .ZN(n585) );
  XNOR2_X1 U537 ( .A(n639), .B(KEYINPUT6), .ZN(n547) );
  AND2_X1 U538 ( .A1(n489), .A2(G214), .ZN(n427) );
  AND2_X1 U539 ( .A1(n598), .A2(n597), .ZN(n429) );
  AND2_X1 U540 ( .A1(n518), .A2(n517), .ZN(n430) );
  XNOR2_X1 U541 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n582) );
  XNOR2_X1 U542 ( .A(n583), .B(n582), .ZN(n598) );
  XNOR2_X1 U543 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U544 ( .A(n442), .B(n441), .ZN(n443) );
  NAND2_X1 U545 ( .A1(n593), .A2(n623), .ZN(n556) );
  XNOR2_X1 U546 ( .A(n480), .B(n479), .ZN(n481) );
  NAND2_X1 U547 ( .A1(n618), .A2(n423), .ZN(n619) );
  XNOR2_X1 U548 ( .A(n619), .B(KEYINPUT119), .ZN(G63) );
  XNOR2_X2 U549 ( .A(G125), .B(KEYINPUT10), .ZN(n433) );
  INV_X1 U550 ( .A(n433), .ZN(n432) );
  NAND2_X1 U551 ( .A1(G140), .A2(n432), .ZN(n435) );
  NAND2_X1 U552 ( .A1(n369), .A2(n433), .ZN(n434) );
  NAND2_X1 U553 ( .A1(n435), .A2(n434), .ZN(n706) );
  XNOR2_X1 U554 ( .A(n436), .B(n492), .ZN(n444) );
  XOR2_X1 U555 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n438) );
  NAND2_X1 U556 ( .A1(G234), .A2(n715), .ZN(n437) );
  XNOR2_X1 U557 ( .A(n438), .B(n437), .ZN(n498) );
  NAND2_X1 U558 ( .A1(G221), .A2(n498), .ZN(n442) );
  XNOR2_X1 U559 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U560 ( .A(n444), .B(n443), .ZN(n689) );
  NOR2_X1 U561 ( .A1(G902), .A2(n689), .ZN(n448) );
  XNOR2_X1 U562 ( .A(KEYINPUT25), .B(KEYINPUT73), .ZN(n446) );
  INV_X1 U563 ( .A(KEYINPUT91), .ZN(n445) );
  NAND2_X1 U564 ( .A1(G234), .A2(n605), .ZN(n449) );
  NAND2_X1 U565 ( .A1(n460), .A2(G217), .ZN(n450) );
  NAND2_X1 U566 ( .A1(G227), .A2(n715), .ZN(n455) );
  NAND2_X1 U567 ( .A1(n460), .A2(G221), .ZN(n461) );
  XNOR2_X1 U568 ( .A(n461), .B(KEYINPUT21), .ZN(n462) );
  NAND2_X1 U569 ( .A1(G237), .A2(G234), .ZN(n463) );
  XNOR2_X1 U570 ( .A(n463), .B(KEYINPUT14), .ZN(n465) );
  NAND2_X1 U571 ( .A1(G952), .A2(n465), .ZN(n653) );
  NOR2_X1 U572 ( .A1(G953), .A2(n653), .ZN(n545) );
  NOR2_X1 U573 ( .A1(G898), .A2(n715), .ZN(n464) );
  XOR2_X1 U574 ( .A(KEYINPUT86), .B(n464), .Z(n696) );
  NAND2_X1 U575 ( .A1(G902), .A2(n465), .ZN(n542) );
  NOR2_X1 U576 ( .A1(n696), .A2(n542), .ZN(n466) );
  NOR2_X1 U577 ( .A1(n545), .A2(n466), .ZN(n467) );
  XNOR2_X1 U578 ( .A(KEYINPUT87), .B(n467), .ZN(n486) );
  AND2_X1 U579 ( .A1(G224), .A2(n715), .ZN(n470) );
  INV_X1 U580 ( .A(n471), .ZN(n472) );
  XNOR2_X1 U581 ( .A(n501), .B(n494), .ZN(n475) );
  NOR2_X2 U582 ( .A1(n612), .A2(n478), .ZN(n482) );
  NAND2_X1 U583 ( .A1(G210), .A2(n483), .ZN(n480) );
  XNOR2_X2 U584 ( .A(n482), .B(n481), .ZN(n593) );
  NAND2_X1 U585 ( .A1(G214), .A2(n483), .ZN(n623) );
  INV_X1 U586 ( .A(KEYINPUT19), .ZN(n484) );
  INV_X1 U587 ( .A(n585), .ZN(n485) );
  XNOR2_X1 U588 ( .A(KEYINPUT13), .B(G475), .ZN(n497) );
  XOR2_X1 U589 ( .A(G131), .B(KEYINPUT12), .Z(n488) );
  XNOR2_X1 U590 ( .A(n488), .B(n487), .ZN(n490) );
  XNOR2_X1 U591 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U592 ( .A(n494), .B(G143), .ZN(n495) );
  NOR2_X1 U593 ( .A1(G902), .A2(n687), .ZN(n496) );
  XOR2_X1 U594 ( .A(KEYINPUT9), .B(KEYINPUT95), .Z(n500) );
  NAND2_X1 U595 ( .A1(G217), .A2(n498), .ZN(n499) );
  XNOR2_X1 U596 ( .A(n500), .B(n499), .ZN(n505) );
  XNOR2_X1 U597 ( .A(n502), .B(n501), .ZN(n503) );
  NOR2_X1 U598 ( .A1(G902), .A2(n617), .ZN(n506) );
  INV_X1 U599 ( .A(KEYINPUT97), .ZN(n516) );
  INV_X1 U600 ( .A(n532), .ZN(n508) );
  INV_X1 U601 ( .A(n533), .ZN(n509) );
  NOR2_X1 U602 ( .A1(n509), .A2(n532), .ZN(n510) );
  XNOR2_X1 U603 ( .A(n510), .B(KEYINPUT96), .ZN(n680) );
  INV_X1 U604 ( .A(n632), .ZN(n527) );
  NOR2_X1 U605 ( .A1(n529), .A2(n643), .ZN(n513) );
  INV_X1 U606 ( .A(KEYINPUT31), .ZN(n512) );
  XNOR2_X1 U607 ( .A(n513), .B(n512), .ZN(n677) );
  INV_X1 U608 ( .A(n639), .ZN(n514) );
  NAND2_X1 U609 ( .A1(n566), .A2(n514), .ZN(n515) );
  NOR2_X1 U610 ( .A1(n529), .A2(n515), .ZN(n664) );
  INV_X1 U611 ( .A(KEYINPUT70), .ZN(n538) );
  NAND2_X1 U612 ( .A1(n538), .A2(KEYINPUT44), .ZN(n517) );
  NAND2_X1 U613 ( .A1(n451), .A2(n559), .ZN(n519) );
  XNOR2_X1 U614 ( .A(KEYINPUT99), .B(n519), .ZN(n520) );
  XNOR2_X1 U615 ( .A(KEYINPUT76), .B(KEYINPUT32), .ZN(n521) );
  XNOR2_X1 U616 ( .A(KEYINPUT100), .B(n639), .ZN(n562) );
  INV_X1 U617 ( .A(n562), .ZN(n576) );
  NAND2_X1 U618 ( .A1(n365), .A2(n576), .ZN(n523) );
  NOR2_X1 U619 ( .A1(n524), .A2(n523), .ZN(n525) );
  NAND2_X1 U620 ( .A1(n451), .A2(n525), .ZN(n668) );
  NAND2_X1 U621 ( .A1(n723), .A2(n668), .ZN(n526) );
  NAND2_X1 U622 ( .A1(n559), .A2(n527), .ZN(n528) );
  XNOR2_X1 U623 ( .A(KEYINPUT34), .B(KEYINPUT75), .ZN(n530) );
  XNOR2_X1 U624 ( .A(n531), .B(n530), .ZN(n536) );
  NAND2_X1 U625 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U626 ( .A(n534), .B(KEYINPUT102), .ZN(n591) );
  XNOR2_X1 U627 ( .A(KEYINPUT74), .B(n591), .ZN(n535) );
  NOR2_X1 U628 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U629 ( .A1(n538), .A2(KEYINPUT44), .ZN(n539) );
  INV_X1 U630 ( .A(KEYINPUT45), .ZN(n540) );
  NOR2_X2 U631 ( .A1(n701), .A2(n605), .ZN(n541) );
  XNOR2_X1 U632 ( .A(n541), .B(KEYINPUT78), .ZN(n604) );
  INV_X1 U633 ( .A(n593), .ZN(n568) );
  OR2_X1 U634 ( .A1(n715), .A2(n542), .ZN(n543) );
  NOR2_X1 U635 ( .A1(G900), .A2(n543), .ZN(n544) );
  NOR2_X1 U636 ( .A1(n545), .A2(n544), .ZN(n564) );
  NOR2_X1 U637 ( .A1(n564), .A2(n635), .ZN(n546) );
  NAND2_X1 U638 ( .A1(n451), .A2(n546), .ZN(n575) );
  NOR2_X1 U639 ( .A1(n575), .A2(n547), .ZN(n548) );
  XNOR2_X1 U640 ( .A(n548), .B(KEYINPUT103), .ZN(n550) );
  INV_X1 U641 ( .A(n678), .ZN(n549) );
  NAND2_X1 U642 ( .A1(n365), .A2(n623), .ZN(n551) );
  NOR2_X1 U643 ( .A1(n557), .A2(n551), .ZN(n553) );
  XNOR2_X1 U644 ( .A(KEYINPUT105), .B(KEYINPUT43), .ZN(n552) );
  XNOR2_X1 U645 ( .A(n553), .B(n552), .ZN(n554) );
  NAND2_X1 U646 ( .A1(n568), .A2(n554), .ZN(n555) );
  XOR2_X1 U647 ( .A(KEYINPUT106), .B(n555), .Z(n724) );
  NOR2_X1 U648 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U649 ( .A(n558), .B(KEYINPUT36), .ZN(n560) );
  NAND2_X1 U650 ( .A1(n560), .A2(n559), .ZN(n561) );
  INV_X1 U651 ( .A(n720), .ZN(n599) );
  NAND2_X1 U652 ( .A1(n562), .A2(n623), .ZN(n563) );
  INV_X1 U653 ( .A(n564), .ZN(n565) );
  AND2_X1 U654 ( .A1(n566), .A2(n565), .ZN(n567) );
  INV_X1 U655 ( .A(KEYINPUT39), .ZN(n569) );
  AND2_X1 U656 ( .A1(n678), .A2(n602), .ZN(n570) );
  XNOR2_X1 U657 ( .A(n570), .B(KEYINPUT40), .ZN(n725) );
  INV_X1 U658 ( .A(n571), .ZN(n624) );
  NAND2_X1 U659 ( .A1(n624), .A2(n623), .ZN(n627) );
  INV_X1 U660 ( .A(n572), .ZN(n626) );
  NOR2_X1 U661 ( .A1(n627), .A2(n626), .ZN(n574) );
  XNOR2_X1 U662 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n573) );
  NOR2_X1 U663 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U664 ( .A(n577), .B(KEYINPUT28), .ZN(n580) );
  XNOR2_X1 U665 ( .A(n578), .B(KEYINPUT107), .ZN(n579) );
  NAND2_X1 U666 ( .A1(n580), .A2(n579), .ZN(n586) );
  NOR2_X1 U667 ( .A1(n655), .A2(n586), .ZN(n581) );
  XNOR2_X1 U668 ( .A(KEYINPUT42), .B(n581), .ZN(n726) );
  NOR2_X1 U669 ( .A1(n628), .A2(KEYINPUT47), .ZN(n584) );
  XNOR2_X1 U670 ( .A(n584), .B(KEYINPUT72), .ZN(n587) );
  NOR2_X1 U671 ( .A1(n586), .A2(n585), .ZN(n674) );
  NAND2_X1 U672 ( .A1(n587), .A2(n674), .ZN(n588) );
  XNOR2_X1 U673 ( .A(n588), .B(KEYINPUT71), .ZN(n596) );
  NAND2_X1 U674 ( .A1(n382), .A2(n674), .ZN(n589) );
  NAND2_X1 U675 ( .A1(n589), .A2(KEYINPUT47), .ZN(n594) );
  NOR2_X1 U676 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U677 ( .A1(n593), .A2(n592), .ZN(n672) );
  NAND2_X1 U678 ( .A1(n594), .A2(n672), .ZN(n595) );
  NOR2_X1 U679 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U680 ( .A1(n599), .A2(n429), .ZN(n600) );
  XNOR2_X1 U681 ( .A(n600), .B(KEYINPUT48), .ZN(n601) );
  NAND2_X1 U682 ( .A1(n602), .A2(n680), .ZN(n682) );
  NAND2_X1 U683 ( .A1(n603), .A2(n682), .ZN(n609) );
  INV_X1 U684 ( .A(n609), .ZN(n713) );
  NAND2_X1 U685 ( .A1(n604), .A2(n713), .ZN(n608) );
  XNOR2_X1 U686 ( .A(KEYINPUT79), .B(n605), .ZN(n606) );
  NAND2_X1 U687 ( .A1(n606), .A2(KEYINPUT2), .ZN(n607) );
  NAND2_X1 U688 ( .A1(n620), .A2(KEYINPUT2), .ZN(n610) );
  XNOR2_X1 U689 ( .A(KEYINPUT55), .B(KEYINPUT82), .ZN(n614) );
  XNOR2_X1 U690 ( .A(n612), .B(KEYINPUT54), .ZN(n613) );
  NAND2_X1 U691 ( .A1(G478), .A2(n690), .ZN(n616) );
  INV_X1 U692 ( .A(KEYINPUT2), .ZN(n622) );
  NOR2_X1 U693 ( .A1(n620), .A2(KEYINPUT77), .ZN(n621) );
  XNOR2_X1 U694 ( .A(n622), .B(n621), .ZN(n659) );
  NOR2_X1 U695 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U696 ( .A1(n626), .A2(n625), .ZN(n630) );
  NOR2_X1 U697 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U698 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U699 ( .A1(n631), .A2(n654), .ZN(n649) );
  NAND2_X1 U700 ( .A1(n365), .A2(n632), .ZN(n634) );
  XNOR2_X1 U701 ( .A(KEYINPUT50), .B(n634), .ZN(n641) );
  NAND2_X1 U702 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U703 ( .A(KEYINPUT49), .B(n637), .ZN(n638) );
  NOR2_X1 U704 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U705 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U706 ( .A(n642), .B(KEYINPUT114), .ZN(n644) );
  NAND2_X1 U707 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U708 ( .A(KEYINPUT51), .B(n645), .ZN(n646) );
  NOR2_X1 U709 ( .A1(n655), .A2(n646), .ZN(n647) );
  XOR2_X1 U710 ( .A(KEYINPUT115), .B(n647), .Z(n648) );
  NOR2_X1 U711 ( .A1(n649), .A2(n648), .ZN(n650) );
  XOR2_X1 U712 ( .A(KEYINPUT116), .B(n650), .Z(n651) );
  XOR2_X1 U713 ( .A(KEYINPUT52), .B(n651), .Z(n652) );
  NOR2_X1 U714 ( .A1(n653), .A2(n652), .ZN(n657) );
  NOR2_X1 U715 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U716 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U717 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U718 ( .A(n662), .B(G101), .Z(G3) );
  NAND2_X1 U719 ( .A1(n664), .A2(n678), .ZN(n663) );
  XNOR2_X1 U720 ( .A(n663), .B(G104), .ZN(G6) );
  XOR2_X1 U721 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n666) );
  NAND2_X1 U722 ( .A1(n664), .A2(n680), .ZN(n665) );
  XNOR2_X1 U723 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U724 ( .A(G107), .B(n667), .ZN(G9) );
  XNOR2_X1 U725 ( .A(G110), .B(n668), .ZN(G12) );
  XOR2_X1 U726 ( .A(KEYINPUT29), .B(KEYINPUT111), .Z(n670) );
  NAND2_X1 U727 ( .A1(n674), .A2(n680), .ZN(n669) );
  XNOR2_X1 U728 ( .A(n670), .B(n669), .ZN(n671) );
  XOR2_X1 U729 ( .A(G128), .B(n671), .Z(G30) );
  XNOR2_X1 U730 ( .A(G143), .B(KEYINPUT112), .ZN(n673) );
  XNOR2_X1 U731 ( .A(n673), .B(n672), .ZN(G45) );
  XOR2_X1 U732 ( .A(G146), .B(KEYINPUT113), .Z(n676) );
  NAND2_X1 U733 ( .A1(n674), .A2(n678), .ZN(n675) );
  XNOR2_X1 U734 ( .A(n676), .B(n675), .ZN(G48) );
  NAND2_X1 U735 ( .A1(n677), .A2(n678), .ZN(n679) );
  XNOR2_X1 U736 ( .A(n679), .B(G113), .ZN(G15) );
  NAND2_X1 U737 ( .A1(n680), .A2(n677), .ZN(n681) );
  XNOR2_X1 U738 ( .A(n681), .B(G116), .ZN(G18) );
  XNOR2_X1 U739 ( .A(G134), .B(n682), .ZN(G36) );
  XOR2_X1 U740 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n683) );
  NOR2_X1 U741 ( .A1(n694), .A2(n685), .ZN(G54) );
  XOR2_X1 U742 ( .A(KEYINPUT59), .B(KEYINPUT83), .Z(n686) );
  XNOR2_X1 U743 ( .A(n689), .B(KEYINPUT120), .ZN(n692) );
  NAND2_X1 U744 ( .A1(G217), .A2(n690), .ZN(n691) );
  XNOR2_X1 U745 ( .A(n692), .B(n691), .ZN(n693) );
  NOR2_X1 U746 ( .A1(n694), .A2(n693), .ZN(G66) );
  XNOR2_X1 U747 ( .A(n695), .B(KEYINPUT121), .ZN(n697) );
  NAND2_X1 U748 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U749 ( .A(n698), .B(KEYINPUT122), .ZN(n705) );
  NAND2_X1 U750 ( .A1(G953), .A2(G224), .ZN(n699) );
  XNOR2_X1 U751 ( .A(KEYINPUT61), .B(n699), .ZN(n700) );
  NAND2_X1 U752 ( .A1(n700), .A2(G898), .ZN(n703) );
  OR2_X1 U753 ( .A1(n701), .A2(G953), .ZN(n702) );
  NAND2_X1 U754 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U755 ( .A(n705), .B(n704), .Z(G69) );
  XNOR2_X1 U756 ( .A(G227), .B(KEYINPUT123), .ZN(n708) );
  XOR2_X1 U757 ( .A(n707), .B(n706), .Z(n714) );
  XNOR2_X1 U758 ( .A(n708), .B(n714), .ZN(n709) );
  NAND2_X1 U759 ( .A1(G900), .A2(n709), .ZN(n710) );
  XOR2_X1 U760 ( .A(KEYINPUT124), .B(n710), .Z(n711) );
  NOR2_X1 U761 ( .A1(n715), .A2(n711), .ZN(n712) );
  XNOR2_X1 U762 ( .A(KEYINPUT125), .B(n712), .ZN(n718) );
  XNOR2_X1 U763 ( .A(n714), .B(n713), .ZN(n716) );
  NAND2_X1 U764 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U765 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U766 ( .A(n719), .B(KEYINPUT126), .ZN(G72) );
  XNOR2_X1 U767 ( .A(n720), .B(G125), .ZN(n721) );
  XNOR2_X1 U768 ( .A(n721), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U769 ( .A(n722), .B(G122), .ZN(G24) );
  XNOR2_X1 U770 ( .A(n723), .B(G119), .ZN(G21) );
  XOR2_X1 U771 ( .A(G140), .B(n724), .Z(G42) );
  XOR2_X1 U772 ( .A(n725), .B(G131), .Z(G33) );
  XNOR2_X1 U773 ( .A(G137), .B(KEYINPUT127), .ZN(n727) );
  XNOR2_X1 U774 ( .A(n727), .B(n726), .ZN(G39) );
endmodule

