//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 0 1 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n537, new_n538, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n564, new_n565, new_n566, new_n568, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT65), .B(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT66), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI211_X1 g042(.A(G137), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n467), .A2(new_n470), .ZN(G160));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(G2105), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n479));
  INV_X1    g054(.A(G124), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n474), .A2(new_n475), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n477), .B(new_n479), .C1(new_n480), .C2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  OAI211_X1 g059(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n485));
  OR2_X1    g060(.A1(G102), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G114), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n486), .A2(new_n488), .A3(G2104), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g065(.A(G138), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n481), .A2(new_n493), .A3(G138), .A4(new_n462), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n490), .B1(new_n492), .B2(new_n494), .ZN(G164));
  INV_X1    g070(.A(KEYINPUT5), .ZN(new_n496));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n500), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT6), .B(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G50), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n505), .A2(new_n506), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n503), .A2(new_n513), .ZN(G166));
  INV_X1    g089(.A(G51), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT67), .B(G89), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n505), .A2(new_n515), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n500), .A2(G63), .A3(G651), .ZN(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n517), .A2(new_n521), .ZN(G168));
  AOI22_X1  g097(.A1(new_n500), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n523), .A2(new_n502), .ZN(new_n524));
  INV_X1    g099(.A(G52), .ZN(new_n525));
  INV_X1    g100(.A(G90), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n505), .A2(new_n525), .B1(new_n511), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n524), .A2(new_n527), .ZN(G171));
  AOI22_X1  g103(.A1(new_n500), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n502), .ZN(new_n530));
  INV_X1    g105(.A(G43), .ZN(new_n531));
  INV_X1    g106(.A(G81), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n505), .A2(new_n531), .B1(new_n511), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G860), .ZN(G153));
  NAND4_X1  g110(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g111(.A1(G1), .A2(G3), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT8), .ZN(new_n538));
  NAND4_X1  g113(.A1(G319), .A2(G483), .A3(G661), .A4(new_n538), .ZN(G188));
  NOR2_X1   g114(.A1(new_n509), .A2(new_n510), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n497), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT9), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n541), .A2(new_n542), .A3(G53), .ZN(new_n543));
  INV_X1    g118(.A(G53), .ZN(new_n544));
  OAI21_X1  g119(.A(KEYINPUT9), .B1(new_n505), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT68), .ZN(new_n547));
  INV_X1    g122(.A(G65), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n500), .A2(KEYINPUT70), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n508), .A2(new_n507), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT70), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n548), .B1(new_n549), .B2(new_n552), .ZN(new_n553));
  AND2_X1   g128(.A1(G78), .A2(G543), .ZN(new_n554));
  OAI21_X1  g129(.A(G651), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n511), .A2(KEYINPUT69), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT69), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n500), .A2(new_n504), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n556), .A2(G91), .A3(new_n558), .ZN(new_n559));
  AND2_X1   g134(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n547), .A2(new_n560), .ZN(G299));
  INV_X1    g136(.A(G171), .ZN(G301));
  INV_X1    g137(.A(G168), .ZN(G286));
  INV_X1    g138(.A(KEYINPUT71), .ZN(new_n564));
  NAND2_X1  g139(.A1(G166), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT71), .B1(new_n503), .B2(new_n513), .ZN(new_n566));
  AND2_X1   g141(.A1(new_n565), .A2(new_n566), .ZN(G303));
  INV_X1    g142(.A(G74), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n502), .B1(new_n550), .B2(new_n568), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n569), .B1(G49), .B2(new_n541), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n556), .A2(G87), .A3(new_n558), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(G288));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G61), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n498), .B2(new_n499), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n573), .B1(new_n575), .B2(KEYINPUT72), .ZN(new_n576));
  OAI211_X1 g151(.A(KEYINPUT72), .B(G61), .C1(new_n508), .C2(new_n507), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n556), .A2(G86), .A3(new_n558), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n504), .A2(G48), .A3(G543), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(G305));
  AOI22_X1  g157(.A1(new_n500), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n502), .ZN(new_n584));
  INV_X1    g159(.A(G47), .ZN(new_n585));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n505), .A2(new_n585), .B1(new_n511), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G290));
  INV_X1    g164(.A(G868), .ZN(new_n590));
  NOR2_X1   g165(.A1(G301), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  AND2_X1   g167(.A1(new_n549), .A2(new_n552), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  OAI211_X1 g169(.A(KEYINPUT73), .B(new_n592), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT73), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n594), .B1(new_n549), .B2(new_n552), .ZN(new_n597));
  INV_X1    g172(.A(new_n592), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n595), .A2(new_n599), .A3(G651), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n556), .A2(G92), .A3(new_n558), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n601), .B(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n541), .A2(G54), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n600), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(KEYINPUT74), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n601), .A2(new_n602), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n601), .A2(new_n602), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n607), .A2(new_n608), .B1(G54), .B2(new_n541), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT74), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n609), .A2(new_n610), .A3(new_n600), .ZN(new_n611));
  AND2_X1   g186(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n591), .B1(new_n612), .B2(new_n590), .ZN(G284));
  AOI21_X1  g188(.A(new_n591), .B1(new_n612), .B2(new_n590), .ZN(G321));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  INV_X1    g190(.A(G299), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G297));
  OAI21_X1  g192(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n612), .B1(new_n619), .B2(G860), .ZN(G148));
  OAI21_X1  g195(.A(new_n590), .B1(new_n530), .B2(new_n533), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n606), .A2(new_n611), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n622), .A2(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n621), .B1(new_n623), .B2(new_n590), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g200(.A(KEYINPUT75), .B(KEYINPUT12), .ZN(new_n626));
  NOR3_X1   g201(.A1(new_n472), .A2(new_n473), .A3(G2105), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT13), .Z(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G2100), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT76), .Z(new_n631));
  NAND2_X1  g206(.A1(new_n476), .A2(G135), .ZN(new_n632));
  OR2_X1    g207(.A1(G99), .A2(G2105), .ZN(new_n633));
  OAI211_X1 g208(.A(new_n633), .B(G2104), .C1(G111), .C2(new_n462), .ZN(new_n634));
  INV_X1    g209(.A(G123), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n632), .B(new_n634), .C1(new_n635), .C2(new_n482), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT77), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2096), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n631), .B(new_n638), .C1(G2100), .C2(new_n629), .ZN(G156));
  XOR2_X1   g214(.A(G2427), .B(G2430), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT79), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT78), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(KEYINPUT14), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT80), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n641), .A2(new_n644), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n647), .A2(new_n648), .A3(new_n651), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT81), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G1341), .ZN(new_n658));
  INV_X1    g233(.A(G1348), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n655), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(G14), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n655), .A2(new_n661), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(G401));
  XOR2_X1   g241(.A(KEYINPUT82), .B(KEYINPUT18), .Z(new_n667));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(KEYINPUT17), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n668), .A2(new_n669), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n667), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2072), .B(G2078), .Z(new_n674));
  INV_X1    g249(.A(new_n667), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n674), .B1(new_n670), .B2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n673), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2096), .B(G2100), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G227));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT19), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G1956), .B(G2474), .Z(new_n683));
  XOR2_X1   g258(.A(G1961), .B(G1966), .Z(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT20), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n683), .A2(new_n684), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  MUX2_X1   g265(.A(new_n690), .B(new_n689), .S(new_n682), .Z(new_n691));
  NOR2_X1   g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1981), .B(G1986), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT83), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n694), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1991), .B(G1996), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(G229));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G23), .ZN(new_n701));
  INV_X1    g276(.A(G288), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(new_n700), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT33), .B(G1976), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT84), .B(G16), .Z(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n707), .A2(G22), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G166), .B2(new_n707), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(G1971), .Z(new_n710));
  AND2_X1   g285(.A1(new_n700), .A2(G6), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G305), .B2(G16), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT32), .B(G1981), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n712), .A2(new_n714), .ZN(new_n716));
  NAND4_X1  g291(.A1(new_n705), .A2(new_n710), .A3(new_n715), .A4(new_n716), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n717), .A2(KEYINPUT34), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n707), .A2(G24), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n588), .B2(new_n707), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(G1986), .ZN(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G25), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n476), .A2(G131), .ZN(new_n724));
  OR2_X1    g299(.A1(G95), .A2(G2105), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n725), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n726));
  INV_X1    g301(.A(G119), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n724), .B(new_n726), .C1(new_n727), .C2(new_n482), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n723), .B1(new_n729), .B2(new_n722), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT35), .B(G1991), .Z(new_n731));
  XOR2_X1   g306(.A(new_n730), .B(new_n731), .Z(new_n732));
  INV_X1    g307(.A(KEYINPUT85), .ZN(new_n733));
  AOI211_X1 g308(.A(new_n721), .B(new_n732), .C1(new_n733), .C2(KEYINPUT36), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n718), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(KEYINPUT34), .B2(new_n717), .ZN(new_n736));
  OR3_X1    g311(.A1(new_n736), .A2(new_n733), .A3(KEYINPUT36), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n733), .B2(KEYINPUT36), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n707), .A2(G19), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n534), .B2(new_n707), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G1341), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n722), .A2(G32), .ZN(new_n742));
  NAND3_X1  g317(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT26), .Z(new_n744));
  NAND2_X1  g319(.A1(new_n476), .A2(G141), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n481), .A2(G129), .A3(G2105), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n744), .A2(new_n745), .A3(new_n746), .A4(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n742), .B1(new_n749), .B2(new_n722), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT27), .B(G1996), .Z(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT87), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n750), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n722), .A2(G33), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT25), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n476), .A2(G139), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n481), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n759), .A2(new_n462), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n754), .B1(new_n761), .B2(new_n722), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G2072), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n636), .A2(new_n722), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT30), .B(G28), .ZN(new_n765));
  OR2_X1    g340(.A1(KEYINPUT31), .A2(G11), .ZN(new_n766));
  NAND2_X1  g341(.A1(KEYINPUT31), .A2(G11), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n765), .A2(new_n722), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n753), .A2(new_n763), .A3(new_n764), .A4(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(G2078), .ZN(new_n770));
  NOR2_X1   g345(.A1(G164), .A2(new_n722), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G27), .B2(new_n722), .ZN(new_n772));
  AOI211_X1 g347(.A(new_n741), .B(new_n769), .C1(new_n770), .C2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n700), .A2(G5), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G171), .B2(new_n700), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n775), .A2(G1961), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT90), .Z(new_n777));
  NOR2_X1   g352(.A1(new_n772), .A2(new_n770), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n722), .A2(G26), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT28), .Z(new_n780));
  NAND2_X1  g355(.A1(new_n476), .A2(G140), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n481), .A2(G128), .A3(G2105), .ZN(new_n782));
  OR2_X1    g357(.A1(G104), .A2(G2105), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n783), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n781), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n780), .B1(new_n785), .B2(G29), .ZN(new_n786));
  INV_X1    g361(.A(G2067), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NOR3_X1   g363(.A1(new_n777), .A2(new_n778), .A3(new_n788), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT86), .B(KEYINPUT24), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G34), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n791), .A2(G29), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G29), .B2(G160), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n793), .A2(G2084), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT91), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n793), .A2(G2084), .ZN(new_n796));
  OAI221_X1 g371(.A(new_n796), .B1(G1961), .B2(new_n775), .C1(G2072), .C2(new_n762), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n773), .A2(new_n789), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n700), .A2(G21), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G168), .B2(new_n700), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT88), .ZN(new_n802));
  INV_X1    g377(.A(G1966), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT89), .Z(new_n805));
  NAND2_X1  g380(.A1(new_n706), .A2(G20), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT23), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n616), .B2(new_n700), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G1956), .ZN(new_n809));
  NOR2_X1   g384(.A1(G29), .A2(G35), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G162), .B2(G29), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT92), .B(KEYINPUT29), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n813), .A2(G2090), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(G2090), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n814), .B(new_n815), .C1(new_n803), .C2(new_n802), .ZN(new_n816));
  NOR4_X1   g391(.A1(new_n799), .A2(new_n805), .A3(new_n809), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n700), .A2(G4), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(new_n612), .B2(new_n700), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(new_n659), .ZN(new_n820));
  AND4_X1   g395(.A1(new_n737), .A2(new_n738), .A3(new_n817), .A4(new_n820), .ZN(G311));
  NAND4_X1  g396(.A1(new_n737), .A2(new_n738), .A3(new_n817), .A4(new_n820), .ZN(G150));
  INV_X1    g397(.A(G860), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n500), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n824), .A2(new_n502), .ZN(new_n825));
  INV_X1    g400(.A(G55), .ZN(new_n826));
  INV_X1    g401(.A(G93), .ZN(new_n827));
  OAI22_X1  g402(.A1(new_n505), .A2(new_n826), .B1(new_n511), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n534), .A2(new_n829), .ZN(new_n830));
  OAI22_X1  g405(.A1(new_n530), .A2(new_n533), .B1(new_n825), .B2(new_n828), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n606), .A2(G559), .A3(new_n611), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(KEYINPUT38), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n833), .A2(KEYINPUT38), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n832), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT38), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n612), .A2(new_n838), .A3(G559), .ZN(new_n839));
  INV_X1    g414(.A(new_n832), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n839), .A2(new_n834), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT39), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n823), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NOR3_X1   g419(.A1(new_n835), .A2(new_n832), .A3(new_n836), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n840), .B1(new_n839), .B2(new_n834), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n843), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT93), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n842), .A2(KEYINPUT93), .A3(new_n843), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n844), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n829), .A2(new_n823), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT94), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT37), .Z(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(KEYINPUT95), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT95), .ZN(new_n857));
  AOI21_X1  g432(.A(KEYINPUT93), .B1(new_n842), .B2(new_n843), .ZN(new_n858));
  AOI211_X1 g433(.A(new_n848), .B(KEYINPUT39), .C1(new_n837), .C2(new_n841), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n857), .B(new_n854), .C1(new_n860), .C2(new_n844), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n856), .A2(new_n861), .ZN(G145));
  XNOR2_X1  g437(.A(G160), .B(KEYINPUT96), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(G162), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n636), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n761), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT97), .ZN(new_n868));
  NAND2_X1  g443(.A1(G126), .A2(G2105), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n869), .B1(new_n474), .B2(new_n475), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n462), .A2(G114), .ZN(new_n871));
  OAI21_X1  g446(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n868), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n485), .A2(KEYINPUT97), .A3(new_n489), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n493), .B1(new_n476), .B2(G138), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n877));
  OAI211_X1 g452(.A(new_n874), .B(new_n875), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT98), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n785), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n781), .A2(new_n782), .A3(KEYINPUT98), .A4(new_n784), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n880), .A2(new_n748), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n748), .B1(new_n880), .B2(new_n881), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n878), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n880), .A2(new_n881), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n749), .ZN(new_n886));
  INV_X1    g461(.A(new_n878), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n880), .A2(new_n748), .A3(new_n881), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT100), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n884), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n890), .B1(new_n884), .B2(new_n889), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n867), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT101), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI211_X1 g470(.A(KEYINPUT101), .B(new_n867), .C1(new_n891), .C2(new_n892), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n884), .A2(new_n889), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n867), .B1(new_n897), .B2(KEYINPUT99), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT99), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n884), .A2(new_n889), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n902));
  INV_X1    g477(.A(G118), .ZN(new_n903));
  AOI22_X1  g478(.A1(new_n902), .A2(KEYINPUT102), .B1(new_n903), .B2(G2105), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n904), .B1(KEYINPUT102), .B2(new_n902), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n476), .A2(G142), .ZN(new_n906));
  INV_X1    g481(.A(G130), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n905), .B(new_n906), .C1(new_n907), .C2(new_n482), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n729), .B(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(new_n628), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n895), .A2(new_n896), .A3(new_n901), .A4(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT103), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI22_X1  g488(.A1(new_n893), .A2(new_n894), .B1(new_n900), .B2(new_n898), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n910), .B1(new_n914), .B2(new_n896), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n866), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(G37), .ZN(new_n917));
  INV_X1    g492(.A(new_n910), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n897), .A2(KEYINPUT100), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n884), .A2(new_n889), .A3(new_n890), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n761), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n901), .B1(new_n921), .B2(KEYINPUT101), .ZN(new_n922));
  INV_X1    g497(.A(new_n896), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n918), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n924), .A2(new_n912), .A3(new_n865), .A4(new_n911), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n916), .A2(new_n917), .A3(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g502(.A1(new_n623), .A2(new_n832), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n840), .B1(new_n622), .B2(G559), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(G299), .A2(new_n605), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n609), .A2(new_n547), .A3(new_n560), .A4(new_n600), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT41), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n931), .A2(KEYINPUT41), .A3(new_n932), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n930), .A2(new_n937), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n928), .A2(new_n933), .A3(new_n929), .ZN(new_n939));
  NOR2_X1   g514(.A1(G305), .A2(new_n588), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(G288), .A2(G166), .ZN(new_n942));
  OR2_X1    g517(.A1(G288), .A2(G166), .ZN(new_n943));
  NAND2_X1  g518(.A1(G305), .A2(new_n588), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n941), .A2(new_n942), .A3(new_n943), .A4(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  AOI22_X1  g521(.A1(new_n941), .A2(new_n944), .B1(new_n943), .B2(new_n942), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n946), .A2(KEYINPUT42), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n949), .B1(new_n946), .B2(new_n947), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n943), .A2(new_n942), .ZN(new_n951));
  INV_X1    g526(.A(new_n944), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n951), .B1(new_n952), .B2(new_n940), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n953), .A2(new_n945), .A3(KEYINPUT104), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n950), .A2(new_n954), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n955), .A2(KEYINPUT42), .ZN(new_n956));
  OAI22_X1  g531(.A1(new_n938), .A2(new_n939), .B1(new_n948), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n939), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n948), .B1(new_n955), .B2(KEYINPUT42), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n958), .B(new_n959), .C1(new_n930), .C2(new_n937), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(G868), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n962), .B1(G868), .B2(new_n829), .ZN(G295));
  OAI21_X1  g538(.A(new_n962), .B1(G868), .B2(new_n829), .ZN(G331));
  NAND2_X1  g539(.A1(G171), .A2(G168), .ZN(new_n965));
  OAI22_X1  g540(.A1(new_n524), .A2(new_n527), .B1(new_n517), .B2(new_n521), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OR2_X1    g542(.A1(new_n832), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n832), .A2(new_n967), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n969), .A2(KEYINPUT106), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT106), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n971), .B1(new_n832), .B2(new_n967), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n968), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n935), .A2(new_n973), .A3(new_n936), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n931), .A2(new_n968), .A3(new_n932), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n969), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n955), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n955), .A2(new_n974), .A3(new_n976), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n979), .A2(new_n917), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n968), .A2(new_n969), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n935), .A2(new_n936), .A3(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n975), .B1(new_n972), .B2(new_n970), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n917), .B(new_n980), .C1(new_n986), .C2(new_n955), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n982), .B1(KEYINPUT43), .B2(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT44), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n991), .B1(new_n987), .B2(KEYINPUT43), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT43), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n979), .A2(new_n993), .A3(new_n917), .A4(new_n980), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT107), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n980), .A2(new_n917), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n955), .B1(new_n984), .B2(new_n985), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT43), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AND4_X1   g573(.A1(KEYINPUT107), .A2(new_n998), .A3(KEYINPUT44), .A4(new_n994), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n990), .B1(new_n995), .B2(new_n999), .ZN(G397));
  INV_X1    g575(.A(G1384), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT45), .B1(new_n878), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G40), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n467), .A2(new_n470), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n785), .B(G2067), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n1008), .B(KEYINPUT108), .ZN(new_n1009));
  INV_X1    g584(.A(G1996), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n748), .B(new_n1010), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n729), .A2(new_n731), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n729), .A2(new_n731), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  XOR2_X1   g590(.A(new_n588), .B(G1986), .Z(new_n1016));
  OAI21_X1  g591(.A(new_n1007), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT50), .B1(new_n878), .B2(new_n1001), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n1019));
  NOR3_X1   g594(.A1(G164), .A2(new_n1019), .A3(G1384), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1005), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT119), .ZN(new_n1022));
  INV_X1    g597(.A(G1961), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT119), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1024), .B(new_n1005), .C1(new_n1018), .C2(new_n1020), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1022), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT45), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1027), .A2(G1384), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1005), .B1(G164), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1002), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1032), .A2(G2078), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n878), .A2(new_n1028), .ZN(new_n1035));
  NOR2_X1   g610(.A1(G164), .A2(G1384), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1035), .B(new_n1005), .C1(new_n1036), .C2(KEYINPUT45), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1032), .B1(new_n1037), .B2(G2078), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1026), .A2(G301), .A3(new_n1034), .A4(new_n1038), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n1039), .A2(KEYINPUT54), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1003), .A2(new_n1005), .A3(new_n1035), .A4(new_n1033), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1026), .A2(new_n1038), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT125), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1042), .A2(new_n1043), .A3(G171), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1043), .B1(new_n1042), .B2(G171), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1040), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1026), .A2(new_n1038), .A3(new_n1034), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n1048), .A2(G171), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1042), .A2(G171), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1047), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1006), .A2(G2084), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1052), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n803), .B1(new_n1002), .B2(new_n1030), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(G286), .A2(KEYINPUT122), .A3(G8), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT122), .ZN(new_n1057));
  INV_X1    g632(.A(G8), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1057), .B1(G168), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1055), .A2(new_n1060), .ZN(new_n1061));
  XOR2_X1   g636(.A(KEYINPUT123), .B(KEYINPUT51), .Z(new_n1062));
  NAND2_X1  g637(.A1(new_n1055), .A2(G8), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1056), .A2(new_n1059), .A3(KEYINPUT124), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT124), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1062), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1058), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n1068), .A2(KEYINPUT51), .A3(new_n1060), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1061), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  XOR2_X1   g645(.A(KEYINPUT109), .B(G1971), .Z(new_n1071));
  NAND2_X1  g646(.A1(new_n1037), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G2090), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1073), .B(new_n1005), .C1(new_n1018), .C2(new_n1020), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1058), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n565), .A2(G8), .A3(new_n566), .ZN(new_n1076));
  NAND2_X1  g651(.A1(KEYINPUT110), .A2(KEYINPUT55), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  XOR2_X1   g653(.A(KEYINPUT110), .B(KEYINPUT55), .Z(new_n1079));
  OAI21_X1  g654(.A(new_n1078), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1075), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1006), .B1(new_n1036), .B2(new_n1019), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n878), .A2(new_n1001), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT50), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1082), .A2(new_n1073), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1058), .B1(new_n1072), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1081), .B1(new_n1080), .B2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n878), .A2(new_n1005), .A3(new_n1001), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1088), .A2(G8), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n570), .A2(new_n571), .A3(G1976), .ZN(new_n1090));
  AND2_X1   g665(.A1(new_n1090), .A2(KEYINPUT111), .ZN(new_n1091));
  INV_X1    g666(.A(G1976), .ZN(new_n1092));
  NAND2_X1  g667(.A1(G288), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1089), .B(new_n1091), .C1(KEYINPUT52), .C2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1088), .A2(KEYINPUT111), .A3(G8), .A4(new_n1090), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT52), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1088), .A2(G8), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1096), .B(new_n1097), .C1(new_n1098), .C2(new_n1093), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1095), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT112), .ZN(new_n1101));
  OAI21_X1  g676(.A(G61), .B1(new_n508), .B2(new_n507), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT72), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1102), .A2(new_n1103), .B1(G73), .B2(G543), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n502), .B1(new_n1104), .B2(new_n577), .ZN(new_n1105));
  INV_X1    g680(.A(G86), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n581), .B1(new_n1106), .B2(new_n511), .ZN(new_n1107));
  OAI21_X1  g682(.A(G1981), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(G1981), .B1(new_n541), .B2(G48), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n579), .A2(new_n580), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT49), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1111), .A2(new_n1098), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1108), .A2(new_n1110), .A3(KEYINPUT49), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1101), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT49), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n579), .A2(new_n580), .A3(new_n1109), .ZN(new_n1116));
  INV_X1    g691(.A(G1981), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1107), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1117), .B1(new_n579), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1115), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1120));
  AND4_X1   g695(.A1(new_n1101), .A2(new_n1120), .A3(new_n1113), .A4(new_n1089), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1100), .B1(new_n1114), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT115), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT115), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1124), .B(new_n1100), .C1(new_n1114), .C2(new_n1121), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1087), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1046), .A2(new_n1051), .A3(new_n1070), .A4(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT57), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT118), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n560), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n555), .A2(new_n1129), .A3(new_n559), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n546), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1128), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n547), .A2(KEYINPUT57), .A3(new_n560), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  XOR2_X1   g710(.A(KEYINPUT56), .B(G2072), .Z(new_n1136));
  NOR2_X1   g711(.A1(new_n1037), .A2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g712(.A(KEYINPUT117), .B(G1956), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1139), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1135), .A2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1133), .B(new_n1134), .C1(new_n1137), .C2(new_n1140), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1142), .B1(new_n1144), .B2(KEYINPUT121), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT121), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1135), .A2(new_n1146), .A3(new_n1141), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1145), .A2(KEYINPUT61), .A3(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1022), .A2(new_n659), .A3(new_n1025), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1088), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n787), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n605), .B1(new_n1152), .B2(KEYINPUT60), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1153), .B1(KEYINPUT60), .B2(new_n1152), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT61), .ZN(new_n1156));
  XNOR2_X1  g731(.A(KEYINPUT58), .B(G1341), .ZN(new_n1157));
  OAI22_X1  g732(.A1(new_n1037), .A2(G1996), .B1(new_n1150), .B2(new_n1157), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1158), .A2(new_n534), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT59), .ZN(new_n1160));
  OR2_X1    g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1162));
  AOI22_X1  g737(.A1(new_n1155), .A2(new_n1156), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1152), .A2(KEYINPUT60), .A3(new_n605), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1148), .A2(new_n1154), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n605), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1142), .B1(new_n1144), .B2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT120), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1127), .B1(new_n1165), .B2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1122), .A2(new_n1081), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n702), .A2(new_n1092), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT113), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1172), .B1(new_n1114), .B2(new_n1121), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(new_n1110), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT114), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1098), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1173), .A2(KEYINPUT114), .A3(new_n1110), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1170), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1070), .A2(KEYINPUT62), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT62), .ZN(new_n1180));
  OAI211_X1 g755(.A(new_n1180), .B(new_n1061), .C1(new_n1067), .C2(new_n1069), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1126), .A2(new_n1179), .A3(new_n1049), .A4(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1068), .A2(G168), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(KEYINPUT63), .B1(new_n1126), .B2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1184), .A2(KEYINPUT63), .A3(new_n1081), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT116), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1075), .A2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1075), .A2(new_n1187), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n1189), .A2(new_n1080), .ZN(new_n1190));
  AOI211_X1 g765(.A(new_n1122), .B(new_n1186), .C1(new_n1188), .C2(new_n1190), .ZN(new_n1191));
  OAI211_X1 g766(.A(new_n1178), .B(new_n1182), .C1(new_n1185), .C2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1017), .B1(new_n1169), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1194));
  OR2_X1    g769(.A1(new_n1194), .A2(KEYINPUT46), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1194), .A2(KEYINPUT46), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1009), .A2(new_n749), .ZN(new_n1197));
  AOI22_X1  g772(.A1(new_n1195), .A2(new_n1196), .B1(new_n1007), .B2(new_n1197), .ZN(new_n1198));
  XOR2_X1   g773(.A(new_n1198), .B(KEYINPUT47), .Z(new_n1199));
  INV_X1    g774(.A(new_n1012), .ZN(new_n1200));
  OAI22_X1  g775(.A1(new_n1200), .A2(new_n1013), .B1(G2067), .B2(new_n785), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1201), .A2(new_n1007), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1015), .A2(new_n1007), .ZN(new_n1203));
  XOR2_X1   g778(.A(new_n1203), .B(KEYINPUT126), .Z(new_n1204));
  NOR4_X1   g779(.A1(new_n1003), .A2(G1986), .A3(G290), .A4(new_n1006), .ZN(new_n1205));
  XNOR2_X1  g780(.A(new_n1205), .B(KEYINPUT48), .ZN(new_n1206));
  OAI211_X1 g781(.A(new_n1199), .B(new_n1202), .C1(new_n1204), .C2(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1193), .A2(new_n1208), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g784(.A1(G227), .A2(new_n460), .ZN(new_n1211));
  NAND2_X1  g785(.A1(new_n665), .A2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g786(.A(G229), .B1(new_n1212), .B2(KEYINPUT127), .ZN(new_n1213));
  INV_X1    g787(.A(KEYINPUT127), .ZN(new_n1214));
  NAND3_X1  g788(.A1(new_n665), .A2(new_n1214), .A3(new_n1211), .ZN(new_n1215));
  NAND4_X1  g789(.A1(new_n988), .A2(new_n1213), .A3(new_n926), .A4(new_n1215), .ZN(G225));
  INV_X1    g790(.A(G225), .ZN(G308));
endmodule


