//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 0 0 0 0 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 1 1 1 1 0 1 0 1 1 0 0 0 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1260, new_n1261, new_n1262, new_n1263;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G250), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G257), .ZN(new_n210));
  INV_X1    g0010(.A(G264), .ZN(new_n211));
  AOI211_X1 g0011(.A(new_n206), .B(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(new_n212), .A2(KEYINPUT0), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n218), .B1(KEYINPUT0), .B2(new_n212), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT65), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G87), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n206), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  INV_X1    g0026(.A(G77), .ZN(new_n227));
  INV_X1    g0027(.A(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G107), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n226), .B1(new_n227), .B2(new_n228), .C1(new_n229), .C2(new_n211), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n207), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT1), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n220), .A2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT67), .ZN(new_n246));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G58), .ZN(new_n248));
  XOR2_X1   g0048(.A(KEYINPUT66), .B(G50), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n246), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(KEYINPUT84), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT18), .ZN(new_n253));
  NOR2_X1   g0053(.A1(KEYINPUT8), .A2(G58), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT70), .B(G58), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n254), .B1(new_n255), .B2(KEYINPUT8), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G13), .A3(G20), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n213), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n262), .B1(new_n257), .B2(G20), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n260), .B1(new_n256), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n262), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT78), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT7), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT3), .B(G33), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n268), .B1(new_n269), .B2(G20), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT3), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G33), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT3), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n268), .A2(KEYINPUT76), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT76), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT7), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n275), .A2(new_n279), .A3(new_n214), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT77), .ZN(new_n281));
  AND3_X1   g0081(.A1(new_n270), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n275), .A2(new_n279), .A3(KEYINPUT77), .A4(new_n214), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G68), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n267), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  AND2_X1   g0085(.A1(new_n283), .A2(G68), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n270), .A2(new_n280), .A3(new_n281), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n286), .A2(KEYINPUT78), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G159), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT79), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n291), .B(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n202), .B1(new_n255), .B2(G68), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n293), .B1(new_n214), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT16), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n266), .B1(new_n289), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n272), .A2(KEYINPUT80), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(new_n274), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n272), .A2(KEYINPUT80), .ZN(new_n301));
  OAI211_X1 g0101(.A(KEYINPUT7), .B(new_n214), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n276), .B(new_n278), .C1(new_n269), .C2(G20), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n222), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n296), .B1(new_n304), .B2(new_n295), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n265), .B1(new_n298), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT81), .ZN(new_n307));
  NAND2_X1  g0107(.A1(G33), .A2(G41), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n308), .A2(G1), .A3(G13), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n307), .B1(new_n311), .B2(new_n235), .ZN(new_n312));
  INV_X1    g0112(.A(G41), .ZN(new_n313));
  INV_X1    g0113(.A(G45), .ZN(new_n314));
  AOI21_X1  g0114(.A(G1), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n315), .A2(new_n309), .A3(G274), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n309), .A2(new_n310), .A3(KEYINPUT81), .A4(G232), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n312), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT82), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n269), .A2(G226), .A3(G1698), .ZN(new_n320));
  NAND2_X1  g0120(.A1(G33), .A2(G87), .ZN(new_n321));
  INV_X1    g0121(.A(G1698), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT68), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT68), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G1698), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n272), .A2(new_n274), .A3(new_n323), .A4(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G223), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n320), .B(new_n321), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n309), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT82), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n312), .A2(new_n331), .A3(new_n316), .A4(new_n317), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n319), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(KEYINPUT83), .B1(new_n333), .B2(G179), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n318), .A2(KEYINPUT82), .B1(new_n328), .B2(new_n329), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT83), .ZN(new_n336));
  INV_X1    g0136(.A(G179), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n335), .A2(new_n336), .A3(new_n337), .A4(new_n332), .ZN(new_n338));
  INV_X1    g0138(.A(G169), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n333), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n334), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n252), .B(new_n253), .C1(new_n306), .C2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G190), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n333), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G200), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n345), .B1(new_n335), .B2(new_n332), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NOR3_X1   g0147(.A1(new_n282), .A2(new_n267), .A3(new_n284), .ZN(new_n348));
  AOI21_X1  g0148(.A(KEYINPUT78), .B1(new_n286), .B2(new_n287), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n297), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n350), .A2(new_n305), .A3(new_n262), .ZN(new_n351));
  INV_X1    g0151(.A(new_n265), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n347), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT17), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n306), .A2(KEYINPUT17), .A3(new_n347), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n342), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NOR3_X1   g0157(.A1(new_n306), .A2(KEYINPUT18), .A3(new_n341), .ZN(new_n358));
  AND3_X1   g0158(.A1(new_n334), .A2(new_n338), .A3(new_n340), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n351), .A2(new_n352), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n253), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT84), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n263), .A2(G50), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n256), .A2(new_n214), .A3(G33), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n290), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI221_X1 g0168(.A(new_n365), .B1(G50), .B2(new_n258), .C1(new_n368), .C2(new_n266), .ZN(new_n369));
  XNOR2_X1  g0169(.A(KEYINPUT68), .B(G1698), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n269), .A2(new_n370), .A3(G222), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n269), .A2(G1698), .ZN(new_n372));
  OAI221_X1 g0172(.A(new_n371), .B1(new_n227), .B2(new_n269), .C1(new_n327), .C2(new_n372), .ZN(new_n373));
  OR2_X1    g0173(.A1(new_n373), .A2(KEYINPUT69), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n309), .B1(new_n373), .B2(KEYINPUT69), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G226), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n316), .B1(new_n377), .B2(new_n311), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n369), .B1(new_n379), .B2(G169), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n380), .B1(new_n337), .B2(new_n379), .ZN(new_n381));
  XNOR2_X1  g0181(.A(new_n369), .B(KEYINPUT9), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n379), .A2(G190), .ZN(new_n383));
  OAI21_X1  g0183(.A(G200), .B1(new_n376), .B2(new_n378), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT10), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT10), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n382), .A2(new_n383), .A3(new_n387), .A4(new_n384), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n381), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G33), .A2(G97), .ZN(new_n390));
  OAI221_X1 g0190(.A(new_n390), .B1(new_n326), .B2(new_n377), .C1(new_n235), .C2(new_n372), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n316), .B1(new_n223), .B2(new_n311), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT72), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT72), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n316), .B(new_n394), .C1(new_n223), .C2(new_n311), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n391), .A2(new_n329), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT13), .ZN(new_n397));
  XNOR2_X1  g0197(.A(new_n396), .B(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT14), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(new_n399), .A3(G169), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n396), .A2(new_n397), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n391), .A2(new_n329), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n393), .A2(new_n395), .ZN(new_n403));
  AND3_X1   g0203(.A1(new_n402), .A2(new_n397), .A3(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(G169), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT14), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n401), .A2(KEYINPUT73), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT73), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n396), .B2(new_n397), .ZN(new_n409));
  INV_X1    g0209(.A(new_n404), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n407), .A2(G179), .A3(new_n409), .A4(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n400), .A2(new_n406), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n259), .A2(KEYINPUT12), .A3(new_n222), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT12), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(new_n258), .B2(G68), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n413), .B(new_n415), .C1(new_n264), .C2(new_n222), .ZN(new_n416));
  XOR2_X1   g0216(.A(new_n416), .B(KEYINPUT75), .Z(new_n417));
  NAND2_X1  g0217(.A1(new_n290), .A2(G50), .ZN(new_n418));
  XOR2_X1   g0218(.A(new_n418), .B(KEYINPUT74), .Z(new_n419));
  NAND2_X1  g0219(.A1(new_n214), .A2(G33), .ZN(new_n420));
  OAI22_X1  g0220(.A1(new_n420), .A2(new_n227), .B1(new_n214), .B2(G68), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n262), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT11), .ZN(new_n423));
  AND2_X1   g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n422), .A2(new_n423), .ZN(new_n425));
  NOR3_X1   g0225(.A1(new_n417), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n412), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n407), .A2(G190), .A3(new_n409), .A4(new_n410), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n398), .A2(G200), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(new_n430), .A3(new_n426), .ZN(new_n431));
  XOR2_X1   g0231(.A(KEYINPUT8), .B(G58), .Z(new_n432));
  AOI22_X1  g0232(.A1(new_n432), .A2(new_n290), .B1(G20), .B2(G77), .ZN(new_n433));
  XNOR2_X1  g0233(.A(KEYINPUT15), .B(G87), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n433), .B1(new_n420), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n262), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n263), .A2(G77), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n436), .B(new_n437), .C1(G77), .C2(new_n258), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n316), .B1(new_n228), .B2(new_n311), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n275), .A2(G107), .ZN(new_n441));
  OAI221_X1 g0241(.A(new_n441), .B1(new_n326), .B2(new_n235), .C1(new_n223), .C2(new_n372), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n440), .B1(new_n442), .B2(new_n329), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n439), .B1(new_n345), .B2(new_n443), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n443), .A2(G190), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n438), .B1(G169), .B2(new_n443), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n447), .A2(KEYINPUT71), .B1(new_n337), .B2(new_n443), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT71), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n438), .B(new_n449), .C1(G169), .C2(new_n443), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n446), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n428), .A2(new_n431), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n364), .A2(new_n389), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT5), .B(G41), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n314), .A2(G1), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n457), .A2(G257), .A3(new_n309), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n455), .A2(G274), .A3(new_n309), .A4(new_n456), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT4), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n461), .B1(new_n326), .B2(new_n228), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n269), .A2(new_n370), .A3(KEYINPUT4), .A4(G244), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n269), .A2(G250), .A3(G1698), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G283), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n462), .A2(new_n463), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n460), .B1(new_n466), .B2(new_n329), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(KEYINPUT87), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT87), .ZN(new_n469));
  AOI211_X1 g0269(.A(new_n469), .B(new_n460), .C1(new_n466), .C2(new_n329), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n339), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n302), .A2(new_n303), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G107), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n229), .A2(KEYINPUT6), .A3(G97), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT85), .ZN(new_n475));
  OR2_X1    g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n474), .A2(new_n475), .ZN(new_n477));
  XOR2_X1   g0277(.A(G97), .B(G107), .Z(new_n478));
  OAI211_X1 g0278(.A(new_n476), .B(new_n477), .C1(new_n478), .C2(KEYINPUT6), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n479), .A2(G20), .B1(G77), .B2(new_n290), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n473), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n262), .ZN(new_n482));
  INV_X1    g0282(.A(G97), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n259), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n257), .A2(G33), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n258), .A2(new_n485), .A3(new_n213), .A4(new_n261), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n484), .B1(new_n486), .B2(new_n483), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n482), .A2(KEYINPUT88), .A3(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT88), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n266), .B1(new_n473), .B2(new_n480), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n490), .B1(new_n491), .B2(new_n487), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n467), .A2(new_n337), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n471), .A2(new_n489), .A3(new_n492), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n466), .A2(new_n329), .ZN(new_n495));
  INV_X1    g0295(.A(new_n460), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT86), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n497), .A2(new_n498), .A3(G200), .ZN(new_n499));
  OAI21_X1  g0299(.A(KEYINPUT86), .B1(new_n467), .B2(new_n345), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n497), .A2(new_n469), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n467), .A2(KEYINPUT87), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n502), .A2(G190), .A3(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n491), .A2(new_n487), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n501), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n434), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n507), .A2(new_n258), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n269), .A2(new_n214), .A3(G68), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT19), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n214), .B1(new_n390), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n224), .A2(new_n483), .A3(new_n229), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n510), .B1(new_n420), .B2(new_n483), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n509), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n508), .B1(new_n515), .B2(new_n262), .ZN(new_n516));
  INV_X1    g0316(.A(new_n486), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n507), .ZN(new_n518));
  AND2_X1   g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n309), .A2(G274), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n456), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n309), .B(G250), .C1(G1), .C2(new_n314), .ZN(new_n522));
  INV_X1    g0322(.A(G116), .ZN(new_n523));
  OAI22_X1  g0323(.A1(new_n372), .A2(new_n228), .B1(new_n273), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT89), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n269), .A2(new_n370), .A3(new_n525), .A4(G238), .ZN(new_n526));
  OAI21_X1  g0326(.A(KEYINPUT89), .B1(new_n326), .B2(new_n223), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n521), .B(new_n522), .C1(new_n528), .C2(new_n309), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n519), .B1(new_n529), .B2(new_n339), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n521), .A2(new_n522), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n527), .A2(new_n526), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n273), .A2(new_n523), .ZN(new_n533));
  INV_X1    g0333(.A(new_n372), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n533), .B1(new_n534), .B2(G244), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n531), .B1(new_n536), .B2(new_n329), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n337), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n516), .B1(new_n224), .B2(new_n486), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n539), .B1(new_n537), .B2(G190), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n529), .A2(G200), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n530), .A2(new_n538), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT90), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n494), .A2(new_n506), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n494), .A2(new_n506), .A3(new_n542), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT90), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT94), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(new_n326), .B2(new_n206), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n269), .A2(new_n370), .A3(KEYINPUT94), .A4(G250), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n275), .A2(new_n210), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G1698), .ZN(new_n552));
  NAND2_X1  g0352(.A1(G33), .A2(G294), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n329), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n329), .B1(new_n456), .B2(new_n455), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(G264), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n555), .A2(new_n337), .A3(new_n459), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n269), .A2(G257), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n553), .B1(new_n559), .B2(new_n322), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n560), .B1(new_n548), .B2(new_n549), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n459), .B(new_n557), .C1(new_n561), .C2(new_n309), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n339), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n272), .A2(new_n274), .A3(new_n214), .A4(G87), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(KEYINPUT22), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT22), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n269), .A2(new_n566), .A3(new_n214), .A4(G87), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT24), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT23), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(new_n214), .B2(G107), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n229), .A2(KEYINPUT23), .A3(G20), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n571), .A2(new_n572), .B1(new_n533), .B2(new_n214), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n568), .A2(new_n569), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n569), .B1(new_n568), .B2(new_n573), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n262), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n259), .A2(KEYINPUT25), .A3(new_n229), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT25), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n258), .B2(G107), .ZN(new_n579));
  AOI22_X1  g0379(.A1(G107), .A2(new_n517), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n558), .A2(new_n563), .A3(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT95), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n563), .A2(new_n558), .A3(new_n581), .A4(KEYINPUT95), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n554), .A2(new_n329), .B1(G264), .B2(new_n556), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n586), .A2(G190), .A3(new_n459), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n562), .A2(G200), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n587), .A2(new_n576), .A3(new_n580), .A4(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n584), .A2(new_n585), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT21), .ZN(new_n591));
  INV_X1    g0391(.A(G303), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n592), .B1(new_n272), .B2(new_n274), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n593), .B1(new_n551), .B2(new_n370), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n534), .A2(G264), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n309), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n556), .A2(G270), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n459), .ZN(new_n598));
  OAI21_X1  g0398(.A(G169), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n465), .B(new_n214), .C1(G33), .C2(new_n483), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n523), .A2(G20), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n600), .A2(new_n262), .A3(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT20), .ZN(new_n603));
  XNOR2_X1  g0403(.A(new_n602), .B(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT91), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n517), .A2(new_n605), .A3(G116), .ZN(new_n606));
  OAI21_X1  g0406(.A(KEYINPUT91), .B1(new_n486), .B2(new_n523), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n259), .A2(new_n523), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n604), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n591), .B1(new_n599), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT93), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT93), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n613), .B(new_n591), .C1(new_n599), .C2(new_n610), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n370), .ZN(new_n616));
  OAI22_X1  g0416(.A1(new_n559), .A2(new_n616), .B1(new_n592), .B2(new_n269), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n372), .A2(new_n211), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n329), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n457), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n556), .A2(G270), .B1(new_n620), .B2(new_n520), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n619), .A2(G179), .A3(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(KEYINPUT92), .B1(new_n610), .B2(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n596), .A2(new_n598), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT92), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n604), .A2(new_n608), .A3(new_n609), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n624), .A2(new_n625), .A3(G179), .A4(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n599), .A2(new_n610), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n623), .A2(new_n627), .B1(new_n628), .B2(KEYINPUT21), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n624), .A2(G190), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n630), .B(new_n610), .C1(new_n345), .C2(new_n624), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n615), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n590), .A2(new_n632), .ZN(new_n633));
  AND4_X1   g0433(.A1(new_n454), .A2(new_n544), .A3(new_n546), .A4(new_n633), .ZN(G372));
  INV_X1    g0434(.A(new_n589), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n615), .A2(new_n629), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  AOI211_X1 g0437(.A(new_n635), .B(new_n545), .C1(new_n582), .C2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n542), .ZN(new_n639));
  OAI21_X1  g0439(.A(KEYINPUT26), .B1(new_n639), .B2(new_n494), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n530), .A2(new_n538), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n471), .A2(new_n493), .ZN(new_n642));
  INV_X1    g0442(.A(new_n505), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(new_n542), .A3(new_n643), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n640), .B(new_n641), .C1(KEYINPUT26), .C2(new_n644), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n638), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n454), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n647), .B(KEYINPUT96), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n359), .A2(new_n360), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(KEYINPUT18), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n359), .A2(new_n360), .A3(new_n253), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n448), .A2(new_n450), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n653), .A2(new_n431), .B1(new_n412), .B2(new_n427), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n355), .A2(new_n356), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n650), .B(new_n651), .C1(new_n654), .C2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n386), .A2(new_n388), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n381), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n648), .A2(new_n658), .ZN(G369));
  NAND3_X1  g0459(.A1(new_n257), .A2(new_n214), .A3(G13), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(G213), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(G343), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n610), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n636), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n632), .B2(new_n667), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G330), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n666), .B1(new_n576), .B2(new_n580), .ZN(new_n672));
  OAI22_X1  g0472(.A1(new_n590), .A2(new_n672), .B1(new_n582), .B2(new_n666), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n637), .A2(new_n665), .ZN(new_n676));
  INV_X1    g0476(.A(new_n590), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n582), .B2(new_n665), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n675), .A2(new_n679), .ZN(G399));
  NOR2_X1   g0480(.A1(new_n209), .A2(G41), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n512), .A2(G116), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G1), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n216), .B2(new_n682), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT28), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT29), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n644), .A2(KEYINPUT26), .ZN(new_n688));
  INV_X1    g0488(.A(new_n494), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT26), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(new_n690), .A3(new_n542), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n641), .B(KEYINPUT97), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n688), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT98), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n688), .A2(new_n691), .A3(KEYINPUT98), .A4(new_n692), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n545), .A2(new_n635), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n584), .A2(new_n585), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n697), .B1(new_n698), .B2(new_n636), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n695), .A2(new_n696), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n687), .B1(new_n700), .B2(new_n666), .ZN(new_n701));
  INV_X1    g0501(.A(G330), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n502), .A2(new_n503), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n586), .A2(G179), .A3(new_n537), .A4(new_n624), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n557), .B1(new_n561), .B2(new_n309), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n529), .A2(new_n707), .A3(new_n622), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n468), .A2(new_n470), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(new_n709), .A3(KEYINPUT30), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n624), .A2(new_n467), .A3(G179), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n711), .A2(new_n529), .A3(new_n562), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n706), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  AND3_X1   g0513(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n665), .ZN(new_n714));
  AOI21_X1  g0514(.A(KEYINPUT31), .B1(new_n713), .B2(new_n665), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n633), .A2(new_n546), .A3(new_n544), .A4(new_n666), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n702), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n687), .B(new_n666), .C1(new_n638), .C2(new_n645), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n701), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n686), .B1(new_n721), .B2(G1), .ZN(G364));
  INV_X1    g0522(.A(G13), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G20), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n257), .B1(new_n724), .B2(G45), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  OR3_X1    g0526(.A1(new_n681), .A2(new_n726), .A3(KEYINPUT99), .ZN(new_n727));
  OAI21_X1  g0527(.A(KEYINPUT99), .B1(new_n681), .B2(new_n726), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n671), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n731), .B1(G330), .B2(new_n669), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G13), .A2(G33), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(G20), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n213), .B1(G20), .B2(new_n339), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n250), .A2(G45), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n275), .A2(new_n208), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n740), .B1(new_n314), .B2(new_n217), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT102), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n269), .A2(new_n208), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n743), .B(KEYINPUT100), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  XOR2_X1   g0545(.A(G355), .B(KEYINPUT101), .Z(new_n746));
  OAI22_X1  g0546(.A1(new_n745), .A2(new_n746), .B1(G116), .B2(new_n208), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n739), .A2(new_n741), .B1(new_n742), .B2(new_n747), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n747), .A2(new_n742), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n738), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n214), .A2(G179), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G190), .A2(G200), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g0553(.A(KEYINPUT103), .B(G159), .ZN(new_n754));
  OAI21_X1  g0554(.A(KEYINPUT32), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n214), .A2(new_n337), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G200), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n343), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G50), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n757), .A2(G190), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI221_X1 g0562(.A(new_n755), .B1(new_n759), .B2(new_n760), .C1(new_n222), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n756), .A2(new_n752), .ZN(new_n764));
  INV_X1    g0564(.A(new_n255), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n756), .A2(G190), .A3(new_n345), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n269), .B1(new_n764), .B2(new_n227), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n343), .A2(G179), .A3(G200), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n214), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G97), .ZN(new_n771));
  OR3_X1    g0571(.A1(new_n753), .A2(new_n754), .A3(KEYINPUT32), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n751), .A2(G190), .A3(G200), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G87), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n751), .A2(new_n343), .A3(G200), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G107), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n771), .A2(new_n772), .A3(new_n775), .A4(new_n778), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n763), .A2(new_n767), .A3(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n766), .ZN(new_n781));
  INV_X1    g0581(.A(new_n753), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n781), .A2(G322), .B1(new_n782), .B2(G329), .ZN(new_n783));
  INV_X1    g0583(.A(G311), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n783), .B(new_n275), .C1(new_n784), .C2(new_n764), .ZN(new_n785));
  INV_X1    g0585(.A(G317), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(KEYINPUT33), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n786), .A2(KEYINPUT33), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n761), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n758), .A2(G326), .ZN(new_n790));
  INV_X1    g0590(.A(G294), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n789), .B(new_n790), .C1(new_n791), .C2(new_n769), .ZN(new_n792));
  INV_X1    g0592(.A(G283), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n793), .A2(new_n776), .B1(new_n773), .B2(new_n592), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n785), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n780), .A2(new_n795), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n729), .B(new_n750), .C1(new_n736), .C2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n735), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n669), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n732), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(G396));
  NAND2_X1  g0601(.A1(new_n646), .A2(new_n666), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n439), .A2(new_n666), .ZN(new_n803));
  AND3_X1   g0603(.A1(new_n448), .A2(new_n450), .A3(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n803), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n804), .B1(new_n451), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n806), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n666), .B(new_n808), .C1(new_n638), .C2(new_n645), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n718), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(new_n727), .B2(new_n728), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n807), .A2(new_n718), .A3(new_n809), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n736), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n734), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(G77), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n729), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n781), .A2(G143), .ZN(new_n818));
  INV_X1    g0618(.A(G150), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n818), .B1(new_n764), .B2(new_n754), .C1(new_n762), .C2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(G137), .B2(new_n758), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n821), .A2(KEYINPUT34), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n821), .A2(KEYINPUT34), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n777), .A2(G68), .ZN(new_n824));
  INV_X1    g0624(.A(G132), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n824), .B(new_n269), .C1(new_n825), .C2(new_n753), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n769), .A2(new_n765), .B1(new_n773), .B2(new_n760), .ZN(new_n827));
  NOR4_X1   g0627(.A1(new_n822), .A2(new_n823), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n764), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n758), .A2(G303), .B1(new_n829), .B2(G116), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n793), .B2(new_n762), .ZN(new_n831));
  XOR2_X1   g0631(.A(new_n831), .B(KEYINPUT104), .Z(new_n832));
  OAI221_X1 g0632(.A(new_n275), .B1(new_n753), .B2(new_n784), .C1(new_n766), .C2(new_n791), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n771), .B1(new_n224), .B2(new_n776), .C1(new_n229), .C2(new_n773), .ZN(new_n834));
  NOR3_X1   g0634(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n828), .A2(new_n835), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n817), .B1(new_n814), .B2(new_n836), .C1(new_n808), .C2(new_n734), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n813), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(G384));
  NOR2_X1   g0639(.A1(new_n724), .A2(new_n257), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n716), .A2(new_n717), .ZN(new_n841));
  INV_X1    g0641(.A(new_n431), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n427), .B(new_n665), .C1(new_n842), .C2(new_n412), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n427), .A2(new_n665), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n428), .A2(new_n431), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n806), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n841), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n350), .A2(new_n262), .ZN(new_n849));
  INV_X1    g0649(.A(new_n295), .ZN(new_n850));
  AOI21_X1  g0650(.A(KEYINPUT16), .B1(new_n289), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n352), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT106), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n663), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n295), .B1(new_n285), .B2(new_n288), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n350), .B(new_n262), .C1(new_n856), .C2(KEYINPUT16), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n857), .A2(KEYINPUT106), .A3(new_n352), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n854), .A2(new_n855), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n854), .A2(new_n359), .A3(new_n858), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n859), .A2(new_n860), .A3(new_n353), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT37), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n360), .A2(new_n855), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT37), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n649), .A2(new_n863), .A3(new_n864), .A4(new_n353), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n859), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n252), .B1(new_n650), .B2(new_n651), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n342), .A2(new_n355), .A3(new_n356), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT38), .B1(new_n866), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n865), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n861), .B2(KEYINPUT37), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n859), .B1(new_n357), .B2(new_n362), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT38), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n848), .B1(new_n871), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT107), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT40), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n353), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n850), .B1(new_n348), .B2(new_n349), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n296), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n853), .B(new_n265), .C1(new_n883), .C2(new_n298), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT106), .B1(new_n857), .B2(new_n352), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n881), .B1(new_n886), .B2(new_n359), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n864), .B1(new_n887), .B2(new_n859), .ZN(new_n888));
  OAI211_X1 g0688(.A(KEYINPUT38), .B(new_n870), .C1(new_n888), .C2(new_n872), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n875), .B1(new_n873), .B2(new_n874), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n847), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT107), .B1(new_n891), .B2(KEYINPUT40), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n650), .A2(new_n651), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n360), .B(new_n855), .C1(new_n893), .C2(new_n655), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n649), .A2(new_n863), .A3(new_n353), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT37), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n865), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n889), .B1(KEYINPUT38), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n841), .A2(new_n846), .A3(KEYINPUT40), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n880), .A2(new_n892), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n453), .B1(new_n717), .B2(new_n716), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n702), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n902), .B2(new_n903), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT39), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n899), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n428), .A2(new_n665), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n889), .A2(new_n890), .A3(KEYINPUT39), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n843), .A2(new_n845), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n652), .A2(new_n665), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n912), .B1(new_n809), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n889), .A2(new_n890), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n915), .A2(new_n916), .B1(new_n893), .B2(new_n663), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n910), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n454), .B1(new_n701), .B2(new_n720), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n658), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n918), .B(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n840), .B1(new_n905), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n921), .B2(new_n905), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n479), .A2(KEYINPUT35), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n479), .A2(KEYINPUT35), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n924), .A2(G116), .A3(new_n215), .A4(new_n925), .ZN(new_n926));
  XOR2_X1   g0726(.A(KEYINPUT105), .B(KEYINPUT36), .Z(new_n927));
  XNOR2_X1  g0727(.A(new_n926), .B(new_n927), .ZN(new_n928));
  OAI211_X1 g0728(.A(G77), .B(new_n217), .C1(new_n765), .C2(new_n222), .ZN(new_n929));
  INV_X1    g0729(.A(new_n201), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n929), .B1(new_n222), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(G1), .A3(new_n723), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n923), .A2(new_n928), .A3(new_n932), .ZN(G367));
  NAND2_X1  g0733(.A1(new_n777), .A2(G77), .ZN(new_n934));
  OAI221_X1 g0734(.A(new_n934), .B1(new_n765), .B2(new_n773), .C1(new_n762), .C2(new_n754), .ZN(new_n935));
  INV_X1    g0735(.A(G143), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n759), .A2(new_n936), .B1(new_n222), .B2(new_n769), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n269), .B1(new_n764), .B2(new_n201), .ZN(new_n938));
  INV_X1    g0738(.A(G137), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n766), .A2(new_n819), .B1(new_n753), .B2(new_n939), .ZN(new_n940));
  NOR4_X1   g0740(.A1(new_n935), .A2(new_n937), .A3(new_n938), .A4(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT112), .ZN(new_n942));
  OAI221_X1 g0742(.A(new_n275), .B1(new_n753), .B2(new_n786), .C1(new_n793), .C2(new_n764), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n762), .A2(new_n791), .B1(new_n776), .B2(new_n483), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n943), .B(new_n944), .C1(G107), .C2(new_n770), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n759), .A2(new_n784), .B1(new_n592), .B2(new_n766), .ZN(new_n946));
  OR3_X1    g0746(.A1(new_n773), .A2(KEYINPUT46), .A3(new_n523), .ZN(new_n947));
  OAI21_X1  g0747(.A(KEYINPUT46), .B1(new_n773), .B2(new_n523), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n946), .A2(KEYINPUT111), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n945), .B(new_n949), .C1(KEYINPUT111), .C2(new_n946), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n942), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT47), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n736), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n539), .A2(new_n665), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n641), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n542), .B2(new_n954), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n735), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n737), .B1(new_n208), .B2(new_n434), .C1(new_n241), .C2(new_n740), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n953), .A2(new_n730), .A3(new_n957), .A4(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n494), .A2(new_n506), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n643), .A2(new_n665), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n642), .A2(new_n961), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n679), .A2(new_n964), .ZN(new_n965));
  XOR2_X1   g0765(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n966));
  XNOR2_X1  g0766(.A(new_n965), .B(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n679), .A2(new_n964), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT44), .ZN(new_n969));
  OR3_X1    g0769(.A1(new_n967), .A2(new_n969), .A3(new_n675), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n675), .B1(new_n967), .B2(new_n969), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n678), .A2(KEYINPUT110), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n676), .A2(new_n673), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n678), .A2(KEYINPUT110), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(new_n670), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n721), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n721), .B1(new_n972), .B2(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n681), .B(KEYINPUT41), .Z(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n726), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n678), .A2(new_n964), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT42), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n964), .B1(new_n584), .B2(new_n585), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n666), .B1(new_n985), .B2(new_n689), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n988));
  NAND2_X1  g0788(.A1(new_n956), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT43), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n987), .B(new_n989), .C1(new_n990), .C2(new_n956), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n987), .B2(new_n989), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n674), .A2(new_n964), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n992), .B(new_n993), .Z(new_n994));
  OAI21_X1  g0794(.A(new_n959), .B1(new_n982), .B2(new_n994), .ZN(G387));
  AOI21_X1  g0795(.A(new_n682), .B1(new_n977), .B2(new_n721), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n721), .B2(new_n977), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n673), .A2(new_n798), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n745), .A2(new_n683), .B1(G107), .B2(new_n208), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n238), .A2(new_n314), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT113), .Z(new_n1001));
  NAND2_X1  g0801(.A1(new_n432), .A2(new_n760), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT50), .Z(new_n1003));
  INV_X1    g0803(.A(new_n683), .ZN(new_n1004));
  AOI211_X1 g0804(.A(G45), .B(new_n1004), .C1(G68), .C2(G77), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n740), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n999), .B1(new_n1001), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n730), .B1(new_n1007), .B2(new_n738), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n770), .A2(new_n507), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n760), .B2(new_n766), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT114), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n776), .A2(new_n483), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n773), .A2(new_n227), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1012), .B(new_n1013), .C1(G159), .C2(new_n758), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n269), .B1(new_n753), .B2(new_n819), .C1(new_n222), .C2(new_n764), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(new_n256), .B2(new_n761), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1011), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n766), .A2(new_n786), .B1(new_n764), .B2(new_n592), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1018), .A2(KEYINPUT115), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(KEYINPUT115), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n761), .A2(G311), .B1(new_n758), .B2(G322), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT48), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n769), .A2(new_n793), .B1(new_n773), .B2(new_n791), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1024), .A2(KEYINPUT49), .A3(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n269), .B1(new_n782), .B2(G326), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1027), .B(new_n1028), .C1(new_n523), .C2(new_n776), .ZN(new_n1029));
  AOI21_X1  g0829(.A(KEYINPUT49), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1017), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1008), .B1(new_n736), .B2(new_n1031), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n977), .A2(new_n726), .B1(new_n998), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n997), .A2(new_n1033), .ZN(G393));
  OR2_X1    g0834(.A1(new_n972), .A2(new_n978), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n972), .A2(new_n978), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1035), .A2(new_n681), .A3(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n972), .A2(new_n725), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n964), .A2(new_n735), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n737), .B1(new_n483), .B2(new_n208), .C1(new_n245), .C2(new_n740), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n730), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n759), .A2(new_n786), .B1(new_n784), .B2(new_n766), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT52), .Z(new_n1043));
  AOI21_X1  g0843(.A(new_n269), .B1(new_n782), .B2(G322), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n791), .B2(new_n764), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n778), .B1(new_n762), .B2(new_n592), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n769), .A2(new_n523), .B1(new_n773), .B2(new_n793), .ZN(new_n1047));
  OR4_X1    g0847(.A1(new_n1043), .A2(new_n1045), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT116), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(G159), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n759), .A2(new_n819), .B1(new_n1051), .B2(new_n766), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT51), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n269), .B1(new_n753), .B2(new_n936), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n432), .B2(new_n829), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n761), .A2(new_n930), .B1(new_n777), .B2(G87), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n769), .A2(new_n227), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(G68), .B2(new_n774), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .A4(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1050), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1041), .B1(new_n1061), .B2(new_n736), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1038), .B1(new_n1039), .B2(new_n1062), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1037), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(G390));
  NAND2_X1  g0865(.A1(new_n718), .A2(new_n808), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n912), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n718), .A2(new_n808), .A3(new_n911), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n809), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1069), .B1(new_n1070), .B2(new_n913), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n700), .A2(new_n666), .A3(new_n808), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1067), .A2(new_n914), .A3(new_n1068), .A4(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n454), .A2(new_n718), .ZN(new_n1075));
  AND3_X1   g0875(.A1(new_n919), .A2(new_n658), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n915), .A2(new_n908), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n907), .B2(new_n909), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n899), .B1(new_n428), .B2(new_n665), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n912), .B1(new_n1072), .B2(new_n914), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1068), .ZN(new_n1083));
  NOR3_X1   g0883(.A1(new_n1079), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1085));
  AOI21_X1  g0885(.A(KEYINPUT38), .B1(new_n894), .B2(new_n897), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n873), .A2(new_n874), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1086), .B1(new_n1087), .B2(KEYINPUT38), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1088), .A2(KEYINPUT39), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n909), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n1089), .A2(new_n1090), .B1(new_n915), .B2(new_n908), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1068), .B1(new_n1085), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1077), .B1(new_n1084), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1085), .A2(new_n1091), .A3(new_n1068), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1083), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1094), .A2(new_n1095), .A3(new_n1076), .A4(new_n1074), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1093), .A2(new_n681), .A3(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1094), .A2(new_n1095), .A3(new_n726), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n733), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n730), .B1(new_n256), .B2(new_n815), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n764), .A2(new_n483), .B1(new_n753), .B2(new_n791), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n269), .B(new_n1101), .C1(G116), .C2(new_n781), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1102), .A2(new_n775), .A3(new_n824), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1057), .B1(G283), .B2(new_n758), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n229), .B2(new_n762), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n774), .A2(G150), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT53), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G159), .A2(new_n770), .B1(new_n758), .B2(G128), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n275), .B1(new_n782), .B2(G125), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(KEYINPUT54), .B(G143), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n781), .A2(G132), .B1(new_n829), .B2(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n761), .A2(G137), .B1(new_n777), .B2(new_n930), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1108), .A2(new_n1109), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n1103), .A2(new_n1105), .B1(new_n1107), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1100), .B1(new_n1115), .B2(new_n736), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1099), .A2(new_n1116), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n1098), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1097), .A2(new_n1118), .ZN(G378));
  INV_X1    g0919(.A(new_n918), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n369), .A2(new_n855), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT55), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n389), .B(new_n1122), .ZN(new_n1123));
  XOR2_X1   g0923(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  OR2_X1    g0925(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n880), .A2(new_n892), .ZN(new_n1130));
  OAI21_X1  g0930(.A(G330), .B1(new_n1088), .B2(new_n900), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1129), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1128), .B(new_n1131), .C1(new_n880), .C2(new_n892), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1120), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n878), .B1(new_n877), .B2(new_n879), .ZN(new_n1136));
  NOR3_X1   g0936(.A1(new_n891), .A2(KEYINPUT107), .A3(KEYINPUT40), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1132), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n1128), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1130), .A2(new_n1132), .A3(new_n1129), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1139), .A2(new_n918), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT119), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1135), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  OAI211_X1 g0943(.A(KEYINPUT119), .B(new_n1120), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1096), .A2(new_n1076), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT57), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT120), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1146), .A2(KEYINPUT120), .A3(new_n1147), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1147), .B1(new_n1096), .B2(new_n1076), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1135), .A2(new_n1141), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n682), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1150), .A2(new_n1151), .A3(new_n1154), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1129), .A2(new_n733), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n730), .B1(new_n930), .B2(new_n815), .ZN(new_n1158));
  AOI211_X1 g0958(.A(G33), .B(G41), .C1(new_n782), .C2(G124), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n776), .B2(new_n754), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n758), .A2(G125), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n762), .B2(new_n825), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n781), .A2(G128), .B1(new_n829), .B2(G137), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n773), .B2(new_n1110), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1162), .B(new_n1164), .C1(G150), .C2(new_n770), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1160), .B1(new_n1166), .B2(KEYINPUT59), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(KEYINPUT59), .B2(new_n1166), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n758), .A2(G116), .B1(new_n777), .B2(new_n255), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n483), .B2(new_n762), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n766), .A2(new_n229), .B1(new_n753), .B2(new_n793), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n313), .B(new_n275), .C1(new_n764), .C2(new_n434), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n769), .A2(new_n222), .B1(new_n773), .B2(new_n227), .ZN(new_n1173));
  NOR4_X1   g0973(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1174), .B(KEYINPUT58), .Z(new_n1175));
  AOI21_X1  g0975(.A(G50), .B1(new_n273), .B2(new_n313), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n269), .B2(G41), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1168), .A2(new_n1175), .A3(new_n1177), .ZN(new_n1178));
  OR2_X1    g0978(.A1(new_n1178), .A2(KEYINPUT117), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n814), .B1(new_n1178), .B2(KEYINPUT117), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1158), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1156), .A2(new_n726), .B1(new_n1157), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1155), .A2(new_n1182), .ZN(G375));
  NAND2_X1  g0983(.A1(new_n912), .A2(new_n733), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n730), .B1(G68), .B2(new_n815), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n523), .A2(new_n762), .B1(new_n759), .B2(new_n791), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(G97), .B2(new_n774), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n766), .A2(new_n793), .B1(new_n764), .B2(new_n229), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n269), .B(new_n1188), .C1(G303), .C2(new_n782), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1187), .A2(new_n934), .A3(new_n1009), .A4(new_n1189), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n769), .A2(new_n760), .B1(new_n773), .B2(new_n1051), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(G132), .B2(new_n758), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n275), .B1(new_n782), .B2(G128), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n781), .A2(G137), .B1(new_n829), .B2(G150), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n761), .A2(new_n1111), .B1(new_n777), .B2(new_n255), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1190), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1185), .B1(new_n1197), .B2(new_n736), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n1074), .A2(new_n726), .B1(new_n1184), .B2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT121), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1077), .A2(new_n981), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1199), .B1(new_n1201), .B2(new_n1202), .ZN(G381));
  INV_X1    g1003(.A(G378), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1155), .A2(new_n1204), .A3(new_n1182), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n997), .A2(new_n800), .A3(new_n1033), .ZN(new_n1206));
  OR3_X1    g1006(.A1(G390), .A2(G384), .A3(new_n1206), .ZN(new_n1207));
  OR4_X1    g1007(.A1(G387), .A2(new_n1205), .A3(G381), .A4(new_n1207), .ZN(G407));
  OAI211_X1 g1008(.A(G407), .B(G213), .C1(G343), .C2(new_n1205), .ZN(G409));
  AND2_X1   g1009(.A1(new_n664), .A2(G213), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1155), .A2(G378), .A3(new_n1182), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1143), .A2(new_n1145), .A3(new_n981), .A4(new_n1144), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1153), .A2(new_n726), .B1(new_n1157), .B2(new_n1181), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n1214), .A2(KEYINPUT122), .A3(new_n1204), .ZN(new_n1215));
  AOI21_X1  g1015(.A(KEYINPUT122), .B1(new_n1214), .B2(new_n1204), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1210), .B1(new_n1211), .B2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n682), .B1(new_n1200), .B2(KEYINPUT60), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1077), .A2(KEYINPUT60), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1219), .B1(new_n1201), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n1199), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(G384), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1218), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT63), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  OR2_X1    g1026(.A1(new_n1064), .A2(G387), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1064), .A2(G387), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(G393), .A2(G396), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1230), .A2(new_n1206), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1231), .A2(KEYINPUT123), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(KEYINPUT123), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1229), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n1234), .A2(KEYINPUT124), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT125), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1064), .A2(G387), .A3(new_n1237), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1227), .A2(new_n1236), .A3(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1228), .A2(KEYINPUT125), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1234), .A2(KEYINPUT124), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(KEYINPUT61), .B1(new_n1235), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1210), .A2(G2897), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1223), .B(new_n1243), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1244), .A2(new_n1218), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1222), .B(new_n838), .ZN(new_n1246));
  AOI211_X1 g1046(.A(new_n1210), .B(new_n1246), .C1(new_n1211), .C2(new_n1217), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(KEYINPUT63), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1226), .A2(new_n1242), .A3(new_n1245), .A4(new_n1248), .ZN(new_n1249));
  XOR2_X1   g1049(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n1244), .B2(new_n1218), .ZN(new_n1251));
  AND2_X1   g1051(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1252), .B1(new_n1247), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1224), .A2(new_n1253), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1251), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1235), .A2(new_n1241), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1249), .B1(new_n1257), .B2(new_n1258), .ZN(G405));
  NAND2_X1  g1059(.A1(G375), .A2(new_n1204), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1260), .A2(new_n1211), .A3(new_n1246), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1246), .B1(new_n1260), .B2(new_n1211), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1263), .B(new_n1258), .ZN(G402));
endmodule


