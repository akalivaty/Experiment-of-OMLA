//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n845, new_n846, new_n847, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965;
  INV_X1    g000(.A(KEYINPUT40), .ZN(new_n202));
  XOR2_X1   g001(.A(G127gat), .B(G134gat), .Z(new_n203));
  INV_X1    g002(.A(KEYINPUT68), .ZN(new_n204));
  XOR2_X1   g003(.A(G113gat), .B(G120gat), .Z(new_n205));
  AOI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT1), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  OR2_X1    g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n206), .A2(new_n208), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G155gat), .ZN(new_n213));
  INV_X1    g012(.A(G162gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n216));
  NOR2_X1   g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  XOR2_X1   g017(.A(KEYINPUT75), .B(G141gat), .Z(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G148gat), .ZN(new_n220));
  INV_X1    g019(.A(G148gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G141gat), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n218), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(G141gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G148gat), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT2), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  NOR3_X1   g025(.A1(new_n226), .A2(new_n215), .A3(new_n217), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n223), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G225gat), .A2(G233gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n231), .B(KEYINPUT76), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n211), .A2(new_n228), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n230), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT39), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n228), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT3), .B1(new_n223), .B2(new_n227), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n212), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT4), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n234), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n211), .A2(KEYINPUT4), .A3(new_n228), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n240), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n236), .B1(new_n232), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT39), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n244), .A2(new_n246), .A3(new_n232), .ZN(new_n247));
  XNOR2_X1  g046(.A(G1gat), .B(G29gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(KEYINPUT0), .ZN(new_n249));
  XNOR2_X1  g048(.A(G57gat), .B(G85gat), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n249), .B(new_n250), .Z(new_n251));
  NAND2_X1  g050(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n202), .B1(new_n245), .B2(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n233), .B1(new_n230), .B2(new_n234), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT5), .ZN(new_n255));
  OAI22_X1  g054(.A1(new_n244), .A2(new_n232), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n242), .A2(new_n243), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n257), .A2(KEYINPUT5), .A3(new_n233), .A4(new_n240), .ZN(new_n258));
  INV_X1    g057(.A(new_n251), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n256), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n232), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n261), .A2(KEYINPUT39), .A3(new_n235), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n262), .A2(KEYINPUT40), .A3(new_n251), .A4(new_n247), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n253), .A2(new_n260), .A3(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G8gat), .B(G36gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(G64gat), .B(G92gat), .ZN(new_n266));
  XOR2_X1   g065(.A(new_n265), .B(new_n266), .Z(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G226gat), .A2(G233gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT64), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n273));
  INV_X1    g072(.A(G183gat), .ZN(new_n274));
  INV_X1    g073(.A(G190gat), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  OR2_X1    g076(.A1(new_n277), .A2(KEYINPUT65), .ZN(new_n278));
  NOR2_X1   g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  OR2_X1    g078(.A1(new_n279), .A2(KEYINPUT23), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(KEYINPUT23), .ZN(new_n281));
  NAND2_X1  g080(.A1(G169gat), .A2(G176gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n283), .B1(new_n277), .B2(KEYINPUT65), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n278), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT25), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n283), .A2(new_n286), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n276), .A2(new_n270), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT27), .B(G183gat), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT66), .B1(new_n292), .B2(new_n275), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n293), .A2(KEYINPUT28), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n294), .B1(G183gat), .B2(G190gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT26), .ZN(new_n296));
  NOR4_X1   g095(.A1(KEYINPUT67), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT67), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n298), .B1(new_n279), .B2(new_n296), .ZN(new_n299));
  OAI221_X1 g098(.A(new_n282), .B1(new_n296), .B2(new_n279), .C1(new_n297), .C2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n293), .A2(KEYINPUT28), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n295), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n269), .B1(new_n291), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT29), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n285), .A2(new_n286), .B1(new_n289), .B2(new_n288), .ZN(new_n307));
  INV_X1    g106(.A(new_n303), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(new_n269), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT72), .B(G197gat), .ZN(new_n311));
  INV_X1    g110(.A(G204gat), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n311), .A2(new_n312), .ZN(new_n314));
  AND2_X1   g113(.A1(G211gat), .A2(G218gat), .ZN(new_n315));
  OAI22_X1  g114(.A1(new_n313), .A2(new_n314), .B1(KEYINPUT22), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(KEYINPUT73), .ZN(new_n317));
  NOR2_X1   g116(.A1(G211gat), .A2(G218gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  OR2_X1    g119(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n317), .A2(new_n320), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n305), .A2(new_n310), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT74), .B(KEYINPUT29), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n326), .B1(new_n307), .B2(new_n308), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(new_n269), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n323), .B1(new_n305), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n268), .B1(new_n325), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n304), .B1(new_n327), .B2(new_n269), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n324), .B(new_n267), .C1(new_n331), .C2(new_n323), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n330), .A2(KEYINPUT30), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n329), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT30), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n334), .A2(new_n335), .A3(new_n267), .A4(new_n324), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n264), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(G228gat), .A2(G233gat), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n238), .A2(new_n326), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n321), .A2(new_n322), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT3), .B1(new_n323), .B2(new_n306), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n339), .B(new_n341), .C1(new_n342), .C2(new_n228), .ZN(new_n343));
  XNOR2_X1  g142(.A(G78gat), .B(G106gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT31), .B(G50gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(G22gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n347), .A2(KEYINPUT77), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n348), .B1(new_n350), .B2(new_n346), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n326), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n353), .B1(new_n321), .B2(new_n322), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n229), .B1(new_n354), .B2(KEYINPUT3), .ZN(new_n355));
  AND2_X1   g154(.A1(new_n355), .A2(new_n341), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n343), .B(new_n352), .C1(new_n356), .C2(new_n339), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n339), .ZN(new_n358));
  INV_X1    g157(.A(new_n342), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n358), .B1(new_n359), .B2(new_n229), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n339), .B1(new_n355), .B2(new_n341), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n351), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AND2_X1   g161(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n337), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n256), .A2(new_n258), .A3(KEYINPUT6), .A4(new_n259), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n366), .A2(KEYINPUT79), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT6), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n260), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n259), .B1(new_n256), .B2(new_n258), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n365), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n367), .B1(new_n371), .B2(KEYINPUT79), .ZN(new_n372));
  INV_X1    g171(.A(new_n323), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n373), .A2(new_n305), .A3(new_n310), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n374), .B(KEYINPUT37), .C1(new_n331), .C2(new_n373), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT78), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT38), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n268), .A2(KEYINPUT37), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n330), .A2(new_n378), .ZN(new_n379));
  OR2_X1    g178(.A1(new_n331), .A2(new_n373), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n380), .A2(KEYINPUT78), .A3(KEYINPUT37), .A4(new_n374), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n377), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n324), .B1(new_n331), .B2(new_n323), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n383), .A2(KEYINPUT37), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n268), .B1(new_n383), .B2(KEYINPUT37), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT38), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n372), .A2(new_n382), .A3(new_n386), .A4(new_n332), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT80), .B1(new_n364), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT36), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n291), .A2(new_n212), .A3(new_n303), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n211), .B1(new_n307), .B2(new_n308), .ZN(new_n391));
  INV_X1    g190(.A(G227gat), .ZN(new_n392));
  INV_X1    g191(.A(G233gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n390), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(KEYINPUT69), .B(KEYINPUT33), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n395), .A2(KEYINPUT32), .ZN(new_n398));
  XOR2_X1   g197(.A(G15gat), .B(G43gat), .Z(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT70), .ZN(new_n400));
  XNOR2_X1  g199(.A(G71gat), .B(G99gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n397), .A2(new_n398), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n396), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n403), .B(KEYINPUT71), .C1(new_n398), .C2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT71), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n397), .A2(new_n398), .A3(new_n407), .A4(new_n402), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n390), .A2(new_n391), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n409), .B1(new_n392), .B2(new_n393), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n410), .A2(KEYINPUT34), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n410), .A2(KEYINPUT34), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n406), .A2(new_n408), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n413), .B1(new_n406), .B2(new_n408), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n389), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n333), .A2(new_n336), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n371), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n357), .A2(new_n362), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n403), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT71), .B1(new_n398), .B2(new_n405), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n408), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n424), .B1(new_n411), .B2(new_n412), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n425), .A2(KEYINPUT36), .A3(new_n414), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n417), .A2(new_n421), .A3(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n388), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n364), .A2(new_n387), .A3(KEYINPUT80), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n425), .A2(new_n414), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n430), .A2(new_n418), .A3(new_n363), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n372), .A2(KEYINPUT35), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n430), .A2(new_n371), .A3(new_n418), .A4(new_n363), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT35), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n428), .A2(new_n429), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(G229gat), .A2(G233gat), .ZN(new_n438));
  XOR2_X1   g237(.A(new_n438), .B(KEYINPUT13), .Z(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(G50gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT83), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT83), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(G50gat), .ZN(new_n444));
  INV_X1    g243(.A(G43gat), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n442), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(G43gat), .A2(G50gat), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT15), .ZN(new_n448));
  OR2_X1    g247(.A1(new_n448), .A2(KEYINPUT82), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(KEYINPUT82), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n446), .A2(new_n447), .A3(new_n449), .A4(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n445), .A2(new_n441), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n447), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT15), .ZN(new_n454));
  INV_X1    g253(.A(G36gat), .ZN(new_n455));
  AND2_X1   g254(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n456));
  NOR2_X1   g255(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(G29gat), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n459), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n451), .A2(new_n454), .A3(new_n461), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n459), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT14), .B(G29gat), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n463), .B1(new_n464), .B2(new_n455), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n448), .B1(new_n452), .B2(new_n447), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT81), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AND4_X1   g266(.A1(KEYINPUT81), .A2(new_n466), .A3(new_n458), .A4(new_n460), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n347), .A2(G15gat), .ZN(new_n470));
  INV_X1    g269(.A(G15gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(G22gat), .ZN(new_n472));
  AOI21_X1  g271(.A(G1gat), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT86), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n473), .B1(new_n474), .B2(G8gat), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT84), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT16), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n477), .B1(new_n478), .B2(G1gat), .ZN(new_n479));
  INV_X1    g278(.A(G1gat), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n480), .A2(KEYINPUT84), .A3(KEYINPUT16), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(G15gat), .B(G22gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT87), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT87), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n482), .A2(new_n486), .A3(new_n483), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(G8gat), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n476), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT85), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n484), .A2(new_n491), .B1(new_n474), .B2(new_n473), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n482), .A2(KEYINPUT85), .A3(new_n483), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n489), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n469), .B1(new_n490), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n487), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n486), .B1(new_n482), .B2(new_n483), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n489), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n475), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n491), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n473), .A2(new_n474), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n500), .A2(new_n493), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(G8gat), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT81), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n504), .B1(new_n461), .B2(new_n454), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n465), .A2(KEYINPUT81), .A3(new_n466), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n466), .B1(new_n458), .B2(new_n460), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n505), .A2(new_n506), .B1(new_n507), .B2(new_n451), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n499), .A2(new_n503), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n440), .B1(new_n495), .B2(new_n509), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n462), .B(KEYINPUT17), .C1(new_n467), .C2(new_n468), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n499), .A2(new_n511), .A3(new_n503), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n508), .A2(KEYINPUT17), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n495), .B(new_n438), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT18), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n510), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G113gat), .B(G141gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n517), .B(G197gat), .ZN(new_n518));
  XOR2_X1   g317(.A(KEYINPUT11), .B(G169gat), .Z(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(KEYINPUT12), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n490), .A2(new_n494), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT17), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n469), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n522), .A2(new_n524), .A3(new_n511), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n525), .A2(KEYINPUT18), .A3(new_n438), .A4(new_n495), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n516), .A2(new_n521), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n521), .B1(new_n516), .B2(new_n526), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n437), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT90), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(G134gat), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT91), .ZN(new_n535));
  AND3_X1   g334(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT92), .ZN(new_n537));
  AND2_X1   g336(.A1(G99gat), .A2(G106gat), .ZN(new_n538));
  NOR2_X1   g337(.A1(G99gat), .A2(G106gat), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(G99gat), .ZN(new_n541));
  INV_X1    g340(.A(G106gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(G99gat), .A2(G106gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n543), .A2(KEYINPUT92), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT93), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n540), .A2(new_n545), .A3(KEYINPUT93), .ZN(new_n549));
  NAND2_X1  g348(.A1(G85gat), .A2(G92gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT7), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT7), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n552), .A2(G85gat), .A3(G92gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(G85gat), .ZN(new_n555));
  INV_X1    g354(.A(G92gat), .ZN(new_n556));
  AOI22_X1  g355(.A1(KEYINPUT8), .A2(new_n544), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n548), .A2(new_n549), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n554), .A2(new_n557), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n546), .A2(new_n560), .A3(new_n547), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n536), .B1(new_n562), .B2(new_n469), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n511), .A2(new_n561), .A3(new_n559), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n563), .B1(new_n564), .B2(new_n513), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(G190gat), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n559), .A2(new_n561), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n524), .A2(new_n511), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n568), .A2(new_n275), .A3(new_n563), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(G218gat), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n535), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n566), .A2(G218gat), .A3(new_n569), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n214), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n568), .A2(new_n275), .A3(new_n563), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n275), .B1(new_n568), .B2(new_n563), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n571), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n577), .A2(new_n573), .A3(KEYINPUT91), .A4(new_n214), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n534), .B1(new_n574), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n577), .A2(KEYINPUT91), .A3(new_n573), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(G162gat), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n582), .A2(new_n533), .A3(new_n578), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(G71gat), .A2(G78gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT9), .ZN(new_n586));
  NAND2_X1  g385(.A1(G71gat), .A2(G78gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT89), .ZN(new_n589));
  NAND2_X1  g388(.A1(G57gat), .A2(G64gat), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(G57gat), .A2(G64gat), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n589), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  OR2_X1    g392(.A1(G57gat), .A2(G64gat), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n594), .A2(KEYINPUT89), .A3(new_n590), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n588), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT88), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n587), .B1(new_n585), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(KEYINPUT88), .A2(G71gat), .A3(G78gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n594), .A2(new_n590), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n598), .B(new_n599), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n596), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT21), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G231gat), .A2(G233gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n607), .B(G127gat), .Z(new_n608));
  OAI21_X1  g407(.A(new_n522), .B1(new_n604), .B2(new_n603), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(G155gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(G183gat), .B(G211gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n610), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n584), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT94), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n584), .A2(new_n615), .A3(KEYINPUT94), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n559), .A2(new_n603), .A3(new_n561), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n596), .A2(new_n602), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT95), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n546), .B1(new_n558), .B2(new_n626), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n560), .A2(KEYINPUT95), .A3(new_n540), .A4(new_n545), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n625), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g428(.A(KEYINPUT96), .B(KEYINPUT10), .Z(new_n630));
  NAND3_X1  g429(.A1(new_n624), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n562), .A2(KEYINPUT10), .A3(new_n625), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n623), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT97), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n624), .A2(new_n629), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n634), .B1(new_n635), .B2(new_n623), .ZN(new_n636));
  AOI211_X1 g435(.A(KEYINPUT97), .B(new_n622), .C1(new_n624), .C2(new_n629), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n633), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(G120gat), .B(G148gat), .Z(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT98), .ZN(new_n640));
  XNOR2_X1  g439(.A(G176gat), .B(G204gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n642), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n622), .B1(new_n624), .B2(new_n629), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(new_n634), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n644), .B1(new_n646), .B2(new_n633), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  NOR3_X1   g447(.A1(new_n619), .A2(new_n621), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n530), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n650), .A2(new_n371), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(new_n480), .ZN(G1324gat));
  NOR2_X1   g451(.A1(new_n650), .A2(new_n418), .ZN(new_n653));
  XOR2_X1   g452(.A(KEYINPUT16), .B(G8gat), .Z(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n655), .B1(new_n489), .B2(new_n653), .ZN(new_n656));
  MUX2_X1   g455(.A(new_n655), .B(new_n656), .S(KEYINPUT42), .Z(G1325gat));
  AND2_X1   g456(.A1(new_n417), .A2(new_n426), .ZN(new_n658));
  OAI21_X1  g457(.A(G15gat), .B1(new_n650), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n430), .A2(new_n471), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n659), .B1(new_n650), .B2(new_n660), .ZN(G1326gat));
  NAND3_X1  g460(.A1(new_n530), .A2(new_n420), .A3(new_n649), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n662), .A2(KEYINPUT99), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(KEYINPUT99), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT43), .B(G22gat), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n665), .B(new_n666), .Z(G1327gat));
  NOR3_X1   g466(.A1(new_n584), .A2(new_n615), .A3(new_n648), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n530), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n371), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n669), .A2(new_n459), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT45), .ZN(new_n672));
  AND3_X1   g471(.A1(new_n364), .A2(new_n387), .A3(KEYINPUT80), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n673), .A2(new_n388), .A3(new_n427), .ZN(new_n674));
  AOI22_X1  g473(.A1(new_n432), .A2(new_n433), .B1(new_n435), .B2(KEYINPUT35), .ZN(new_n675));
  OAI21_X1  g474(.A(KEYINPUT100), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n364), .A2(new_n387), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT80), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n679), .A2(new_n658), .A3(new_n429), .A4(new_n421), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n434), .A2(new_n436), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT100), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n584), .A2(KEYINPUT44), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n676), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(KEYINPUT44), .B1(new_n437), .B2(new_n584), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n615), .ZN(new_n688));
  INV_X1    g487(.A(new_n529), .ZN(new_n689));
  INV_X1    g488(.A(new_n648), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n687), .A2(new_n371), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n672), .B1(new_n692), .B2(new_n459), .ZN(G1328gat));
  INV_X1    g492(.A(KEYINPUT101), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n687), .A2(new_n418), .A3(new_n691), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(new_n455), .ZN(new_n696));
  INV_X1    g495(.A(new_n418), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n530), .A2(new_n455), .A3(new_n697), .A4(new_n668), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT46), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n694), .B1(new_n696), .B2(new_n699), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n698), .B(KEYINPUT46), .Z(new_n701));
  OAI211_X1 g500(.A(new_n701), .B(KEYINPUT101), .C1(new_n455), .C2(new_n695), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n702), .ZN(G1329gat));
  AND3_X1   g502(.A1(new_n669), .A2(new_n445), .A3(new_n430), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT47), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AOI211_X1 g505(.A(new_n658), .B(new_n691), .C1(new_n685), .C2(new_n686), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n707), .A2(KEYINPUT103), .ZN(new_n708));
  OAI21_X1  g507(.A(G43gat), .B1(new_n707), .B2(KEYINPUT103), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n706), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT102), .B(KEYINPUT47), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n707), .A2(new_n445), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n711), .B1(new_n712), .B2(new_n704), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n710), .A2(new_n713), .ZN(G1330gat));
  AND2_X1   g513(.A1(new_n442), .A2(new_n444), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n420), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g515(.A(new_n716), .B(KEYINPUT104), .Z(new_n717));
  NAND2_X1  g516(.A1(new_n669), .A2(new_n717), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n687), .A2(new_n363), .A3(new_n691), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n719), .B2(new_n715), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT48), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OAI211_X1 g521(.A(KEYINPUT48), .B(new_n718), .C1(new_n719), .C2(new_n715), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(G1331gat));
  AND2_X1   g523(.A1(new_n676), .A2(new_n683), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n689), .A2(new_n690), .ZN(new_n726));
  AND3_X1   g525(.A1(new_n618), .A2(new_n620), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(new_n371), .ZN(new_n729));
  XOR2_X1   g528(.A(KEYINPUT105), .B(G57gat), .Z(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(G1332gat));
  NOR2_X1   g530(.A1(new_n728), .A2(new_n418), .ZN(new_n732));
  NOR2_X1   g531(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n733));
  AND2_X1   g532(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n735), .B1(new_n732), .B2(new_n733), .ZN(G1333gat));
  INV_X1    g535(.A(new_n430), .ZN(new_n737));
  OR3_X1    g536(.A1(new_n728), .A2(G71gat), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(G71gat), .B1(new_n728), .B2(new_n658), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT50), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n738), .A2(KEYINPUT50), .A3(new_n739), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(G1334gat));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n363), .ZN(new_n745));
  XNOR2_X1  g544(.A(KEYINPUT106), .B(G78gat), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1335gat));
  NAND2_X1  g546(.A1(new_n685), .A2(new_n686), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n688), .A2(new_n726), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT107), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(G85gat), .B1(new_n751), .B2(new_n371), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n680), .A2(new_n681), .ZN(new_n753));
  INV_X1    g552(.A(new_n584), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n615), .A2(new_n689), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n753), .A2(KEYINPUT51), .A3(new_n754), .A4(new_n755), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n690), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n760), .A2(new_n555), .A3(new_n670), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n752), .A2(new_n761), .ZN(G1336gat));
  NOR2_X1   g561(.A1(new_n418), .A2(G92gat), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT108), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n760), .A2(new_n763), .B1(new_n764), .B2(KEYINPUT52), .ZN(new_n765));
  OAI21_X1  g564(.A(G92gat), .B1(new_n751), .B2(new_n418), .ZN(new_n766));
  OR2_X1    g565(.A1(new_n764), .A2(KEYINPUT52), .ZN(new_n767));
  AND3_X1   g566(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n767), .B1(new_n765), .B2(new_n766), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n768), .A2(new_n769), .ZN(G1337gat));
  OAI21_X1  g569(.A(G99gat), .B1(new_n751), .B2(new_n658), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n760), .A2(new_n541), .A3(new_n430), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(G1338gat));
  NOR2_X1   g572(.A1(new_n363), .A2(G106gat), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n760), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n750), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n776), .B1(new_n685), .B2(new_n686), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n542), .B1(new_n777), .B2(new_n420), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n775), .B1(new_n778), .B2(KEYINPUT109), .ZN(new_n779));
  AOI211_X1 g578(.A(new_n363), .B(new_n776), .C1(new_n685), .C2(new_n686), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT109), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n780), .A2(new_n781), .A3(new_n542), .ZN(new_n782));
  OAI21_X1  g581(.A(KEYINPUT53), .B1(new_n779), .B2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT110), .ZN(new_n785));
  OAI21_X1  g584(.A(G106gat), .B1(new_n780), .B2(new_n785), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n751), .A2(KEYINPUT110), .A3(new_n363), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n784), .B(new_n775), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n783), .A2(new_n788), .ZN(G1339gat));
  NAND4_X1  g588(.A1(new_n618), .A2(new_n529), .A3(new_n620), .A4(new_n690), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n582), .A2(new_n533), .A3(new_n578), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n533), .B1(new_n582), .B2(new_n578), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n631), .A2(new_n623), .A3(new_n632), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT111), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n631), .A2(new_n632), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n622), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n631), .A2(new_n632), .A3(KEYINPUT111), .A4(new_n623), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n795), .A2(new_n797), .A3(KEYINPUT54), .A4(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n642), .B1(new_n633), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AOI211_X1 g603(.A(new_n803), .B(new_n642), .C1(new_n633), .C2(new_n800), .ZN(new_n805));
  AOI22_X1  g604(.A1(new_n805), .A2(new_n799), .B1(new_n638), .B2(new_n642), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n495), .A2(new_n509), .A3(new_n440), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT112), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n495), .A2(new_n509), .A3(KEYINPUT112), .A4(new_n440), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n525), .A2(new_n495), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n809), .B(new_n810), .C1(new_n811), .C2(new_n438), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n520), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n516), .A2(new_n521), .A3(new_n526), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n804), .A2(new_n806), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n791), .A2(new_n792), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n813), .A2(new_n648), .A3(new_n814), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n804), .A2(new_n806), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n817), .B1(new_n818), .B2(new_n529), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT113), .ZN(new_n820));
  AOI22_X1  g619(.A1(new_n819), .A2(new_n820), .B1(new_n580), .B2(new_n583), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n817), .B(KEYINPUT113), .C1(new_n818), .C2(new_n529), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n816), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n688), .B1(new_n823), .B2(KEYINPUT114), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT114), .ZN(new_n825));
  AOI211_X1 g624(.A(new_n825), .B(new_n816), .C1(new_n822), .C2(new_n821), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n790), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n828), .A2(new_n371), .A3(new_n431), .ZN(new_n829));
  AOI21_X1  g628(.A(G113gat), .B1(new_n829), .B2(new_n689), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n828), .A2(new_n420), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n697), .A2(new_n371), .ZN(new_n832));
  AND3_X1   g631(.A1(new_n831), .A2(new_n430), .A3(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n689), .A2(G113gat), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n830), .B1(new_n833), .B2(new_n834), .ZN(G1340gat));
  AOI21_X1  g634(.A(G120gat), .B1(new_n829), .B2(new_n648), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n648), .A2(G120gat), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n836), .B1(new_n833), .B2(new_n837), .ZN(G1341gat));
  AND3_X1   g637(.A1(new_n833), .A2(G127gat), .A3(new_n615), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n829), .A2(new_n615), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n841), .A2(KEYINPUT115), .ZN(new_n842));
  AOI21_X1  g641(.A(G127gat), .B1(new_n841), .B2(KEYINPUT115), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n839), .B1(new_n842), .B2(new_n843), .ZN(G1342gat));
  AND2_X1   g643(.A1(new_n833), .A2(new_n754), .ZN(new_n845));
  INV_X1    g644(.A(G134gat), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n829), .A2(new_n846), .A3(new_n754), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n847), .B1(KEYINPUT56), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n849), .B1(KEYINPUT56), .B2(new_n848), .ZN(G1343gat));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n827), .A2(new_n420), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n851), .B1(new_n852), .B2(KEYINPUT57), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT57), .B1(new_n827), .B2(new_n420), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT116), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n689), .A2(new_n806), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n802), .A2(KEYINPUT117), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n802), .A2(KEYINPUT117), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n857), .A2(new_n858), .A3(KEYINPUT55), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n817), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n584), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(KEYINPUT118), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT118), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n816), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n615), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n790), .ZN(new_n867));
  OAI211_X1 g666(.A(KEYINPUT57), .B(new_n420), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n853), .A2(new_n855), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n658), .A2(new_n832), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n869), .A2(KEYINPUT121), .A3(new_n689), .A4(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n868), .B1(new_n854), .B2(KEYINPUT116), .ZN(new_n873));
  AOI211_X1 g672(.A(new_n851), .B(KEYINPUT57), .C1(new_n827), .C2(new_n420), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n689), .B(new_n871), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT121), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(new_n219), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n872), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n658), .A2(new_n420), .ZN(new_n880));
  NOR4_X1   g679(.A1(new_n828), .A2(new_n371), .A3(new_n697), .A4(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n224), .A3(new_n689), .ZN(new_n882));
  XOR2_X1   g681(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n883));
  NAND3_X1  g682(.A1(new_n879), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n875), .A2(new_n885), .A3(new_n878), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n885), .B1(new_n875), .B2(new_n878), .ZN(new_n887));
  INV_X1    g686(.A(new_n882), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT58), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n884), .B1(new_n889), .B2(new_n890), .ZN(G1344gat));
  NAND3_X1  g690(.A1(new_n881), .A2(new_n221), .A3(new_n648), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n867), .A2(KEYINPUT122), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n867), .A2(KEYINPUT122), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n688), .B1(new_n862), .B2(new_n816), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT57), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n897), .A2(new_n898), .A3(new_n420), .ZN(new_n899));
  OAI21_X1  g698(.A(KEYINPUT57), .B1(new_n828), .B2(new_n363), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n870), .A2(new_n690), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT123), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT123), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n899), .A2(new_n905), .A3(new_n900), .A4(new_n902), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n906), .A2(G148gat), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n893), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n871), .B1(new_n873), .B2(new_n874), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(new_n690), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n910), .A2(KEYINPUT59), .A3(new_n221), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n892), .B1(new_n908), .B2(new_n911), .ZN(G1345gat));
  OAI21_X1  g711(.A(G155gat), .B1(new_n909), .B2(new_n688), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n881), .A2(new_n213), .A3(new_n615), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1346gat));
  NAND2_X1  g714(.A1(new_n754), .A2(G162gat), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n881), .A2(new_n754), .ZN(new_n917));
  OAI22_X1  g716(.A1(new_n909), .A2(new_n916), .B1(new_n917), .B2(G162gat), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT124), .ZN(G1347gat));
  NAND2_X1  g718(.A1(new_n697), .A2(new_n371), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT125), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n921), .A2(new_n737), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n831), .A2(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(G169gat), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n923), .A2(new_n924), .A3(new_n529), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n828), .A2(new_n670), .ZN(new_n926));
  AND4_X1   g725(.A1(new_n697), .A2(new_n926), .A3(new_n363), .A4(new_n430), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n689), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n925), .B1(new_n928), .B2(new_n924), .ZN(G1348gat));
  INV_X1    g728(.A(G176gat), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n927), .A2(new_n930), .A3(new_n648), .ZN(new_n931));
  OAI21_X1  g730(.A(G176gat), .B1(new_n923), .B2(new_n690), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1349gat));
  NAND3_X1  g732(.A1(new_n927), .A2(new_n292), .A3(new_n615), .ZN(new_n934));
  OAI21_X1  g733(.A(G183gat), .B1(new_n923), .B2(new_n688), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g736(.A(G190gat), .B1(new_n923), .B2(new_n584), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT61), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n927), .A2(new_n275), .A3(new_n754), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(G1351gat));
  NOR2_X1   g740(.A1(new_n880), .A2(new_n418), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n942), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n943), .A2(G197gat), .A3(new_n529), .ZN(new_n944));
  INV_X1    g743(.A(new_n658), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n945), .A2(new_n921), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n899), .A2(new_n689), .A3(new_n900), .A4(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n944), .B1(new_n947), .B2(G197gat), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT126), .ZN(G1352gat));
  INV_X1    g748(.A(new_n943), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n950), .A2(new_n312), .A3(new_n648), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT62), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n901), .A2(new_n946), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n312), .B1(new_n953), .B2(new_n648), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n952), .A2(new_n954), .ZN(G1353gat));
  NOR3_X1   g754(.A1(new_n943), .A2(G211gat), .A3(new_n688), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n899), .A2(new_n615), .A3(new_n900), .A4(new_n946), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT63), .B1(new_n957), .B2(G211gat), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT127), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n958), .A2(new_n959), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n957), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(G1354gat));
  NAND3_X1  g762(.A1(new_n950), .A2(new_n571), .A3(new_n754), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n953), .A2(new_n754), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n965), .B2(new_n571), .ZN(G1355gat));
endmodule


