//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 1 1 1 0 1 0 1 0 1 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 1 0 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0007(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n211));
  NAND4_X1  g0011(.A1(new_n208), .A2(new_n209), .A3(new_n210), .A4(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G1), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n212), .A2(new_n216), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT65), .Z(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT66), .Z(new_n221));
  NOR2_X1   g0021(.A1(new_n216), .A2(G13), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT0), .Z(new_n224));
  INV_X1    g0024(.A(new_n201), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G50), .ZN(new_n226));
  NAND3_X1  g0026(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NOR4_X1   g0028(.A1(new_n219), .A2(new_n221), .A3(new_n224), .A4(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G226), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT67), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n234), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G68), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n202), .ZN(new_n241));
  INV_X1    g0041(.A(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  INV_X1    g0047(.A(KEYINPUT3), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G222), .ZN(new_n254));
  INV_X1    g0054(.A(G223), .ZN(new_n255));
  OAI211_X1 g0055(.A(new_n252), .B(new_n254), .C1(new_n255), .C2(new_n253), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G1), .A2(G13), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n257), .B1(G33), .B2(G41), .ZN(new_n258));
  OAI211_X1 g0058(.A(new_n256), .B(new_n258), .C1(G77), .C2(new_n252), .ZN(new_n259));
  INV_X1    g0059(.A(G45), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT68), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT68), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G45), .ZN(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n261), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(new_n213), .A3(G274), .ZN(new_n266));
  INV_X1    g0066(.A(G226), .ZN(new_n267));
  OAI211_X1 g0067(.A(G1), .B(G13), .C1(new_n249), .C2(new_n264), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n213), .B1(G41), .B2(G45), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n259), .B(new_n266), .C1(new_n267), .C2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G169), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n273), .B1(G179), .B2(new_n271), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n213), .A2(G13), .A3(G20), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n202), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n257), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n213), .A2(G20), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n277), .B1(new_n282), .B2(new_n202), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT69), .ZN(new_n284));
  NOR3_X1   g0084(.A1(new_n284), .A2(new_n242), .A3(KEYINPUT8), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n285), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n287), .A2(new_n214), .A3(G33), .ZN(new_n288));
  INV_X1    g0088(.A(G150), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  OAI221_X1 g0091(.A(new_n288), .B1(new_n289), .B2(new_n291), .C1(new_n214), .C2(new_n204), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n283), .B1(new_n292), .B2(new_n279), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n274), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G190), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n271), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(G200), .B2(new_n271), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT9), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n293), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n293), .A2(new_n298), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n297), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT10), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT10), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n303), .B(new_n297), .C1(new_n299), .C2(new_n300), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n294), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT70), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n275), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n275), .A2(new_n306), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(KEYINPUT12), .B1(new_n310), .B2(G68), .ZN(new_n311));
  INV_X1    g0111(.A(G13), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n312), .A2(G1), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT12), .ZN(new_n314));
  INV_X1    g0114(.A(G68), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n313), .A2(new_n314), .A3(G20), .A4(new_n315), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n316), .B(KEYINPUT73), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n311), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(KEYINPUT70), .B1(new_n313), .B2(G20), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n319), .A2(new_n307), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(new_n279), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n315), .B1(new_n213), .B2(G20), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT74), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT74), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n318), .A2(new_n326), .A3(new_n323), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n315), .A2(G20), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n214), .A2(G33), .ZN(new_n329));
  OAI221_X1 g0129(.A(new_n328), .B1(new_n329), .B2(new_n205), .C1(new_n291), .C2(new_n202), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n279), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n331), .B(KEYINPUT11), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n325), .A2(new_n327), .A3(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT14), .ZN(new_n334));
  INV_X1    g0134(.A(G238), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n266), .B1(new_n335), .B2(new_n270), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n267), .A2(G1698), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n252), .A2(new_n337), .B1(G33), .B2(G97), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT72), .ZN(new_n339));
  AND2_X1   g0139(.A1(G232), .A2(G1698), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n339), .B1(new_n252), .B2(new_n340), .ZN(new_n341));
  AND2_X1   g0141(.A1(KEYINPUT3), .A2(G33), .ZN(new_n342));
  NOR2_X1   g0142(.A1(KEYINPUT3), .A2(G33), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n339), .B(new_n340), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n338), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n336), .B1(new_n346), .B2(new_n258), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT13), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n340), .B1(new_n342), .B2(new_n343), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT72), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n344), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n268), .B1(new_n352), .B2(new_n338), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n353), .A2(KEYINPUT13), .A3(new_n336), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n334), .B(G169), .C1(new_n349), .C2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n347), .A2(new_n348), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT13), .B1(new_n353), .B2(new_n336), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n356), .A2(G179), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n356), .A2(new_n357), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n334), .B1(new_n360), .B2(G169), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n333), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  AND3_X1   g0162(.A1(new_n325), .A2(new_n327), .A3(new_n332), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n360), .A2(G200), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n363), .B(new_n364), .C1(new_n295), .C2(new_n360), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n321), .A2(G77), .A3(new_n281), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n320), .A2(new_n205), .ZN(new_n367));
  NAND2_X1  g0167(.A1(G20), .A2(G77), .ZN(new_n368));
  XNOR2_X1  g0168(.A(KEYINPUT15), .B(G87), .ZN(new_n369));
  OAI221_X1 g0169(.A(new_n368), .B1(new_n286), .B2(new_n291), .C1(new_n329), .C2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n279), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n366), .A2(new_n367), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT71), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT71), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n366), .A2(new_n374), .A3(new_n367), .A4(new_n371), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G238), .A2(G1698), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n252), .B(new_n377), .C1(new_n233), .C2(G1698), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n378), .B(new_n258), .C1(G107), .C2(new_n252), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n268), .A2(G244), .A3(new_n269), .ZN(new_n380));
  AND2_X1   g0180(.A1(new_n266), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(G169), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  AND2_X1   g0182(.A1(new_n379), .A2(new_n381), .ZN(new_n383));
  INV_X1    g0183(.A(G179), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n376), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n383), .A2(G190), .ZN(new_n388));
  INV_X1    g0188(.A(G200), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n388), .B1(new_n389), .B2(new_n383), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n376), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n305), .A2(new_n362), .A3(new_n365), .A4(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n287), .A2(new_n275), .ZN(new_n394));
  INV_X1    g0194(.A(new_n282), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n394), .B1(new_n287), .B2(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n242), .A2(new_n315), .ZN(new_n397));
  OAI21_X1  g0197(.A(G20), .B1(new_n397), .B2(new_n201), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n290), .A2(G159), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n250), .A2(new_n214), .A3(new_n251), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT7), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT75), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n250), .A2(KEYINPUT7), .A3(new_n214), .A4(new_n251), .ZN(new_n406));
  AND3_X1   g0206(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(G68), .B1(new_n404), .B2(new_n405), .ZN(new_n408));
  OAI211_X1 g0208(.A(KEYINPUT16), .B(new_n401), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n279), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT76), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n404), .A2(new_n411), .A3(new_n406), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n402), .A2(KEYINPUT76), .A3(new_n403), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(G68), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(KEYINPUT16), .B1(new_n414), .B2(new_n401), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n396), .B1(new_n410), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n255), .A2(new_n253), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n267), .A2(G1698), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n417), .B(new_n418), .C1(new_n342), .C2(new_n343), .ZN(new_n419));
  NAND2_X1  g0219(.A1(G33), .A2(G87), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT77), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT77), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n419), .A2(new_n423), .A3(new_n420), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n422), .A2(new_n424), .A3(new_n258), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n268), .A2(G232), .A3(new_n269), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n266), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n425), .A2(new_n295), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n268), .B1(new_n421), .B2(KEYINPUT77), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n427), .B1(new_n430), .B2(new_n424), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n429), .B1(G200), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT17), .ZN(new_n434));
  AND2_X1   g0234(.A1(new_n434), .A2(KEYINPUT79), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n434), .A2(KEYINPUT79), .ZN(new_n436));
  OAI22_X1  g0236(.A1(new_n416), .A2(new_n433), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n396), .ZN(new_n438));
  INV_X1    g0238(.A(new_n415), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n342), .A2(new_n343), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT7), .B1(new_n440), .B2(new_n214), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n315), .B1(new_n441), .B2(KEYINPUT75), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n400), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n280), .B1(new_n444), .B2(KEYINPUT16), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n438), .B1(new_n439), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n436), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n446), .A2(new_n432), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n437), .A2(new_n448), .ZN(new_n449));
  AOI211_X1 g0249(.A(new_n384), .B(new_n427), .C1(new_n430), .C2(new_n424), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n272), .B1(new_n425), .B2(new_n428), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT78), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  AND3_X1   g0253(.A1(new_n419), .A2(new_n423), .A3(new_n420), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n423), .B1(new_n419), .B2(new_n420), .ZN(new_n455));
  NOR3_X1   g0255(.A1(new_n454), .A2(new_n455), .A3(new_n268), .ZN(new_n456));
  OAI21_X1  g0256(.A(G169), .B1(new_n456), .B2(new_n427), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n425), .A2(G179), .A3(new_n428), .ZN(new_n458));
  AOI21_X1  g0258(.A(KEYINPUT78), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  OAI211_X1 g0259(.A(KEYINPUT18), .B(new_n416), .C1(new_n453), .C2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n452), .B1(new_n450), .B2(new_n451), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n457), .A2(KEYINPUT78), .A3(new_n458), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT18), .B1(new_n464), .B2(new_n416), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n449), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n260), .A2(G1), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n264), .A2(KEYINPUT5), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT5), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G41), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n467), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n471), .A2(G257), .A3(new_n268), .ZN(new_n472));
  XNOR2_X1  g0272(.A(KEYINPUT5), .B(G41), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n473), .A2(new_n268), .A3(G274), .A4(new_n467), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(G250), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n476), .B1(new_n250), .B2(new_n251), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT4), .ZN(new_n478));
  OAI21_X1  g0278(.A(G1698), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G283), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(G244), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n482), .B1(new_n250), .B2(new_n251), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n478), .A2(G1698), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n478), .B1(new_n440), .B2(new_n482), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n479), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n475), .B1(new_n487), .B2(new_n258), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n295), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n489), .B1(G200), .B2(new_n488), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n412), .A2(G107), .A3(new_n413), .ZN(new_n491));
  INV_X1    g0291(.A(G107), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n492), .A2(KEYINPUT6), .A3(G97), .ZN(new_n493));
  INV_X1    g0293(.A(G97), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n494), .A2(new_n492), .ZN(new_n495));
  NOR2_X1   g0295(.A1(G97), .A2(G107), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n493), .B1(new_n497), .B2(KEYINPUT6), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n498), .A2(G20), .B1(G77), .B2(new_n290), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n491), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n279), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n275), .A2(G97), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n280), .B(new_n275), .C1(G1), .C2(new_n249), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n502), .B1(new_n504), .B2(G97), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n501), .A2(KEYINPUT80), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT80), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n280), .B1(new_n491), .B2(new_n499), .ZN(new_n508));
  INV_X1    g0308(.A(new_n505), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n490), .A2(new_n506), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(G87), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(new_n494), .A3(new_n492), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G97), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n214), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n513), .A2(new_n515), .A3(KEYINPUT19), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n214), .B(G68), .C1(new_n342), .C2(new_n343), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT19), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n329), .B2(new_n494), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n516), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n279), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n320), .A2(new_n369), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT82), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT82), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n525), .A2(new_n526), .B1(G87), .B2(new_n504), .ZN(new_n527));
  INV_X1    g0327(.A(G274), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n467), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n476), .B1(new_n260), .B2(G1), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n529), .A2(new_n268), .A3(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(G238), .A2(G1698), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(new_n482), .B2(G1698), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n533), .A2(new_n252), .B1(G33), .B2(G116), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n531), .B1(new_n534), .B2(new_n268), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n535), .A2(new_n295), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n536), .B1(G200), .B2(new_n535), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT82), .ZN(new_n538));
  AOI21_X1  g0338(.A(KEYINPUT82), .B1(new_n521), .B2(new_n522), .ZN(new_n539));
  OAI22_X1  g0339(.A1(new_n538), .A2(new_n539), .B1(new_n369), .B2(new_n503), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n535), .A2(new_n272), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n384), .B(new_n531), .C1(new_n534), .C2(new_n268), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n527), .A2(new_n537), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  AOI211_X1 g0344(.A(new_n384), .B(new_n475), .C1(new_n487), .C2(new_n258), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n484), .B(G244), .C1(new_n343), .C2(new_n342), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n546), .B(new_n480), .C1(new_n483), .C2(KEYINPUT4), .ZN(new_n547));
  OAI21_X1  g0347(.A(G250), .B1(new_n342), .B2(new_n343), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n253), .B1(new_n548), .B2(KEYINPUT4), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n258), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n475), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n272), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI22_X1  g0352(.A1(new_n545), .A2(new_n552), .B1(new_n508), .B2(new_n509), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n553), .A2(KEYINPUT81), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT81), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n501), .A2(new_n505), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n550), .A2(new_n551), .A3(G179), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(new_n488), .B2(new_n272), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n555), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n511), .B(new_n544), .C1(new_n554), .C2(new_n559), .ZN(new_n560));
  XNOR2_X1  g0360(.A(KEYINPUT84), .B(KEYINPUT24), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n214), .B(G87), .C1(new_n342), .C2(new_n343), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT22), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT22), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n252), .A2(new_n564), .A3(new_n214), .A4(G87), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(KEYINPUT85), .B(KEYINPUT23), .C1(new_n214), .C2(G107), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n214), .A2(G33), .A3(G116), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n492), .A2(G20), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n567), .B(new_n568), .C1(KEYINPUT23), .C2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(KEYINPUT85), .B1(new_n569), .B2(KEYINPUT23), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n561), .B1(new_n566), .B2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n566), .A2(new_n572), .A3(new_n561), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n280), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n276), .A2(new_n492), .ZN(new_n577));
  OR2_X1    g0377(.A1(new_n577), .A2(KEYINPUT25), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(KEYINPUT25), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n578), .B(new_n579), .C1(new_n492), .C2(new_n503), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n471), .A2(G264), .A3(new_n268), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n474), .ZN(new_n582));
  AND2_X1   g0382(.A1(G257), .A2(G1698), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n252), .A2(new_n583), .B1(G33), .B2(G294), .ZN(new_n584));
  OAI211_X1 g0384(.A(G250), .B(new_n253), .C1(new_n342), .C2(new_n343), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n268), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT86), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n582), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n583), .B1(new_n342), .B2(new_n343), .ZN(new_n589));
  NAND2_X1  g0389(.A1(G33), .A2(G294), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n585), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n258), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT86), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n272), .B1(new_n588), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(new_n474), .A3(new_n581), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n595), .A2(new_n384), .ZN(new_n596));
  OAI22_X1  g0396(.A1(new_n576), .A2(new_n580), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(G116), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n308), .A2(new_n598), .A3(new_n309), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n598), .B1(new_n213), .B2(G33), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n280), .B(new_n600), .C1(new_n319), .C2(new_n307), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n278), .A2(new_n257), .B1(G20), .B2(new_n598), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n480), .B(new_n214), .C1(G33), .C2(new_n494), .ZN(new_n603));
  AOI21_X1  g0403(.A(KEYINPUT20), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n602), .A2(KEYINPUT20), .A3(new_n603), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n599), .B(new_n601), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n253), .A2(G257), .ZN(new_n607));
  NAND2_X1  g0407(.A1(G264), .A2(G1698), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n607), .B(new_n608), .C1(new_n342), .C2(new_n343), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n609), .B(new_n258), .C1(G303), .C2(new_n252), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n471), .A2(G270), .A3(new_n268), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(new_n474), .A3(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n606), .A2(KEYINPUT21), .A3(G169), .A4(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n612), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n614), .A2(new_n606), .A3(G179), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(G303), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n268), .B1(new_n440), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n258), .A2(new_n528), .ZN(new_n619));
  INV_X1    g0419(.A(new_n471), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n618), .A2(new_n609), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n272), .B1(new_n621), .B2(new_n611), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT21), .B1(new_n622), .B2(new_n606), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n616), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n591), .A2(new_n587), .A3(new_n258), .ZN(new_n625));
  INV_X1    g0425(.A(new_n582), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n593), .A2(new_n295), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n595), .A2(new_n389), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n575), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n279), .B1(new_n630), .B2(new_n573), .ZN(new_n631));
  INV_X1    g0431(.A(new_n580), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n629), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n389), .B1(new_n621), .B2(new_n611), .ZN(new_n634));
  OAI21_X1  g0434(.A(KEYINPUT83), .B1(new_n634), .B2(new_n606), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n612), .A2(G200), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT83), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n605), .A2(new_n604), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n599), .A2(new_n601), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n636), .A2(new_n637), .A3(new_n638), .A4(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n614), .A2(G190), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n635), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n597), .A2(new_n624), .A3(new_n633), .A4(new_n642), .ZN(new_n643));
  NOR4_X1   g0443(.A1(new_n393), .A2(new_n466), .A3(new_n560), .A4(new_n643), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n644), .B(KEYINPUT87), .ZN(G372));
  INV_X1    g0445(.A(new_n449), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n365), .A2(new_n387), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n646), .B1(new_n647), .B2(new_n362), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT18), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n457), .A2(new_n458), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n416), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n649), .B1(new_n416), .B2(new_n650), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n648), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n655), .B1(new_n302), .B2(new_n304), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n656), .A2(new_n294), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n393), .A2(new_n466), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n540), .A2(new_n543), .ZN(new_n659));
  INV_X1    g0459(.A(new_n624), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n588), .A2(new_n593), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(G169), .ZN(new_n662));
  INV_X1    g0462(.A(new_n596), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n662), .A2(new_n663), .B1(new_n631), .B2(new_n632), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n633), .B1(new_n660), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n659), .B1(new_n560), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n553), .A2(KEYINPUT81), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n556), .A2(new_n558), .A3(new_n555), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n544), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(KEYINPUT26), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT88), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(new_n545), .B2(new_n552), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n557), .B(KEYINPUT88), .C1(new_n488), .C2(new_n272), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n506), .A2(new_n510), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n544), .A2(new_n674), .A3(new_n675), .A4(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n670), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n658), .B1(new_n666), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n657), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT89), .ZN(G369));
  NAND2_X1  g0481(.A1(new_n313), .A2(new_n214), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G213), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT90), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n687), .A2(G343), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(G343), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n664), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT91), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n692), .B1(new_n576), .B2(new_n580), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n597), .A2(new_n695), .A3(new_n633), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n624), .A2(new_n692), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n697), .A2(new_n698), .B1(new_n664), .B2(new_n691), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n692), .A2(new_n606), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n624), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n624), .A2(new_n642), .A3(new_n700), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G330), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n697), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n699), .A2(new_n706), .ZN(G399));
  OR2_X1    g0507(.A1(new_n513), .A2(G116), .ZN(new_n708));
  XOR2_X1   g0508(.A(new_n708), .B(KEYINPUT92), .Z(new_n709));
  NAND2_X1  g0509(.A1(new_n222), .A2(new_n264), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n709), .A2(new_n213), .A3(new_n711), .ZN(new_n712));
  OAI22_X1  g0512(.A1(new_n712), .A2(KEYINPUT93), .B1(new_n226), .B2(new_n710), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n713), .B1(KEYINPUT93), .B2(new_n712), .ZN(new_n714));
  XOR2_X1   g0514(.A(new_n714), .B(KEYINPUT28), .Z(new_n715));
  OAI21_X1  g0515(.A(new_n691), .B1(new_n666), .B2(new_n678), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT29), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(KEYINPUT94), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT94), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n716), .A2(new_n720), .A3(new_n717), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n544), .A2(new_n674), .A3(new_n676), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT26), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n544), .A2(new_n667), .A3(new_n675), .A4(new_n668), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OAI211_X1 g0525(.A(KEYINPUT29), .B(new_n691), .C1(new_n666), .C2(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n719), .A2(new_n721), .A3(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(G330), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n506), .A2(new_n510), .ZN(new_n729));
  AOI22_X1  g0529(.A1(new_n729), .A2(new_n490), .B1(new_n667), .B2(new_n668), .ZN(new_n730));
  AND4_X1   g0530(.A1(new_n597), .A2(new_n624), .A3(new_n633), .A4(new_n642), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n730), .A2(new_n544), .A3(new_n731), .A4(new_n691), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT30), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n620), .A2(new_n258), .ZN(new_n734));
  AOI22_X1  g0534(.A1(new_n734), .A2(G264), .B1(new_n591), .B2(new_n258), .ZN(new_n735));
  INV_X1    g0535(.A(new_n531), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n533), .A2(new_n252), .ZN(new_n737));
  NAND2_X1  g0537(.A1(G33), .A2(G116), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n736), .B1(new_n739), .B2(new_n258), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n614), .A2(new_n735), .A3(G179), .A4(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n488), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n733), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n614), .A2(new_n740), .A3(G179), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(new_n742), .A3(new_n595), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n735), .A2(new_n740), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n612), .A2(new_n384), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n746), .A2(KEYINPUT30), .A3(new_n488), .A4(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n743), .A2(new_n745), .A3(new_n748), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n749), .A2(KEYINPUT31), .A3(new_n692), .ZN(new_n750));
  AOI21_X1  g0550(.A(KEYINPUT31), .B1(new_n749), .B2(new_n692), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n728), .B1(new_n732), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n727), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n715), .B1(new_n756), .B2(G1), .ZN(G364));
  NOR2_X1   g0557(.A1(new_n312), .A2(G20), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n213), .B1(new_n758), .B2(G45), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n711), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n705), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n762), .B1(G330), .B2(new_n703), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n222), .A2(new_n252), .ZN(new_n764));
  INV_X1    g0564(.A(G355), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n764), .A2(new_n765), .B1(G116), .B2(new_n222), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n243), .A2(G45), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n222), .A2(new_n440), .ZN(new_n768));
  INV_X1    g0568(.A(new_n226), .ZN(new_n769));
  AND2_X1   g0569(.A1(new_n261), .A2(new_n263), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n766), .B1(new_n767), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G13), .A2(G33), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n257), .B1(G20), .B2(new_n272), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n761), .B1(new_n772), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT95), .ZN(new_n780));
  AND2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n295), .ZN(new_n783));
  AND2_X1   g0583(.A1(new_n783), .A2(G326), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n214), .A2(new_n295), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n384), .A2(G200), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n252), .B(new_n784), .C1(G322), .C2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n214), .A2(G190), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n389), .A2(G179), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(G311), .A2(new_n792), .B1(new_n795), .B2(G283), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n785), .A2(new_n793), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(G179), .A2(G200), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n790), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(G303), .A2(new_n798), .B1(new_n801), .B2(G329), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n214), .B1(new_n799), .B2(G190), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n782), .A2(G190), .ZN(new_n805));
  XNOR2_X1  g0605(.A(KEYINPUT33), .B(G317), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n804), .A2(G294), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n789), .A2(new_n796), .A3(new_n802), .A4(new_n807), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n787), .A2(new_n242), .B1(new_n791), .B2(new_n205), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT96), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n252), .B1(new_n794), .B2(new_n492), .C1(new_n512), .C2(new_n797), .ZN(new_n811));
  INV_X1    g0611(.A(new_n783), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n812), .A2(new_n202), .B1(new_n803), .B2(new_n494), .ZN(new_n813));
  OR3_X1    g0613(.A1(new_n810), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(G159), .ZN(new_n815));
  OR3_X1    g0615(.A1(new_n800), .A2(KEYINPUT32), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(KEYINPUT32), .B1(new_n800), .B2(new_n815), .ZN(new_n817));
  INV_X1    g0617(.A(new_n805), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n816), .B(new_n817), .C1(new_n315), .C2(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n808), .B1(new_n814), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n781), .B1(new_n776), .B2(new_n820), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n775), .B(KEYINPUT97), .Z(new_n822));
  OAI221_X1 g0622(.A(new_n821), .B1(new_n780), .B2(new_n779), .C1(new_n703), .C2(new_n822), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n763), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(G396));
  AOI21_X1  g0625(.A(new_n691), .B1(new_n373), .B2(new_n375), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n386), .B1(new_n391), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n376), .A2(new_n385), .A3(new_n691), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n716), .A2(new_n829), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n827), .A2(new_n828), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n691), .B(new_n831), .C1(new_n666), .C2(new_n678), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n761), .B1(new_n833), .B2(new_n754), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n754), .B2(new_n833), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n776), .A2(new_n773), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n760), .B(new_n711), .C1(new_n205), .C2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n776), .ZN(new_n838));
  AOI22_X1  g0638(.A1(G143), .A2(new_n788), .B1(new_n792), .B2(G159), .ZN(new_n839));
  INV_X1    g0639(.A(G137), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n839), .B1(new_n812), .B2(new_n840), .C1(new_n289), .C2(new_n818), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT34), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n252), .B1(new_n794), .B2(new_n315), .ZN(new_n843));
  INV_X1    g0643(.A(G132), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n797), .A2(new_n202), .B1(new_n800), .B2(new_n844), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n843), .B(new_n845), .C1(G58), .C2(new_n804), .ZN(new_n846));
  INV_X1    g0646(.A(G283), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n440), .B1(new_n794), .B2(new_n512), .C1(new_n818), .C2(new_n847), .ZN(new_n848));
  AOI22_X1  g0648(.A1(G107), .A2(new_n798), .B1(new_n792), .B2(G116), .ZN(new_n849));
  INV_X1    g0649(.A(G311), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n849), .B1(new_n850), .B2(new_n800), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n848), .B(new_n851), .C1(G303), .C2(new_n783), .ZN(new_n852));
  INV_X1    g0652(.A(G294), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n787), .A2(new_n853), .B1(new_n803), .B2(new_n494), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT98), .Z(new_n855));
  AOI22_X1  g0655(.A1(new_n842), .A2(new_n846), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n837), .B1(new_n838), .B2(new_n856), .C1(new_n831), .C2(new_n774), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n835), .A2(new_n857), .ZN(G384));
  NAND2_X1  g0658(.A1(new_n498), .A2(KEYINPUT35), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n227), .A2(new_n598), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n498), .B2(KEYINPUT35), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT99), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n859), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n862), .B2(new_n861), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT36), .ZN(new_n865));
  OR3_X1    g0665(.A1(new_n226), .A2(new_n205), .A3(new_n397), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n202), .A2(G68), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n213), .B(G13), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT101), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n333), .A2(new_n692), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n362), .A2(new_n365), .A3(new_n871), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n333), .B(new_n692), .C1(new_n359), .C2(new_n361), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  XOR2_X1   g0675(.A(new_n828), .B(KEYINPUT100), .Z(new_n876));
  AOI21_X1  g0676(.A(new_n875), .B1(new_n832), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT38), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n444), .A2(KEYINPUT16), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n396), .B1(new_n410), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n686), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n416), .B1(new_n453), .B2(new_n459), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n649), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n460), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n881), .B1(new_n884), .B2(new_n449), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n880), .A2(new_n650), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n432), .B(new_n396), .C1(new_n415), .C2(new_n410), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n881), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n416), .B1(new_n464), .B2(new_n686), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT37), .B1(new_n446), .B2(new_n432), .ZN(new_n890));
  AOI22_X1  g0690(.A1(KEYINPUT37), .A2(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n878), .B1(new_n885), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n881), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n466), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n888), .A2(KEYINPUT37), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n889), .A2(new_n890), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n894), .A2(KEYINPUT38), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n892), .A2(new_n898), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n877), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n653), .A2(new_n686), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n870), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n885), .A2(new_n878), .A3(new_n891), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT38), .B1(new_n894), .B2(new_n897), .ZN(new_n904));
  OAI21_X1  g0704(.A(KEYINPUT39), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT39), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n416), .A2(new_n686), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n653), .B2(new_n449), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n416), .A2(new_n650), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(new_n907), .A3(new_n887), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(KEYINPUT37), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT102), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n911), .A2(new_n912), .B1(new_n890), .B2(new_n889), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n910), .A2(KEYINPUT102), .A3(KEYINPUT37), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n908), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n906), .B(new_n898), .C1(new_n915), .C2(KEYINPUT38), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n905), .A2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n362), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n691), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n901), .B1(new_n877), .B2(new_n899), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT101), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n902), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n719), .A2(new_n658), .A3(new_n726), .A4(new_n721), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n657), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n924), .B(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT40), .ZN(new_n928));
  INV_X1    g0728(.A(new_n899), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n829), .B1(new_n872), .B2(new_n873), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n732), .A2(new_n752), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n928), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n930), .A2(new_n931), .A3(KEYINPUT40), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n911), .A2(new_n912), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n935), .A2(new_n896), .A3(new_n914), .ZN(new_n936));
  INV_X1    g0736(.A(new_n908), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT38), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n934), .B1(new_n938), .B2(new_n903), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n933), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n658), .A2(new_n931), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n942), .A2(G330), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n927), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n213), .B2(new_n758), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n927), .A2(new_n944), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n869), .B1(new_n946), .B2(new_n947), .ZN(G367));
  NAND2_X1  g0748(.A1(new_n697), .A2(new_n698), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n730), .B1(new_n729), .B2(new_n691), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n674), .A2(new_n676), .A3(new_n692), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n949), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT42), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n953), .A2(new_n597), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n554), .A2(new_n559), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n691), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n527), .A2(new_n691), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n961), .A2(new_n659), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(new_n544), .B2(new_n961), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT43), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n963), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n959), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n955), .A2(new_n964), .A3(new_n963), .A4(new_n958), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n706), .A2(new_n953), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n970), .B(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n710), .B(KEYINPUT41), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT45), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT103), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n699), .A2(new_n975), .A3(new_n952), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n975), .B1(new_n699), .B2(new_n952), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n974), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n978), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n980), .A2(KEYINPUT45), .A3(new_n976), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT44), .ZN(new_n982));
  INV_X1    g0782(.A(new_n699), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n982), .B1(new_n983), .B2(new_n953), .ZN(new_n984));
  NOR3_X1   g0784(.A1(new_n699), .A2(KEYINPUT44), .A3(new_n952), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n979), .A2(new_n981), .A3(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n706), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(KEYINPUT104), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n697), .A2(new_n698), .ZN(new_n992));
  AND3_X1   g0792(.A1(new_n992), .A2(new_n705), .A3(new_n949), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n705), .B1(new_n992), .B2(new_n949), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n756), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n979), .A2(new_n981), .A3(new_n986), .A4(new_n989), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n991), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n973), .B1(new_n999), .B2(new_n756), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n972), .B1(new_n1000), .B2(new_n760), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n237), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n777), .B1(new_n222), .B2(new_n369), .C1(new_n1002), .C2(new_n768), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n761), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT105), .Z(new_n1005));
  NOR2_X1   g0805(.A1(new_n803), .A2(new_n315), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1007), .B(new_n252), .C1(new_n289), .C2(new_n787), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n794), .A2(new_n205), .B1(new_n800), .B2(new_n840), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n797), .A2(new_n242), .B1(new_n791), .B2(new_n202), .ZN(new_n1010));
  INV_X1    g0810(.A(G143), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n818), .A2(new_n815), .B1(new_n812), .B2(new_n1011), .ZN(new_n1012));
  NOR4_X1   g0812(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .A4(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(KEYINPUT46), .B1(new_n798), .B2(G116), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n798), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n812), .B2(new_n850), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n1014), .B(new_n1016), .C1(G107), .C2(new_n804), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n787), .A2(new_n617), .B1(new_n791), .B2(new_n847), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n440), .B1(new_n794), .B2(new_n494), .C1(new_n818), .C2(new_n853), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n1018), .B(new_n1019), .C1(G317), .C2(new_n801), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1013), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g0821(.A(KEYINPUT106), .B(KEYINPUT47), .Z(new_n1022));
  NOR2_X1   g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n776), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1005), .B1(new_n1023), .B2(new_n1025), .C1(new_n966), .C2(new_n822), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1001), .A2(new_n1026), .ZN(G387));
  OAI21_X1  g0827(.A(KEYINPUT111), .B1(new_n997), .B2(new_n710), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT112), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n756), .B2(new_n995), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT111), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n996), .A2(new_n1031), .A3(new_n711), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n755), .B(KEYINPUT112), .C1(new_n993), .C2(new_n994), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1028), .A2(new_n1030), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n697), .A2(new_n822), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n709), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n1036), .A2(new_n764), .B1(G107), .B2(new_n222), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT107), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n770), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n234), .A2(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  NOR3_X1   g0842(.A1(new_n1042), .A2(G50), .A3(new_n286), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n286), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1041), .B1(new_n1044), .B2(new_n202), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n260), .B1(new_n315), .B2(new_n205), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n1043), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n768), .B1(new_n1036), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1038), .B1(new_n1040), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n761), .B1(new_n1049), .B2(new_n778), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n803), .A2(new_n369), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n440), .B(new_n1051), .C1(G97), .C2(new_n795), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n783), .A2(G159), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n287), .A2(new_n805), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n797), .A2(new_n205), .B1(new_n791), .B2(new_n315), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n787), .A2(new_n202), .B1(new_n800), .B2(new_n289), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .A4(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n252), .B1(new_n801), .B2(G326), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n797), .A2(new_n853), .B1(new_n803), .B2(new_n847), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G317), .A2(new_n788), .B1(new_n792), .B2(G303), .ZN(new_n1061));
  XOR2_X1   g0861(.A(KEYINPUT109), .B(G322), .Z(new_n1062));
  OAI221_X1 g0862(.A(new_n1061), .B1(new_n812), .B2(new_n1062), .C1(new_n850), .C2(new_n818), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT48), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1060), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n1064), .B2(new_n1063), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT49), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1059), .B1(new_n598), .B2(new_n794), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1058), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT110), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n838), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1050), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n995), .A2(new_n760), .B1(new_n1035), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1034), .A2(new_n1075), .ZN(G393));
  OR2_X1    g0876(.A1(new_n987), .A2(new_n988), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n987), .A2(new_n988), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n711), .B(new_n999), .C1(new_n1079), .C2(new_n997), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n953), .A2(new_n775), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n797), .A2(new_n315), .B1(new_n800), .B2(new_n1011), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT113), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n252), .B1(new_n512), .B2(new_n794), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n1083), .B2(new_n1082), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT114), .Z(new_n1086));
  AOI22_X1  g0886(.A1(new_n788), .A2(G159), .B1(G150), .B2(new_n783), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT51), .Z(new_n1088));
  AOI22_X1  g0888(.A1(new_n1044), .A2(new_n792), .B1(new_n804), .B2(G77), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1088), .B(new_n1089), .C1(new_n202), .C2(new_n818), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1086), .A2(new_n1090), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n788), .A2(G311), .B1(G317), .B2(new_n783), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT52), .Z(new_n1093));
  OR2_X1    g0893(.A1(new_n1062), .A2(new_n800), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(G283), .A2(new_n798), .B1(new_n792), .B2(G294), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n440), .B1(new_n794), .B2(new_n492), .C1(new_n818), .C2(new_n617), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(G116), .B2(new_n804), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .A4(new_n1097), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT115), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n776), .B1(new_n1091), .B2(new_n1099), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n777), .B1(new_n494), .B2(new_n222), .C1(new_n246), .C2(new_n768), .ZN(new_n1101));
  AND4_X1   g0901(.A1(new_n761), .A2(new_n1081), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n1079), .B2(new_n760), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1080), .A2(new_n1103), .ZN(G390));
  OAI211_X1 g0904(.A(new_n691), .B(new_n831), .C1(new_n666), .C2(new_n725), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n876), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n874), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n898), .B1(new_n915), .B2(KEYINPUT38), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1107), .A2(new_n919), .A3(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n877), .A2(new_n920), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1109), .B1(new_n917), .B2(new_n1110), .ZN(new_n1111));
  NOR3_X1   g0911(.A1(new_n560), .A2(new_n643), .A3(new_n692), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n749), .A2(new_n692), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT31), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n749), .A2(KEYINPUT31), .A3(new_n692), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  OAI211_X1 g0917(.A(G330), .B(new_n831), .C1(new_n1112), .C2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1118), .A2(new_n875), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1111), .A2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n905), .B(new_n916), .C1(new_n877), .C2(new_n920), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n753), .A2(new_n831), .A3(new_n874), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1121), .A2(new_n1122), .A3(new_n1109), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n905), .A2(new_n916), .A3(new_n773), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n836), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n761), .B1(new_n287), .B2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n797), .A2(new_n289), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT53), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(KEYINPUT54), .B(G143), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n792), .A2(new_n1132), .B1(new_n795), .B2(G50), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1130), .B(new_n1133), .C1(new_n844), .C2(new_n787), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n440), .B1(new_n801), .B2(G125), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(G128), .A2(new_n783), .B1(new_n805), .B2(G137), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1135), .B(new_n1136), .C1(new_n815), .C2(new_n803), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n440), .B1(new_n797), .B2(new_n512), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT116), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(G97), .A2(new_n792), .B1(new_n795), .B2(G68), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(G116), .A2(new_n788), .B1(new_n801), .B2(G294), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n805), .A2(G107), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n804), .A2(G77), .B1(G283), .B2(new_n783), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .A4(new_n1143), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n1134), .A2(new_n1137), .B1(new_n1139), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1128), .B1(new_n1145), .B2(new_n776), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1125), .A2(new_n760), .B1(new_n1126), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n832), .A2(new_n876), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n874), .B1(new_n753), .B2(new_n831), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1148), .B1(new_n1119), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1118), .A2(new_n875), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1151), .A2(new_n1122), .A3(new_n876), .A4(new_n1105), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n658), .A2(new_n753), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1153), .A2(new_n657), .A3(new_n925), .A4(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1124), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n925), .A2(new_n657), .A3(new_n1154), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1120), .A2(new_n1158), .A3(new_n1123), .A4(new_n1153), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1156), .A2(new_n711), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1147), .A2(new_n1160), .ZN(G378));
  AOI21_X1  g0961(.A(new_n932), .B1(new_n892), .B2(new_n898), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n939), .B(G330), .C1(KEYINPUT40), .C2(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  OR2_X1    g0965(.A1(new_n305), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n305), .A2(new_n1165), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n293), .A2(new_n685), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1166), .A2(new_n1169), .A3(new_n1167), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1163), .A2(new_n1174), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(KEYINPUT101), .A2(new_n922), .B1(new_n917), .B2(new_n920), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n933), .A2(new_n1173), .A3(G330), .A4(new_n939), .ZN(new_n1177));
  AND4_X1   g0977(.A1(new_n902), .A2(new_n1175), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n1177), .A2(new_n1175), .B1(new_n1176), .B2(new_n902), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1123), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1122), .B1(new_n1121), .B2(new_n1109), .ZN(new_n1182));
  NOR3_X1   g0982(.A1(new_n1181), .A2(new_n1155), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT119), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1157), .B(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(KEYINPUT120), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1157), .B(KEYINPUT119), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT120), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n1159), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1180), .B1(new_n1186), .B2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(KEYINPUT121), .B1(new_n1190), .B2(KEYINPUT57), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n710), .B1(new_n1190), .B2(KEYINPUT57), .ZN(new_n1192));
  OR2_X1    g0992(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1187), .A2(new_n1159), .A3(new_n1188), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1188), .B1(new_n1187), .B2(new_n1159), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1193), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT121), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT57), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1191), .A2(new_n1192), .A3(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n761), .B1(G50), .B2(new_n1127), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1173), .A2(new_n774), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n783), .A2(G125), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n289), .B2(new_n803), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(G128), .A2(new_n788), .B1(new_n798), .B2(new_n1132), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n840), .B2(new_n791), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1204), .B(new_n1206), .C1(G132), .C2(new_n805), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n249), .B(new_n264), .C1(new_n794), .C2(new_n815), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(G124), .B2(new_n801), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1209), .A2(new_n1210), .A3(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1007), .B1(new_n818), .B2(new_n494), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n787), .A2(new_n492), .B1(new_n800), .B2(new_n847), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n369), .A2(new_n791), .B1(new_n794), .B2(new_n242), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n264), .B(new_n440), .C1(new_n797), .C2(new_n205), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1215), .B(new_n1216), .C1(KEYINPUT117), .C2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(KEYINPUT117), .B2(new_n1217), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1214), .B(new_n1219), .C1(G116), .C2(new_n783), .ZN(new_n1220));
  OR2_X1    g1020(.A1(new_n1220), .A2(KEYINPUT58), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(KEYINPUT58), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n202), .B1(new_n342), .B2(G41), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1213), .A2(new_n1221), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1201), .B(new_n1202), .C1(new_n776), .C2(new_n1224), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1225), .B(KEYINPUT118), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n760), .B2(new_n1193), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1200), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT122), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1200), .A2(KEYINPUT122), .A3(new_n1227), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(G375));
  OAI22_X1  g1033(.A1(new_n812), .A2(new_n853), .B1(new_n791), .B2(new_n492), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(G116), .B2(new_n805), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1235), .B(KEYINPUT123), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(G97), .A2(new_n798), .B1(new_n801), .B2(G303), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n847), .B2(new_n787), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n440), .B1(new_n794), .B2(new_n205), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1238), .A2(new_n1051), .A3(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n797), .A2(new_n815), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n787), .A2(new_n840), .B1(new_n791), .B2(new_n289), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1241), .B(new_n1242), .C1(G128), .C2(new_n801), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n252), .B1(new_n794), .B2(new_n242), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n812), .A2(new_n844), .B1(new_n803), .B2(new_n202), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1244), .B(new_n1245), .C1(new_n805), .C2(new_n1132), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1236), .A2(new_n1240), .B1(new_n1243), .B2(new_n1246), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n761), .B1(G68), .B2(new_n1127), .C1(new_n1247), .C2(new_n838), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(new_n875), .B2(new_n773), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n1153), .B2(new_n760), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(KEYINPUT124), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1153), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n1157), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n973), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1253), .A2(new_n1254), .A3(new_n1155), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1251), .A2(new_n1255), .ZN(G381));
  INV_X1    g1056(.A(G378), .ZN(new_n1257));
  NOR4_X1   g1057(.A1(G387), .A2(G390), .A3(G384), .A4(G381), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1034), .A2(new_n824), .A3(new_n1075), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1232), .A2(new_n1257), .A3(new_n1258), .A4(new_n1260), .ZN(G407));
  NAND3_X1  g1061(.A1(new_n688), .A2(new_n689), .A3(G213), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1232), .A2(new_n1257), .A3(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(G407), .A2(G213), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(KEYINPUT125), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT125), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(G407), .A2(new_n1264), .A3(new_n1267), .A4(G213), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(G409));
  INV_X1    g1069(.A(KEYINPUT63), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1200), .A2(G378), .A3(new_n1227), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1254), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1180), .B1(new_n1272), .B2(new_n759), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1257), .B1(new_n1273), .B2(new_n1225), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1271), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1262), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT60), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1253), .A2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1252), .A2(new_n1157), .A3(KEYINPUT60), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1278), .A2(new_n711), .A3(new_n1155), .A4(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1280), .A2(new_n1251), .A3(G384), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(G384), .B1(new_n1280), .B2(new_n1251), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1270), .B1(new_n1276), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1263), .A2(G2897), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1284), .A2(new_n1287), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1284), .A2(new_n1287), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(KEYINPUT61), .B1(new_n1276), .B2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n824), .B1(new_n1034), .B2(new_n1075), .ZN(new_n1292));
  OAI211_X1 g1092(.A(G387), .B(KEYINPUT126), .C1(new_n1260), .C2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1292), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1294), .A2(new_n1001), .A3(new_n1026), .A4(new_n1259), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1293), .A2(G390), .A3(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(G390), .B1(new_n1293), .B2(new_n1295), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1263), .B1(new_n1271), .B2(new_n1274), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1299), .A2(KEYINPUT63), .A3(new_n1284), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1286), .A2(new_n1291), .A3(new_n1298), .A4(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT62), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1299), .A2(new_n1302), .A3(new_n1284), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT61), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1290), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1304), .B1(new_n1299), .B2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1302), .B1(new_n1299), .B2(new_n1284), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1303), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1301), .B1(new_n1308), .B2(new_n1298), .ZN(G405));
  INV_X1    g1109(.A(KEYINPUT127), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1310), .B1(new_n1232), .B2(G378), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1230), .A2(KEYINPUT127), .A3(new_n1257), .A4(new_n1231), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1311), .A2(new_n1271), .A3(new_n1312), .ZN(new_n1313));
  NOR3_X1   g1113(.A1(new_n1296), .A2(new_n1297), .A3(new_n1284), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(G387), .A2(KEYINPUT126), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1260), .A2(new_n1292), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1295), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(G390), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1293), .A2(G390), .A3(new_n1295), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1285), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  OR2_X1    g1121(.A1(new_n1314), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1313), .A2(new_n1322), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1314), .A2(new_n1321), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1324), .A2(new_n1271), .A3(new_n1312), .A4(new_n1311), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1323), .A2(new_n1325), .ZN(G402));
endmodule


