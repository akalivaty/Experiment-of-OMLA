//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 1 1 0 1 1 1 0 0 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  NOR3_X1   g003(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G148gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G141gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT73), .ZN(new_n210));
  OAI22_X1  g009(.A1(new_n205), .A2(new_n207), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G141gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G148gat), .ZN(new_n213));
  AND3_X1   g012(.A1(new_n209), .A2(new_n213), .A3(new_n210), .ZN(new_n214));
  AOI21_X1  g013(.A(KEYINPUT2), .B1(new_n209), .B2(new_n213), .ZN(new_n215));
  NOR2_X1   g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(new_n206), .ZN(new_n218));
  OAI22_X1  g017(.A1(new_n211), .A2(new_n214), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT22), .ZN(new_n220));
  INV_X1    g019(.A(G211gat), .ZN(new_n221));
  INV_X1    g020(.A(G218gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT71), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT71), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n225), .B(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n226));
  XNOR2_X1  g025(.A(G197gat), .B(G204gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n224), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G211gat), .B(G218gat), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n224), .A2(new_n229), .A3(new_n226), .A4(new_n227), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT29), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n219), .B1(new_n233), .B2(KEYINPUT3), .ZN(new_n234));
  AND3_X1   g033(.A1(new_n231), .A2(KEYINPUT72), .A3(new_n232), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT72), .B1(new_n231), .B2(new_n232), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT74), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n238), .B1(new_n219), .B2(KEYINPUT3), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT2), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n216), .A2(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n212), .A2(G148gat), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n241), .A2(new_n206), .B1(new_n242), .B2(KEYINPUT73), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n209), .A2(new_n213), .A3(new_n210), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n208), .A2(G141gat), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n240), .B1(new_n242), .B2(new_n245), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n207), .A2(new_n216), .ZN(new_n247));
  AOI22_X1  g046(.A1(new_n243), .A2(new_n244), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n248), .A2(KEYINPUT74), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT29), .B1(new_n239), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n234), .B1(new_n237), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(G228gat), .A2(G233gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n253), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n255), .B(new_n234), .C1(new_n237), .C2(new_n251), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT78), .B(G22gat), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n254), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n257), .B1(new_n254), .B2(new_n256), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n204), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n254), .A2(KEYINPUT79), .A3(new_n256), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT79), .B1(new_n254), .B2(new_n256), .ZN(new_n263));
  INV_X1    g062(.A(G22gat), .ZN(new_n264));
  NOR3_X1   g063(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n204), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n258), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n261), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G8gat), .B(G36gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(G64gat), .B(G92gat), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n270), .B(new_n271), .Z(new_n272));
  INV_X1    g071(.A(new_n237), .ZN(new_n273));
  NAND2_X1  g072(.A1(G226gat), .A2(G233gat), .ZN(new_n274));
  INV_X1    g073(.A(G169gat), .ZN(new_n275));
  INV_X1    g074(.A(G176gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278));
  NOR3_X1   g077(.A1(new_n277), .A2(KEYINPUT26), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G183gat), .A2(G190gat), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  AND2_X1   g080(.A1(new_n278), .A2(KEYINPUT26), .ZN(new_n282));
  NOR3_X1   g081(.A1(new_n279), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT27), .B(G183gat), .ZN(new_n285));
  INV_X1    g084(.A(G190gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(KEYINPUT28), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n289));
  INV_X1    g088(.A(G183gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT27), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT27), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G183gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n291), .A2(new_n293), .A3(new_n286), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT66), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n285), .A2(KEYINPUT66), .A3(new_n286), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n289), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n288), .B1(new_n298), .B2(KEYINPUT68), .ZN(new_n299));
  INV_X1    g098(.A(new_n289), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT66), .B1(new_n285), .B2(new_n286), .ZN(new_n301));
  AND4_X1   g100(.A1(KEYINPUT66), .A2(new_n291), .A3(new_n293), .A4(new_n286), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT68), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n284), .B1(new_n299), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n278), .A2(KEYINPUT23), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT23), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(G169gat), .B2(G176gat), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n307), .B(new_n309), .C1(new_n275), .C2(new_n276), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT25), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n313), .B1(G183gat), .B2(G190gat), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n280), .B1(KEYINPUT65), .B2(KEYINPUT24), .ZN(new_n315));
  AND2_X1   g114(.A1(KEYINPUT65), .A2(KEYINPUT24), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n312), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT24), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n314), .B1(new_n319), .B2(new_n280), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n311), .B1(new_n320), .B2(new_n310), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n306), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n274), .B1(new_n324), .B2(KEYINPUT29), .ZN(new_n325));
  INV_X1    g124(.A(new_n274), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n326), .B1(new_n306), .B2(new_n323), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n273), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  OAI211_X1 g127(.A(KEYINPUT68), .B(new_n300), .C1(new_n301), .C2(new_n302), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n287), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n296), .A2(new_n297), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT68), .B1(new_n331), .B2(new_n300), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n283), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT29), .B1(new_n333), .B2(new_n322), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n327), .B(new_n273), .C1(new_n334), .C2(new_n326), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n272), .B1(new_n328), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n327), .B1(new_n334), .B2(new_n326), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(new_n237), .ZN(new_n339));
  INV_X1    g138(.A(new_n272), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n339), .A2(new_n340), .A3(new_n335), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n337), .A2(KEYINPUT30), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT30), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n343), .B(new_n272), .C1(new_n328), .C2(new_n336), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n239), .A2(new_n250), .ZN(new_n347));
  XNOR2_X1  g146(.A(G113gat), .B(G120gat), .ZN(new_n348));
  INV_X1    g147(.A(G127gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n349), .A2(G134gat), .ZN(new_n350));
  INV_X1    g149(.A(G134gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n351), .A2(G127gat), .ZN(new_n352));
  OAI22_X1  g151(.A1(new_n348), .A2(KEYINPUT1), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(G120gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(G113gat), .ZN(new_n355));
  INV_X1    g154(.A(G113gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(G120gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G127gat), .B(G134gat), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT1), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  AND2_X1   g160(.A1(new_n353), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n362), .B1(KEYINPUT3), .B2(new_n219), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n362), .A2(new_n248), .A3(KEYINPUT4), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT4), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n353), .A2(new_n361), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n366), .B1(new_n219), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT75), .ZN(new_n369));
  AND3_X1   g168(.A1(new_n365), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n369), .B1(new_n365), .B2(new_n368), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n364), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT39), .ZN(new_n373));
  NAND2_X1  g172(.A1(G225gat), .A2(G233gat), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n372), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G1gat), .B(G29gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(KEYINPUT0), .ZN(new_n378));
  XNOR2_X1  g177(.A(G57gat), .B(G85gat), .ZN(new_n379));
  XOR2_X1   g178(.A(new_n378), .B(new_n379), .Z(new_n380));
  NAND2_X1  g179(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n248), .B(new_n367), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n374), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT39), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n384), .B1(new_n372), .B2(new_n375), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT40), .B1(new_n381), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n385), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT40), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n387), .A2(new_n388), .A3(new_n380), .A4(new_n376), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT5), .B1(new_n382), .B2(new_n374), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT4), .B1(new_n362), .B2(new_n248), .ZN(new_n391));
  NOR3_X1   g190(.A1(new_n219), .A2(new_n367), .A3(new_n366), .ZN(new_n392));
  NOR3_X1   g191(.A1(new_n391), .A2(new_n392), .A3(new_n375), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n390), .B1(new_n364), .B2(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n375), .A2(KEYINPUT5), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n364), .B(new_n395), .C1(new_n370), .C2(new_n371), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT76), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT75), .B1(new_n391), .B2(new_n392), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n365), .A2(new_n368), .A3(new_n369), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT76), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n400), .A2(new_n401), .A3(new_n364), .A4(new_n395), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n394), .B1(new_n397), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n380), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n386), .A2(new_n389), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n269), .B1(new_n346), .B2(new_n406), .ZN(new_n407));
  XOR2_X1   g206(.A(KEYINPUT77), .B(KEYINPUT6), .Z(new_n408));
  NOR2_X1   g207(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n405), .A2(new_n408), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NOR3_X1   g210(.A1(new_n403), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n402), .ZN(new_n413));
  INV_X1    g212(.A(new_n394), .ZN(new_n414));
  AND4_X1   g213(.A1(new_n413), .A2(new_n414), .A3(new_n408), .A4(new_n405), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT38), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT37), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n339), .A2(new_n418), .A3(new_n335), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n418), .B1(new_n339), .B2(new_n335), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n417), .B(new_n340), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n416), .A2(new_n421), .A3(KEYINPUT80), .A4(new_n337), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n340), .B1(new_n419), .B2(new_n420), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT38), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n337), .ZN(new_n426));
  NOR3_X1   g225(.A1(new_n426), .A2(new_n412), .A3(new_n415), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT80), .B1(new_n427), .B2(new_n421), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n407), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  OR3_X1    g228(.A1(new_n403), .A2(new_n409), .A3(new_n411), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n403), .A2(new_n408), .A3(new_n405), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n268), .B1(new_n345), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n367), .B1(new_n306), .B2(new_n323), .ZN(new_n434));
  NAND2_X1  g233(.A1(G227gat), .A2(G233gat), .ZN(new_n435));
  XOR2_X1   g234(.A(new_n435), .B(KEYINPUT64), .Z(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n333), .A2(new_n362), .A3(new_n322), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n434), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n439), .B(KEYINPUT34), .ZN(new_n440));
  XOR2_X1   g239(.A(G15gat), .B(G43gat), .Z(new_n441));
  XNOR2_X1  g240(.A(G71gat), .B(G99gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n437), .B1(new_n434), .B2(new_n438), .ZN(new_n444));
  XOR2_X1   g243(.A(KEYINPUT69), .B(KEYINPUT33), .Z(new_n445));
  OAI21_X1  g244(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT32), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n438), .ZN(new_n450));
  AOI221_X4 g249(.A(new_n447), .B1(new_n445), .B2(new_n443), .C1(new_n450), .C2(new_n436), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n440), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n450), .A2(new_n436), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT32), .ZN(new_n454));
  INV_X1    g253(.A(new_n445), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n456), .A3(new_n443), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT34), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n439), .B(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n446), .A2(new_n448), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n457), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n452), .A2(new_n461), .A3(KEYINPUT70), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT36), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT70), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n464), .B(new_n440), .C1(new_n449), .C2(new_n451), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n462), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n452), .A2(new_n461), .A3(KEYINPUT36), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n433), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n268), .A2(new_n452), .A3(new_n461), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n345), .A2(new_n432), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT35), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n462), .A2(new_n465), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n416), .B1(new_n344), .B2(new_n342), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT35), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n268), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n472), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  AOI22_X1  g275(.A1(new_n429), .A2(new_n468), .B1(new_n471), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G15gat), .B(G22gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT84), .ZN(new_n479));
  INV_X1    g278(.A(G1gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n478), .A2(KEYINPUT84), .A3(G1gat), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT16), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  OR2_X1    g284(.A1(new_n485), .A2(G8gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(G8gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT85), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n486), .A2(KEYINPUT85), .A3(new_n487), .ZN(new_n491));
  XOR2_X1   g290(.A(G43gat), .B(G50gat), .Z(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT81), .ZN(new_n495));
  OR2_X1    g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OR3_X1    g295(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n494), .A2(new_n495), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(G29gat), .ZN(new_n500));
  INV_X1    g299(.A(G36gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g301(.A(KEYINPUT15), .B(new_n493), .C1(new_n499), .C2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT17), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT15), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n492), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT83), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT83), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n492), .A2(new_n508), .A3(new_n505), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n493), .A2(KEYINPUT82), .A3(KEYINPUT15), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT82), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n513), .B1(new_n492), .B2(new_n505), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n502), .B1(new_n497), .B2(new_n494), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n512), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n503), .B(new_n504), .C1(new_n511), .C2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n510), .A2(new_n512), .A3(new_n514), .A4(new_n515), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n504), .B1(new_n519), .B2(new_n503), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n490), .B(new_n491), .C1(new_n518), .C2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(G229gat), .A2(G233gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n519), .A2(new_n503), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n488), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n521), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT18), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n524), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n486), .A2(KEYINPUT85), .A3(new_n487), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT85), .B1(new_n486), .B2(new_n487), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n523), .A2(KEYINPUT17), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n517), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n528), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n534), .A2(KEYINPUT18), .A3(new_n522), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n522), .B(KEYINPUT13), .Z(new_n536));
  NOR2_X1   g335(.A1(new_n488), .A2(new_n523), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n536), .B1(new_n528), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n527), .A2(new_n535), .A3(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G113gat), .B(G141gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(G197gat), .ZN(new_n541));
  XOR2_X1   g340(.A(KEYINPUT11), .B(G169gat), .Z(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT12), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n539), .B(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n477), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT93), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT7), .ZN(new_n548));
  NAND2_X1  g347(.A1(G85gat), .A2(G92gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(G99gat), .A2(G106gat), .ZN(new_n551));
  INV_X1    g350(.A(G85gat), .ZN(new_n552));
  INV_X1    g351(.A(G92gat), .ZN(new_n553));
  AOI22_X1  g352(.A1(KEYINPUT8), .A2(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT94), .ZN(new_n555));
  OR2_X1    g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n555), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n550), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT95), .ZN(new_n559));
  XOR2_X1   g358(.A(G99gat), .B(G106gat), .Z(new_n560));
  NAND3_X1  g359(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n549), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(new_n548), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n554), .A2(new_n555), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n554), .A2(new_n555), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n560), .A2(new_n559), .ZN(new_n567));
  INV_X1    g366(.A(new_n560), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(KEYINPUT95), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n561), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n571), .B1(new_n532), .B2(new_n517), .ZN(new_n572));
  AND2_X1   g371(.A1(G232gat), .A2(G233gat), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n523), .A2(new_n571), .B1(KEYINPUT41), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G190gat), .B(G218gat), .ZN(new_n576));
  OR3_X1    g375(.A1(new_n572), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n576), .B1(new_n572), .B2(new_n575), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT96), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n573), .A2(KEYINPUT41), .ZN(new_n582));
  XNOR2_X1  g381(.A(G134gat), .B(G162gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n579), .B1(new_n581), .B2(new_n585), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n577), .A2(KEYINPUT96), .A3(new_n578), .A4(new_n584), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT21), .ZN(new_n590));
  XNOR2_X1  g389(.A(G71gat), .B(G78gat), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT9), .ZN(new_n593));
  XNOR2_X1  g392(.A(G57gat), .B(G64gat), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT86), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  OR2_X1    g396(.A1(G57gat), .A2(G64gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(G57gat), .A2(G64gat), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n598), .A2(KEYINPUT86), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n597), .A2(new_n591), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT87), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n595), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(KEYINPUT88), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT88), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n606), .B(new_n595), .C1(new_n601), .C2(new_n603), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT91), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n605), .A2(KEYINPUT91), .A3(new_n607), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n590), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OR3_X1    g411(.A1(new_n612), .A2(KEYINPUT92), .A3(new_n488), .ZN(new_n613));
  OAI21_X1  g412(.A(KEYINPUT92), .B1(new_n612), .B2(new_n488), .ZN(new_n614));
  XOR2_X1   g413(.A(G127gat), .B(G155gat), .Z(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT20), .ZN(new_n616));
  NAND2_X1  g415(.A1(G231gat), .A2(G233gat), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n617), .B(KEYINPUT89), .Z(new_n618));
  XNOR2_X1  g417(.A(new_n616), .B(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  AND3_X1   g419(.A1(new_n613), .A2(new_n614), .A3(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n608), .A2(KEYINPUT21), .ZN(new_n622));
  XNOR2_X1  g421(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G183gat), .B(G211gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n620), .B1(new_n613), .B2(new_n614), .ZN(new_n627));
  OR3_X1    g426(.A1(new_n621), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n626), .B1(new_n621), .B2(new_n627), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n589), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(G230gat), .A2(G233gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT98), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  AND3_X1   g433(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n567), .B1(new_n566), .B2(new_n569), .ZN(new_n636));
  OAI21_X1  g435(.A(KEYINPUT10), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n637), .B1(new_n610), .B2(new_n611), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n605), .A2(new_n561), .A3(new_n570), .A4(new_n607), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT10), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT97), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n568), .B1(new_n558), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n604), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n566), .A2(KEYINPUT97), .A3(new_n560), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  AND3_X1   g444(.A1(new_n639), .A2(new_n640), .A3(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n634), .B1(new_n638), .B2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G120gat), .B(G148gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(G176gat), .B(G204gat), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n648), .B(new_n649), .Z(new_n650));
  AOI21_X1  g449(.A(new_n634), .B1(new_n639), .B2(new_n645), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n647), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n647), .A2(new_n654), .ZN(new_n655));
  OAI211_X1 g454(.A(KEYINPUT100), .B(new_n634), .C1(new_n638), .C2(new_n646), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n651), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n650), .B(KEYINPUT99), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n653), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n631), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n546), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT101), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n546), .A2(KEYINPUT101), .A3(new_n661), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n416), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT102), .B(G1gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1324gat));
  XOR2_X1   g468(.A(KEYINPUT16), .B(G8gat), .Z(new_n670));
  NAND3_X1  g469(.A1(new_n666), .A2(new_n346), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n666), .A2(new_n346), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(G8gat), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n671), .ZN(new_n674));
  MUX2_X1   g473(.A(new_n671), .B(new_n674), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g474(.A1(new_n466), .A2(new_n467), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n666), .A2(G15gat), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(G15gat), .B1(new_n666), .B2(new_n472), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n678), .B1(new_n681), .B2(new_n682), .ZN(G1326gat));
  NAND2_X1  g482(.A1(new_n666), .A2(new_n269), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT43), .B(G22gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  NOR3_X1   g485(.A1(new_n589), .A2(new_n630), .A3(new_n660), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n546), .A2(new_n500), .A3(new_n416), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT45), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n429), .A2(new_n468), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n476), .A2(new_n471), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n692), .A2(KEYINPUT105), .A3(new_n588), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n477), .A2(KEYINPUT106), .A3(new_n589), .ZN(new_n694));
  OAI211_X1 g493(.A(KEYINPUT44), .B(new_n693), .C1(new_n694), .C2(KEYINPUT105), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n692), .A2(new_n588), .ZN(new_n698));
  OAI211_X1 g497(.A(new_n696), .B(new_n697), .C1(new_n698), .C2(KEYINPUT106), .ZN(new_n699));
  INV_X1    g498(.A(new_n630), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n700), .A2(KEYINPUT104), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n700), .A2(KEYINPUT104), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n703), .A2(new_n545), .A3(new_n660), .ZN(new_n704));
  AND4_X1   g503(.A1(new_n416), .A2(new_n695), .A3(new_n699), .A4(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n689), .B1(new_n705), .B2(new_n500), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1328gat));
  NAND4_X1  g507(.A1(new_n546), .A2(new_n501), .A3(new_n346), .A4(new_n687), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(KEYINPUT46), .Z(new_n710));
  AND4_X1   g509(.A1(new_n346), .A2(new_n695), .A3(new_n699), .A4(new_n704), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n710), .B1(new_n711), .B2(new_n501), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(G1329gat));
  NAND2_X1  g513(.A1(new_n546), .A2(new_n687), .ZN(new_n715));
  INV_X1    g514(.A(new_n472), .ZN(new_n716));
  OR3_X1    g515(.A1(new_n715), .A2(G43gat), .A3(new_n716), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n695), .A2(new_n677), .A3(new_n699), .A4(new_n704), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT110), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(G43gat), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n718), .A2(KEYINPUT110), .ZN(new_n721));
  OAI211_X1 g520(.A(KEYINPUT47), .B(new_n717), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT109), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n718), .A2(G43gat), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n717), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n723), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  AOI211_X1 g526(.A(KEYINPUT109), .B(KEYINPUT47), .C1(new_n724), .C2(new_n717), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n722), .B1(new_n727), .B2(new_n728), .ZN(G1330gat));
  INV_X1    g528(.A(KEYINPUT112), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n695), .A2(new_n269), .A3(new_n699), .A4(new_n704), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(G50gat), .ZN(new_n732));
  OR2_X1    g531(.A1(new_n268), .A2(G50gat), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n715), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  XOR2_X1   g535(.A(KEYINPUT111), .B(KEYINPUT48), .Z(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n730), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n734), .B1(new_n731), .B2(G50gat), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n740), .A2(KEYINPUT112), .A3(new_n737), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT113), .ZN(new_n742));
  AND4_X1   g541(.A1(new_n742), .A2(new_n732), .A3(KEYINPUT48), .A4(new_n735), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n742), .B1(new_n740), .B2(KEYINPUT48), .ZN(new_n744));
  OAI22_X1  g543(.A1(new_n739), .A2(new_n741), .B1(new_n743), .B2(new_n744), .ZN(G1331gat));
  INV_X1    g544(.A(new_n545), .ZN(new_n746));
  INV_X1    g545(.A(new_n653), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n655), .A2(new_n656), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n652), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n747), .B1(new_n749), .B2(new_n658), .ZN(new_n750));
  NOR4_X1   g549(.A1(new_n477), .A2(new_n746), .A3(new_n631), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n416), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(G57gat), .ZN(G1332gat));
  AND2_X1   g552(.A1(new_n751), .A2(new_n346), .ZN(new_n754));
  NOR2_X1   g553(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n755));
  AND2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(new_n754), .B2(new_n755), .ZN(G1333gat));
  NAND2_X1  g557(.A1(new_n751), .A2(new_n677), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n716), .A2(G71gat), .ZN(new_n760));
  AOI22_X1  g559(.A1(new_n759), .A2(G71gat), .B1(new_n751), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g561(.A1(new_n751), .A2(new_n269), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g563(.A1(new_n630), .A2(new_n746), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n695), .A2(new_n660), .A3(new_n699), .A4(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(G85gat), .B1(new_n766), .B2(new_n432), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n692), .A2(new_n588), .A3(new_n765), .ZN(new_n768));
  XOR2_X1   g567(.A(new_n768), .B(KEYINPUT51), .Z(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n660), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n416), .A2(new_n552), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n767), .B1(new_n770), .B2(new_n771), .ZN(G1336gat));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n750), .A2(new_n345), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n769), .A2(new_n553), .A3(new_n774), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n695), .A2(new_n699), .A3(new_n765), .A4(new_n774), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT114), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(G92gat), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n776), .A2(KEYINPUT114), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n773), .B(new_n775), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n776), .A2(G92gat), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n775), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n780), .B1(new_n773), .B2(new_n782), .ZN(G1337gat));
  OAI21_X1  g582(.A(G99gat), .B1(new_n766), .B2(new_n676), .ZN(new_n784));
  OR2_X1    g583(.A1(new_n716), .A2(G99gat), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n784), .B1(new_n770), .B2(new_n785), .ZN(G1338gat));
  XNOR2_X1  g585(.A(KEYINPUT115), .B(G106gat), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n787), .B1(new_n766), .B2(new_n268), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n750), .A2(G106gat), .A3(new_n268), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(KEYINPUT116), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n769), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g592(.A1(new_n661), .A2(new_n545), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n639), .A2(new_n645), .A3(new_n640), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n605), .A2(KEYINPUT91), .A3(new_n607), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT91), .B1(new_n605), .B2(new_n607), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n633), .B(new_n796), .C1(new_n799), .C2(new_n637), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n647), .A2(KEYINPUT54), .A3(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT117), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n801), .B(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n655), .A2(new_n804), .A3(new_n656), .ZN(new_n805));
  INV_X1    g604(.A(new_n650), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT118), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n805), .A2(new_n809), .A3(new_n806), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n803), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n747), .B1(new_n811), .B2(KEYINPUT55), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n527), .A2(new_n535), .A3(new_n538), .ZN(new_n813));
  OAI21_X1  g612(.A(KEYINPUT119), .B1(new_n534), .B2(new_n522), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n521), .A2(new_n524), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT119), .ZN(new_n816));
  INV_X1    g615(.A(new_n522), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  OR3_X1    g617(.A1(new_n528), .A2(new_n537), .A3(new_n536), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n814), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  AOI22_X1  g619(.A1(new_n813), .A2(new_n544), .B1(new_n820), .B2(new_n543), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n801), .B(KEYINPUT117), .ZN(new_n822));
  AND3_X1   g621(.A1(new_n805), .A2(new_n809), .A3(new_n806), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n809), .B1(new_n805), .B2(new_n806), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n812), .A2(new_n588), .A3(new_n821), .A4(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n522), .B1(new_n521), .B2(new_n524), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n819), .B1(new_n829), .B2(new_n816), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n534), .A2(KEYINPUT119), .A3(new_n522), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n543), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n527), .A2(new_n535), .A3(new_n544), .A4(new_n538), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT120), .B1(new_n750), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT120), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n821), .A2(new_n660), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n545), .B1(new_n825), .B2(new_n826), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n838), .B1(new_n812), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n828), .B1(new_n840), .B2(new_n588), .ZN(new_n841));
  INV_X1    g640(.A(new_n703), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n795), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n346), .A2(new_n432), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n716), .A2(new_n269), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n847), .A2(new_n356), .A3(new_n545), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n843), .A2(new_n432), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n469), .A2(new_n346), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n746), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n848), .B1(new_n853), .B2(new_n356), .ZN(G1340gat));
  NOR3_X1   g653(.A1(new_n847), .A2(new_n354), .A3(new_n750), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n852), .A2(new_n660), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n855), .B1(new_n856), .B2(new_n354), .ZN(G1341gat));
  OAI21_X1  g656(.A(G127gat), .B1(new_n847), .B2(new_n842), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n630), .A2(new_n349), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n858), .B1(new_n851), .B2(new_n859), .ZN(G1342gat));
  NAND3_X1  g659(.A1(new_n852), .A2(new_n351), .A3(new_n588), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n862));
  OAI21_X1  g661(.A(G134gat), .B1(new_n847), .B2(new_n589), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(G1343gat));
  NAND2_X1  g664(.A1(new_n676), .A2(new_n845), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n268), .A2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n869));
  OAI211_X1 g668(.A(KEYINPUT55), .B(new_n822), .C1(new_n823), .C2(new_n824), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n827), .A2(new_n746), .A3(new_n653), .A4(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n750), .A2(new_n834), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n588), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n827), .A2(new_n588), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n870), .A2(new_n653), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n875), .A2(new_n876), .A3(new_n834), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n869), .B(new_n700), .C1(new_n874), .C2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n794), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n872), .B1(new_n812), .B2(new_n839), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n828), .B1(new_n880), .B2(new_n588), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n869), .B1(new_n881), .B2(new_n700), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n868), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n867), .B1(new_n843), .B2(new_n268), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n866), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n212), .B1(new_n885), .B2(new_n746), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n849), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(KEYINPUT122), .B1(new_n843), .B2(new_n432), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n676), .A2(new_n269), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n890), .A2(new_n346), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n545), .A2(G141gat), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n888), .A2(new_n889), .A3(new_n891), .A4(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT58), .B1(new_n886), .B2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT58), .ZN(new_n896));
  AOI211_X1 g695(.A(new_n545), .B(new_n866), .C1(new_n883), .C2(new_n884), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n896), .B(new_n893), .C1(new_n897), .C2(new_n212), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n895), .A2(new_n898), .ZN(G1344gat));
  AOI211_X1 g698(.A(KEYINPUT59), .B(new_n208), .C1(new_n885), .C2(new_n660), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n902), .B1(new_n875), .B2(new_n876), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n812), .A2(KEYINPUT124), .A3(new_n588), .A4(new_n827), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n903), .A2(new_n821), .A3(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n874), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n630), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n867), .B(new_n269), .C1(new_n907), .C2(new_n795), .ZN(new_n908));
  OAI21_X1  g707(.A(KEYINPUT57), .B1(new_n843), .B2(new_n268), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n866), .A2(new_n750), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n901), .B1(new_n911), .B2(G148gat), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT123), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n750), .A2(G148gat), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n917));
  INV_X1    g716(.A(new_n915), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n917), .A2(KEYINPUT123), .A3(new_n918), .ZN(new_n919));
  OAI22_X1  g718(.A1(new_n900), .A2(new_n912), .B1(new_n916), .B2(new_n919), .ZN(G1345gat));
  INV_X1    g719(.A(G155gat), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n914), .A2(new_n921), .A3(new_n630), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n885), .A2(new_n703), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n923), .B2(new_n921), .ZN(G1346gat));
  AOI21_X1  g723(.A(G162gat), .B1(new_n914), .B2(new_n588), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n588), .A2(G162gat), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n925), .B1(new_n885), .B2(new_n926), .ZN(G1347gat));
  NOR2_X1   g726(.A1(new_n345), .A2(new_n416), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n844), .A2(new_n846), .A3(new_n928), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n929), .A2(new_n275), .A3(new_n545), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n844), .A2(new_n432), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n931), .A2(new_n469), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n346), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(new_n746), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n930), .B1(new_n935), .B2(new_n275), .ZN(G1348gat));
  NAND3_X1  g735(.A1(new_n932), .A2(new_n276), .A3(new_n774), .ZN(new_n937));
  OAI21_X1  g736(.A(G176gat), .B1(new_n929), .B2(new_n750), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1349gat));
  OAI21_X1  g738(.A(G183gat), .B1(new_n929), .B2(new_n842), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n630), .A2(new_n285), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n933), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(KEYINPUT60), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT60), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n944), .B(new_n940), .C1(new_n933), .C2(new_n941), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n945), .ZN(G1350gat));
  NAND3_X1  g745(.A1(new_n934), .A2(new_n286), .A3(new_n588), .ZN(new_n947));
  OAI21_X1  g746(.A(G190gat), .B1(new_n929), .B2(new_n589), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n948), .A2(KEYINPUT61), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n948), .A2(KEYINPUT61), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(G1351gat));
  NOR2_X1   g750(.A1(new_n545), .A2(G197gat), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT125), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n843), .A2(new_n416), .A3(new_n890), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n953), .B1(new_n954), .B2(new_n346), .ZN(new_n955));
  INV_X1    g754(.A(new_n890), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n750), .A2(new_n834), .A3(KEYINPUT120), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n836), .B1(new_n821), .B2(new_n660), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n746), .B1(new_n811), .B2(KEYINPUT55), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n959), .B1(new_n960), .B2(new_n876), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(new_n589), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n703), .B1(new_n962), .B2(new_n828), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n432), .B(new_n956), .C1(new_n963), .C2(new_n795), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n964), .A2(KEYINPUT125), .A3(new_n345), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n952), .B1(new_n955), .B2(new_n965), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n676), .A2(new_n928), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n908), .A2(new_n746), .A3(new_n909), .A4(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(KEYINPUT126), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(G197gat), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n968), .A2(KEYINPUT126), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n966), .B1(new_n970), .B2(new_n971), .ZN(G1352gat));
  AND2_X1   g771(.A1(new_n908), .A2(new_n909), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n973), .A2(new_n660), .A3(new_n967), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(G204gat), .ZN(new_n975));
  OR3_X1    g774(.A1(new_n750), .A2(G204gat), .A3(new_n345), .ZN(new_n976));
  OAI21_X1  g775(.A(KEYINPUT62), .B1(new_n964), .B2(new_n976), .ZN(new_n977));
  OR3_X1    g776(.A1(new_n964), .A2(KEYINPUT62), .A3(new_n976), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n975), .A2(new_n977), .A3(new_n978), .ZN(G1353gat));
  OAI211_X1 g778(.A(new_n221), .B(new_n630), .C1(new_n955), .C2(new_n965), .ZN(new_n980));
  NAND4_X1  g779(.A1(new_n908), .A2(new_n630), .A3(new_n909), .A4(new_n967), .ZN(new_n981));
  AND3_X1   g780(.A1(new_n981), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n982));
  AOI21_X1  g781(.A(KEYINPUT63), .B1(new_n981), .B2(G211gat), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(G1354gat));
  AND4_X1   g783(.A1(G218gat), .A2(new_n973), .A3(new_n588), .A4(new_n967), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n588), .B1(new_n955), .B2(new_n965), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT127), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n986), .A2(new_n987), .A3(new_n222), .ZN(new_n988));
  OAI21_X1  g787(.A(KEYINPUT125), .B1(new_n964), .B2(new_n345), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n843), .A2(new_n416), .ZN(new_n990));
  NAND4_X1  g789(.A1(new_n990), .A2(new_n953), .A3(new_n346), .A4(new_n956), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n589), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g791(.A(KEYINPUT127), .B1(new_n992), .B2(G218gat), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n985), .B1(new_n988), .B2(new_n993), .ZN(G1355gat));
endmodule


