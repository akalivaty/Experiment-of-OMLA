//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 1 1 0 0 0 1 1 0 1 0 1 1 0 0 1 1 1 0 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015;
  INV_X1    g000(.A(KEYINPUT29), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT69), .B1(new_n188), .B2(G116), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT69), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n188), .A2(G116), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT2), .ZN(new_n196));
  INV_X1    g010(.A(G113), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n197), .A3(KEYINPUT67), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT67), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n199), .B1(KEYINPUT2), .B2(G113), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(KEYINPUT2), .A2(G113), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT68), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT68), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT2), .A3(G113), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n201), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n195), .A2(new_n207), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n193), .A2(new_n201), .A3(new_n206), .A4(new_n194), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G143), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  OAI211_X1 g029(.A(KEYINPUT65), .B(KEYINPUT1), .C1(new_n213), .C2(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G128), .ZN(new_n217));
  AOI21_X1  g031(.A(KEYINPUT65), .B1(new_n212), .B2(KEYINPUT1), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n215), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n215), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT1), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(G128), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT11), .ZN(new_n224));
  INV_X1    g038(.A(G134), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n224), .B1(new_n225), .B2(G137), .ZN(new_n226));
  INV_X1    g040(.A(G137), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(KEYINPUT11), .A3(G134), .ZN(new_n228));
  INV_X1    g042(.A(G131), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n225), .A2(G137), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n226), .A2(new_n228), .A3(new_n229), .A4(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n227), .A2(G134), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n225), .A2(G137), .ZN(new_n233));
  OAI21_X1  g047(.A(G131), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n226), .A2(new_n230), .A3(new_n228), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G131), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n231), .ZN(new_n239));
  OR2_X1    g053(.A1(KEYINPUT0), .A2(G128), .ZN(new_n240));
  NAND2_X1  g054(.A1(KEYINPUT0), .A2(G128), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n215), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n212), .A2(new_n214), .A3(new_n241), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n223), .A2(new_n236), .B1(new_n239), .B2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT70), .B1(new_n246), .B2(KEYINPUT30), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n235), .B1(new_n219), .B2(new_n222), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n238), .A2(new_n231), .B1(new_n243), .B2(new_n244), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT30), .ZN(new_n251));
  NOR4_X1   g065(.A1(new_n248), .A2(new_n249), .A3(new_n250), .A4(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n223), .A2(new_n236), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n212), .A2(new_n214), .B1(new_n240), .B2(new_n241), .ZN(new_n254));
  AND3_X1   g068(.A1(new_n212), .A2(new_n214), .A3(new_n241), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT64), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT64), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n243), .A2(new_n257), .A3(new_n244), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n239), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n253), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(KEYINPUT66), .B1(new_n260), .B2(new_n251), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT66), .ZN(new_n262));
  AOI211_X1 g076(.A(new_n262), .B(KEYINPUT30), .C1(new_n253), .C2(new_n259), .ZN(new_n263));
  OAI221_X1 g077(.A(new_n210), .B1(new_n247), .B2(new_n252), .C1(new_n261), .C2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n210), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n246), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n267));
  INV_X1    g081(.A(G101), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n267), .B(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(G237), .A2(G953), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G210), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n269), .B(new_n271), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n264), .A2(new_n266), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n265), .B1(new_n253), .B2(new_n259), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT71), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n266), .B1(new_n274), .B2(new_n275), .ZN(new_n278));
  OAI21_X1  g092(.A(KEYINPUT28), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT28), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n266), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n272), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n187), .B1(new_n273), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n210), .B1(new_n248), .B2(new_n249), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n266), .A2(KEYINPUT73), .A3(new_n284), .ZN(new_n285));
  OR3_X1    g099(.A1(new_n246), .A2(KEYINPUT73), .A3(new_n265), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(new_n286), .A3(KEYINPUT28), .ZN(new_n287));
  NOR3_X1   g101(.A1(new_n248), .A2(new_n210), .A3(new_n249), .ZN(new_n288));
  OR3_X1    g102(.A1(new_n288), .A2(KEYINPUT74), .A3(KEYINPUT28), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n281), .A2(KEYINPUT74), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n272), .A2(new_n187), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n287), .A2(new_n289), .A3(new_n290), .A4(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT75), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n292), .B(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G902), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n283), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G472), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n288), .A2(new_n272), .ZN(new_n298));
  OAI22_X1  g112(.A1(new_n261), .A2(new_n263), .B1(new_n247), .B2(new_n252), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n298), .B1(new_n299), .B2(new_n265), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT31), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n260), .A2(new_n210), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n288), .B1(new_n302), .B2(KEYINPUT71), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n280), .B1(new_n303), .B2(new_n276), .ZN(new_n304));
  INV_X1    g118(.A(new_n281), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n272), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT31), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n264), .A2(new_n307), .A3(new_n298), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n301), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(G472), .A2(G902), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(KEYINPUT32), .B1(new_n311), .B2(KEYINPUT72), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT72), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT32), .ZN(new_n314));
  AOI211_X1 g128(.A(new_n313), .B(new_n314), .C1(new_n309), .C2(new_n310), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n297), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(G214), .B1(G237), .B2(G902), .ZN(new_n317));
  NAND2_X1  g131(.A1(G234), .A2(G237), .ZN(new_n318));
  INV_X1    g132(.A(G953), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(G952), .A3(new_n319), .ZN(new_n320));
  XOR2_X1   g134(.A(KEYINPUT21), .B(G898), .Z(new_n321));
  NAND3_X1  g135(.A1(new_n318), .A2(G902), .A3(G953), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n245), .A2(G125), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n219), .A2(new_n222), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n324), .B1(new_n325), .B2(G125), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT85), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT85), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n328), .B(new_n324), .C1(new_n325), .C2(G125), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G224), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n331), .A2(G953), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n330), .B(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT6), .ZN(new_n334));
  XNOR2_X1  g148(.A(G110), .B(G122), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G107), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT81), .B1(new_n337), .B2(G104), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT81), .ZN(new_n339));
  INV_X1    g153(.A(G104), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(new_n340), .A3(G107), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT3), .B1(new_n340), .B2(G107), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT3), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(new_n337), .A3(G104), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n342), .A2(new_n268), .A3(new_n343), .A4(new_n345), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n343), .A2(new_n338), .A3(new_n345), .A4(new_n341), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G101), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(KEYINPUT4), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT4), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n347), .A2(new_n350), .A3(G101), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n349), .A2(new_n210), .A3(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n340), .A2(G107), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n337), .A2(G104), .ZN(new_n354));
  OAI21_X1  g168(.A(G101), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n355), .B1(new_n347), .B2(G101), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT5), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n358), .A2(new_n188), .A3(G116), .ZN(new_n359));
  OAI211_X1 g173(.A(G113), .B(new_n359), .C1(new_n195), .C2(new_n358), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n357), .A2(new_n209), .A3(new_n360), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n352), .A2(KEYINPUT84), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT84), .B1(new_n352), .B2(new_n361), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n336), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n352), .A2(new_n361), .A3(new_n335), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n334), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n352), .A2(new_n361), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT84), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n352), .A2(new_n361), .A3(KEYINPUT84), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT6), .B1(new_n371), .B2(new_n336), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n333), .B1(new_n366), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(G210), .B1(G237), .B2(G902), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n360), .A2(new_n209), .ZN(new_n375));
  OAI211_X1 g189(.A(KEYINPUT86), .B(new_n355), .C1(new_n347), .C2(G101), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n360), .A2(new_n209), .A3(new_n376), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n335), .B(KEYINPUT8), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT7), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n332), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n326), .A2(new_n383), .ZN(new_n384));
  OAI221_X1 g198(.A(new_n324), .B1(new_n382), .B2(new_n332), .C1(new_n325), .C2(G125), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n381), .A2(new_n365), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n295), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT87), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n386), .A2(KEYINPUT87), .A3(new_n295), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n373), .A2(new_n374), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n374), .B1(new_n373), .B2(new_n391), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n317), .B(new_n323), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G237), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(new_n319), .A3(G214), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n213), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n270), .A2(G143), .A3(G214), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(KEYINPUT90), .B1(new_n399), .B2(G131), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT90), .ZN(new_n401));
  AOI211_X1 g215(.A(new_n401), .B(new_n229), .C1(new_n397), .C2(new_n398), .ZN(new_n402));
  OAI21_X1  g216(.A(KEYINPUT17), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT78), .ZN(new_n404));
  INV_X1    g218(.A(G140), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G125), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n404), .B1(new_n406), .B2(KEYINPUT16), .ZN(new_n407));
  INV_X1    g221(.A(G125), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(G140), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n406), .A2(new_n409), .A3(KEYINPUT16), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT16), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n411), .A2(new_n405), .A3(KEYINPUT78), .A4(G125), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n407), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n211), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n407), .A2(new_n410), .A3(G146), .A4(new_n412), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AND4_X1   g230(.A1(G143), .A2(new_n395), .A3(new_n319), .A4(G214), .ZN(new_n417));
  AOI21_X1  g231(.A(G143), .B1(new_n270), .B2(G214), .ZN(new_n418));
  OAI21_X1  g232(.A(G131), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n401), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n399), .A2(KEYINPUT90), .A3(G131), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n417), .A2(new_n418), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n229), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT17), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n420), .A2(new_n421), .A3(new_n423), .A4(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n403), .A2(new_n416), .A3(new_n425), .ZN(new_n426));
  XOR2_X1   g240(.A(G113), .B(G122), .Z(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(KEYINPUT92), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n428), .B(new_n340), .ZN(new_n429));
  NAND3_X1  g243(.A1(KEYINPUT88), .A2(KEYINPUT18), .A3(G131), .ZN(new_n430));
  OR2_X1    g244(.A1(new_n422), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n422), .A2(new_n430), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n406), .A2(new_n409), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G146), .ZN(new_n434));
  XNOR2_X1  g248(.A(G125), .B(G140), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n211), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT89), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n434), .A2(new_n436), .A3(KEYINPUT89), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n431), .B(new_n432), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n426), .A2(new_n429), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n429), .B1(new_n426), .B2(new_n439), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n295), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G475), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT13), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(new_n213), .A3(G128), .ZN(new_n445));
  XOR2_X1   g259(.A(G128), .B(G143), .Z(new_n446));
  OAI211_X1 g260(.A(G134), .B(new_n445), .C1(new_n446), .C2(new_n444), .ZN(new_n447));
  INV_X1    g261(.A(G122), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(G116), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n191), .A2(G122), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(G107), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n449), .A2(new_n450), .A3(new_n337), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n447), .B(new_n454), .C1(G134), .C2(new_n446), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n191), .A2(KEYINPUT14), .A3(G122), .ZN(new_n456));
  OAI211_X1 g270(.A(G107), .B(new_n456), .C1(new_n451), .C2(KEYINPUT14), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n446), .A2(G134), .ZN(new_n458));
  XNOR2_X1  g272(.A(G128), .B(G143), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n459), .A2(new_n225), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n457), .B(new_n453), .C1(new_n458), .C2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  OR2_X1    g276(.A1(KEYINPUT9), .A2(G234), .ZN(new_n463));
  NAND2_X1  g277(.A1(KEYINPUT9), .A2(G234), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n463), .A2(G217), .A3(new_n319), .A4(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT94), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n465), .B(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n462), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n455), .A2(new_n461), .A3(new_n467), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(G478), .ZN(new_n472));
  NOR2_X1   g286(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT96), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n476), .B(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n471), .A2(new_n295), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(G902), .B1(new_n469), .B2(new_n470), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n476), .A2(new_n477), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(G475), .A2(G902), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n420), .A2(new_n421), .A3(new_n423), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n433), .A2(KEYINPUT19), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT19), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n435), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n487), .A2(new_n489), .A3(KEYINPUT91), .A4(new_n211), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT91), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n487), .A2(new_n489), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n491), .B1(new_n492), .B2(G146), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n486), .A2(new_n415), .A3(new_n490), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n439), .ZN(new_n495));
  INV_X1    g309(.A(new_n429), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n426), .A2(new_n429), .A3(new_n439), .ZN(new_n498));
  AOI211_X1 g312(.A(KEYINPUT20), .B(new_n485), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n429), .B1(new_n494), .B2(new_n439), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n484), .B1(new_n440), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT20), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n499), .B1(new_n502), .B2(KEYINPUT93), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT93), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n501), .A2(new_n504), .A3(KEYINPUT20), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n443), .B(new_n483), .C1(new_n503), .C2(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n394), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT79), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT77), .ZN(new_n509));
  INV_X1    g323(.A(G128), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n509), .B1(G119), .B2(new_n510), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n188), .A2(KEYINPUT77), .A3(G128), .ZN(new_n512));
  OAI22_X1  g326(.A1(new_n511), .A2(new_n512), .B1(G119), .B2(new_n510), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT24), .B(G110), .ZN(new_n514));
  OAI21_X1  g328(.A(KEYINPUT23), .B1(new_n188), .B2(G128), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT23), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(new_n510), .A3(G119), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n515), .A2(new_n517), .B1(new_n188), .B2(G128), .ZN(new_n518));
  INV_X1    g332(.A(G110), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n513), .A2(new_n514), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n415), .A2(new_n436), .ZN(new_n521));
  OAI22_X1  g335(.A1(new_n513), .A2(new_n514), .B1(new_n518), .B2(new_n519), .ZN(new_n522));
  OAI221_X1 g336(.A(new_n508), .B1(new_n520), .B2(new_n521), .C1(new_n416), .C2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n522), .B1(new_n414), .B2(new_n415), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n520), .A2(new_n521), .ZN(new_n525));
  OAI21_X1  g339(.A(KEYINPUT79), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n319), .A2(G221), .A3(G234), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(KEYINPUT22), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(G137), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n523), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n524), .A2(new_n525), .ZN(new_n531));
  INV_X1    g345(.A(new_n529), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n508), .A3(new_n532), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT25), .B1(new_n534), .B2(G902), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n530), .A2(new_n533), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT25), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(new_n537), .A3(new_n295), .ZN(new_n538));
  INV_X1    g352(.A(G234), .ZN(new_n539));
  OAI21_X1  g353(.A(G217), .B1(new_n539), .B2(G902), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(KEYINPUT76), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n535), .A2(new_n538), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n540), .A2(new_n295), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n536), .A2(new_n544), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n463), .A2(new_n464), .ZN(new_n547));
  OAI21_X1  g361(.A(G221), .B1(new_n547), .B2(G902), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n349), .A2(new_n245), .A3(new_n351), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n357), .A2(KEYINPUT10), .A3(new_n223), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT10), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n510), .B1(new_n212), .B2(KEYINPUT1), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n220), .A2(new_n553), .ZN(new_n554));
  NOR3_X1   g368(.A1(new_n215), .A2(KEYINPUT1), .A3(new_n510), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n552), .B1(new_n556), .B2(new_n356), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n550), .A2(new_n551), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n239), .ZN(new_n559));
  INV_X1    g373(.A(new_n239), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n550), .A2(new_n557), .A3(new_n551), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(G110), .B(G140), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(KEYINPUT80), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n319), .A2(G227), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n564), .B(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT83), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n562), .A2(KEYINPUT83), .A3(new_n566), .ZN(new_n570));
  INV_X1    g384(.A(new_n566), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n561), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n346), .B(new_n355), .C1(new_n555), .C2(new_n554), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n356), .A2(new_n222), .A3(new_n219), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(new_n574), .A3(KEYINPUT82), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT82), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n325), .A2(new_n576), .A3(new_n356), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n575), .A2(KEYINPUT12), .A3(new_n239), .A4(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT12), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n573), .A2(new_n574), .A3(KEYINPUT82), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n239), .B1(new_n574), .B2(KEYINPUT82), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n572), .B1(new_n578), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n569), .A2(new_n570), .A3(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(G469), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n586), .A3(new_n295), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n586), .A2(new_n295), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n582), .A2(new_n578), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n571), .B1(new_n589), .B2(new_n561), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n559), .A2(new_n561), .A3(new_n571), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n588), .B1(new_n593), .B2(G469), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n549), .B1(new_n587), .B2(new_n594), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n316), .A2(new_n507), .A3(new_n546), .A4(new_n595), .ZN(new_n596));
  XOR2_X1   g410(.A(KEYINPUT97), .B(G101), .Z(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(G3));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n599));
  INV_X1    g413(.A(G472), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n309), .B2(new_n295), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n311), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n587), .A2(new_n594), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n604), .A2(new_n546), .A3(new_n548), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n599), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n309), .A2(new_n310), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n607), .A2(new_n601), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n608), .A2(KEYINPUT98), .A3(new_n546), .A4(new_n595), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n443), .B1(new_n503), .B2(new_n505), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT99), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n455), .A2(new_n461), .A3(new_n467), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n467), .B1(new_n455), .B2(new_n461), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n611), .B(KEYINPUT33), .C1(new_n612), .C2(new_n613), .ZN(new_n617));
  AOI21_X1  g431(.A(G902), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(G478), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n480), .A2(G478), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n610), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n394), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n606), .A2(new_n609), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT34), .B(G104), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G6));
  NAND2_X1  g441(.A1(new_n497), .A2(new_n498), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT20), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n628), .A2(new_n629), .A3(new_n484), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n502), .A2(new_n630), .B1(G475), .B2(new_n442), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n482), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n394), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n606), .A2(new_n609), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT35), .B(G107), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(KEYINPUT100), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n634), .B(new_n636), .ZN(G9));
  NAND2_X1  g451(.A1(new_n604), .A2(new_n548), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n532), .A2(KEYINPUT36), .ZN(new_n639));
  OR2_X1    g453(.A1(new_n531), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n531), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n640), .A2(new_n544), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT101), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n542), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n638), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n507), .A2(new_n646), .A3(new_n608), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT37), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(new_n519), .ZN(G12));
  NOR2_X1   g463(.A1(new_n322), .A2(G900), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT102), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n320), .B(KEYINPUT103), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n632), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n595), .A2(new_n654), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n644), .B(new_n317), .C1(new_n392), .C2(new_n393), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n316), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G128), .ZN(G30));
  XOR2_X1   g473(.A(new_n653), .B(KEYINPUT39), .Z(new_n660));
  NAND2_X1  g474(.A1(new_n595), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT105), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT40), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT104), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n272), .B1(new_n264), .B2(new_n266), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n285), .A2(new_n286), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n668), .A2(new_n272), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n666), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n295), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n667), .A2(new_n666), .A3(new_n669), .ZN(new_n672));
  OAI21_X1  g486(.A(G472), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n673), .B1(new_n312), .B2(new_n315), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n645), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n374), .ZN(new_n677));
  INV_X1    g491(.A(new_n332), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n330), .B(new_n678), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n335), .B1(new_n369), .B2(new_n370), .ZN(new_n680));
  INV_X1    g494(.A(new_n365), .ZN(new_n681));
  OAI21_X1  g495(.A(KEYINPUT6), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n364), .A2(new_n334), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n679), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n390), .ZN(new_n685));
  AOI21_X1  g499(.A(KEYINPUT87), .B1(new_n386), .B2(new_n295), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n677), .B1(new_n684), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n373), .A2(new_n374), .A3(new_n391), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT38), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(KEYINPUT38), .B1(new_n688), .B2(new_n689), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n610), .A2(new_n482), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n665), .A2(new_n317), .A3(new_n676), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G143), .ZN(G45));
  INV_X1    g513(.A(new_n317), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n700), .B1(new_n688), .B2(new_n689), .ZN(new_n701));
  INV_X1    g515(.A(new_n653), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n610), .A2(new_n622), .A3(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n316), .A2(new_n646), .A3(new_n701), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT106), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(new_n211), .ZN(G48));
  AOI21_X1  g521(.A(KEYINPUT83), .B1(new_n562), .B2(new_n566), .ZN(new_n708));
  AOI211_X1 g522(.A(new_n568), .B(new_n571), .C1(new_n559), .C2(new_n561), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n708), .A2(new_n709), .A3(new_n583), .ZN(new_n710));
  OAI21_X1  g524(.A(G469), .B1(new_n710), .B2(G902), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n711), .A2(new_n548), .A3(new_n587), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(KEYINPUT107), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT107), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n711), .A2(new_n714), .A3(new_n548), .A4(new_n587), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n716), .A2(new_n316), .A3(new_n546), .A4(new_n624), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT41), .B(G113), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G15));
  NAND4_X1  g533(.A1(new_n716), .A2(new_n316), .A3(new_n546), .A4(new_n633), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G116), .ZN(G18));
  NOR2_X1   g535(.A1(new_n645), .A2(new_n506), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n317), .B1(new_n392), .B2(new_n393), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n712), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n316), .A2(new_n722), .A3(new_n323), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(KEYINPUT108), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(new_n188), .ZN(G21));
  OAI21_X1  g541(.A(KEYINPUT109), .B1(new_n723), .B2(new_n696), .ZN(new_n728));
  INV_X1    g542(.A(new_n443), .ZN(new_n729));
  INV_X1    g543(.A(new_n505), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n629), .B1(new_n628), .B2(new_n484), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n630), .B1(new_n731), .B2(new_n504), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n729), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n483), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT109), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n701), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n728), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n272), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n301), .A2(new_n308), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n310), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n542), .A2(new_n545), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n742), .A2(new_n601), .A3(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n323), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n745), .B1(new_n713), .B2(new_n715), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n737), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G122), .ZN(G24));
  NOR3_X1   g562(.A1(new_n742), .A2(new_n645), .A3(new_n601), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(new_n724), .A3(new_n704), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G125), .ZN(G27));
  XNOR2_X1  g565(.A(new_n311), .B(new_n314), .ZN(new_n752));
  INV_X1    g566(.A(new_n297), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n546), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n688), .A2(new_n317), .A3(new_n689), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n704), .A2(new_n756), .A3(new_n595), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT42), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n638), .A2(new_n703), .A3(KEYINPUT42), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n759), .A2(new_n316), .A3(new_n546), .A4(new_n756), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(new_n229), .ZN(G33));
  INV_X1    g576(.A(new_n655), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n316), .A2(new_n763), .A3(new_n546), .A4(new_n756), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G134), .ZN(G36));
  OAI211_X1 g579(.A(new_n443), .B(new_n622), .C1(new_n503), .C2(new_n505), .ZN(new_n766));
  AOI211_X1 g580(.A(KEYINPUT111), .B(KEYINPUT43), .C1(new_n766), .C2(KEYINPUT110), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n620), .B1(new_n618), .B2(G478), .ZN(new_n769));
  AOI211_X1 g583(.A(new_n729), .B(new_n769), .C1(new_n730), .C2(new_n732), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT110), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n768), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT43), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n773), .B1(new_n766), .B2(KEYINPUT111), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n767), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(new_n603), .A3(new_n644), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT44), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(KEYINPUT112), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT112), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n776), .A2(new_n780), .A3(new_n777), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n775), .A2(KEYINPUT44), .A3(new_n603), .A4(new_n644), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT45), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n784), .B1(new_n590), .B2(new_n592), .ZN(new_n785));
  INV_X1    g599(.A(new_n561), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n786), .B1(new_n582), .B2(new_n578), .ZN(new_n787));
  OAI211_X1 g601(.A(KEYINPUT45), .B(new_n591), .C1(new_n787), .C2(new_n571), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n785), .A2(G469), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n588), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT46), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n789), .A2(KEYINPUT46), .A3(new_n790), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n793), .A2(new_n587), .A3(new_n794), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n795), .A2(new_n548), .A3(new_n660), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n783), .A2(new_n756), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n782), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G137), .ZN(G39));
  NAND2_X1  g613(.A1(new_n795), .A2(new_n548), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT47), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n795), .A2(KEYINPUT47), .A3(new_n548), .ZN(new_n803));
  AOI211_X1 g617(.A(new_n703), .B(new_n755), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n316), .A2(new_n546), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G140), .ZN(G42));
  AND2_X1   g622(.A1(new_n711), .A2(new_n587), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT49), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n695), .A2(new_n810), .A3(new_n546), .A4(new_n317), .ZN(new_n811));
  OR4_X1    g625(.A1(new_n549), .A2(new_n811), .A3(new_n674), .A4(new_n766), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n771), .B1(new_n733), .B2(new_n622), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n774), .B1(new_n813), .B2(KEYINPUT111), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n768), .B(new_n773), .C1(new_n770), .C2(new_n771), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n814), .A2(new_n652), .A3(new_n744), .A4(new_n815), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n816), .A2(new_n723), .A3(new_n712), .ZN(new_n817));
  INV_X1    g631(.A(new_n754), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n712), .A2(new_n755), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n818), .A2(new_n652), .A3(new_n775), .A4(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(KEYINPUT48), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n674), .A2(new_n712), .A3(new_n755), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n743), .A2(new_n320), .ZN(new_n823));
  AND4_X1   g637(.A1(new_n610), .A2(new_n822), .A3(new_n622), .A4(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(G952), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n824), .A2(new_n825), .A3(G953), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT50), .ZN(new_n827));
  INV_X1    g641(.A(new_n712), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n775), .A2(new_n652), .A3(new_n828), .A4(new_n744), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n700), .B1(new_n692), .B2(new_n693), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n827), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n816), .A2(new_n712), .ZN(new_n832));
  INV_X1    g646(.A(new_n830), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n832), .A2(KEYINPUT50), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n809), .A2(new_n549), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n802), .A2(new_n803), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n816), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n837), .A2(new_n756), .A3(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n775), .A2(new_n652), .A3(new_n749), .A4(new_n819), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n822), .A2(new_n733), .A3(new_n769), .A4(new_n823), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n835), .A2(new_n839), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT50), .B1(new_n832), .B2(new_n833), .ZN(new_n844));
  NOR4_X1   g658(.A1(new_n816), .A2(new_n827), .A3(new_n830), .A4(new_n712), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n839), .B(new_n843), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n842), .B1(KEYINPUT51), .B2(new_n846), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n839), .B(new_n840), .C1(new_n844), .C2(new_n845), .ZN(new_n848));
  INV_X1    g662(.A(new_n841), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n846), .A2(KEYINPUT51), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n821), .B(new_n826), .C1(new_n847), .C2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT53), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n638), .A2(new_n653), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n723), .A2(new_n696), .A3(KEYINPUT109), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n735), .B1(new_n701), .B2(new_n734), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n858), .A2(new_n675), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n705), .A2(new_n658), .A3(new_n750), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT52), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n747), .A2(new_n717), .A3(new_n720), .A4(new_n725), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n758), .A2(new_n760), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n737), .A2(new_n645), .A3(new_n674), .A4(new_n855), .ZN(new_n865));
  NOR4_X1   g679(.A1(new_n703), .A2(new_n742), .A3(new_n645), .A4(new_n601), .ZN(new_n866));
  AOI22_X1  g680(.A1(new_n866), .A2(new_n724), .B1(new_n657), .B2(new_n316), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT52), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n865), .A2(new_n867), .A3(new_n868), .A4(new_n705), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n861), .A2(new_n863), .A3(new_n864), .A4(new_n869), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n506), .B(KEYINPUT113), .C1(new_n733), .C2(new_n622), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT113), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n872), .B1(new_n733), .B2(new_n769), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n394), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n606), .A2(new_n874), .A3(new_n609), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n875), .A2(new_n596), .A3(new_n647), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT115), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n483), .B(new_n443), .C1(new_n731), .C2(new_n499), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT114), .B1(new_n878), .B2(new_n653), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT114), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n631), .A2(new_n880), .A3(new_n483), .A4(new_n702), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n877), .B1(new_n882), .B2(new_n755), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n879), .A2(new_n881), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n392), .A2(new_n393), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n884), .A2(new_n885), .A3(KEYINPUT115), .A4(new_n317), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n883), .A2(new_n316), .A3(new_n646), .A4(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n749), .A2(new_n595), .A3(new_n704), .A4(new_n756), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n887), .A2(new_n764), .A3(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n876), .A2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n854), .B1(new_n870), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n854), .B1(new_n890), .B2(KEYINPUT116), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n859), .A2(new_n860), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n862), .B1(new_n894), .B2(new_n868), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n865), .A2(new_n867), .A3(new_n705), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n761), .B1(new_n896), .B2(KEYINPUT52), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT116), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n898), .B1(new_n876), .B2(new_n889), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n893), .A2(new_n895), .A3(new_n897), .A4(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT54), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n892), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n895), .A2(KEYINPUT53), .A3(new_n897), .A4(new_n890), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n901), .B1(new_n892), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(KEYINPUT117), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n892), .A2(new_n903), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT54), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT117), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n892), .A2(new_n900), .A3(new_n901), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AOI211_X1 g724(.A(new_n817), .B(new_n853), .C1(new_n905), .C2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(G952), .A2(G953), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n812), .B1(new_n911), .B2(new_n912), .ZN(G75));
  NOR2_X1   g727(.A1(new_n366), .A2(new_n372), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(new_n333), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT119), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n295), .B1(new_n892), .B2(new_n900), .ZN(new_n917));
  AOI211_X1 g731(.A(KEYINPUT55), .B(KEYINPUT56), .C1(new_n917), .C2(G210), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT55), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n892), .A2(new_n900), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n920), .A2(G210), .A3(G902), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT56), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n919), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n916), .B1(new_n918), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n319), .A2(G952), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(G210), .ZN(new_n927));
  AOI211_X1 g741(.A(new_n927), .B(new_n295), .C1(new_n892), .C2(new_n900), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT55), .B1(new_n928), .B2(KEYINPUT56), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n921), .A2(new_n919), .A3(new_n922), .ZN(new_n930));
  INV_X1    g744(.A(new_n916), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n924), .A2(new_n926), .A3(new_n932), .ZN(G51));
  NAND2_X1  g747(.A1(new_n920), .A2(KEYINPUT54), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n909), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n790), .A2(KEYINPUT57), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n790), .A2(KEYINPUT57), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n585), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n917), .A2(G469), .A3(new_n785), .A4(new_n788), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n925), .B1(new_n939), .B2(new_n940), .ZN(G54));
  NAND3_X1  g755(.A1(new_n917), .A2(KEYINPUT58), .A3(G475), .ZN(new_n942));
  INV_X1    g756(.A(new_n628), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n942), .A2(new_n943), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n944), .A2(new_n945), .A3(new_n925), .ZN(G60));
  NAND2_X1  g760(.A1(G478), .A2(G902), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT59), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n616), .A2(new_n617), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n949), .B1(new_n934), .B2(new_n909), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n905), .A2(new_n910), .A3(new_n948), .ZN(new_n951));
  AOI221_X4 g765(.A(new_n925), .B1(new_n948), .B2(new_n950), .C1(new_n951), .C2(new_n949), .ZN(G63));
  NAND2_X1  g766(.A1(G217), .A2(G902), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT60), .Z(new_n954));
  NAND4_X1  g768(.A1(new_n920), .A2(new_n641), .A3(new_n640), .A4(new_n954), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n920), .A2(new_n954), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n926), .B(new_n955), .C1(new_n956), .C2(new_n536), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT61), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n957), .B(new_n958), .ZN(G66));
  INV_X1    g773(.A(new_n321), .ZN(new_n960));
  OAI21_X1  g774(.A(G953), .B1(new_n960), .B2(new_n331), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n862), .A2(new_n876), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n961), .B1(new_n962), .B2(G953), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n914), .B1(G898), .B2(new_n319), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n963), .B(new_n964), .ZN(G69));
  NAND2_X1  g779(.A1(new_n871), .A2(new_n873), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n966), .A2(KEYINPUT122), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n663), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n316), .A2(new_n546), .A3(new_n756), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n966), .A2(KEYINPUT122), .ZN(new_n971));
  OAI21_X1  g785(.A(KEYINPUT123), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OR4_X1    g786(.A1(KEYINPUT123), .A2(new_n968), .A3(new_n969), .A4(new_n971), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT62), .ZN(new_n974));
  AOI22_X1  g788(.A1(new_n972), .A2(new_n973), .B1(KEYINPUT121), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n860), .B(KEYINPUT120), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n698), .A2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT121), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n977), .A2(new_n978), .A3(KEYINPUT62), .ZN(new_n979));
  AOI22_X1  g793(.A1(new_n782), .A2(new_n797), .B1(new_n806), .B2(new_n804), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n698), .B(new_n976), .C1(KEYINPUT121), .C2(new_n974), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n975), .A2(new_n979), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n319), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n299), .B(new_n492), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n319), .B1(G227), .B2(G900), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n983), .A2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(G900), .ZN(new_n988));
  OAI21_X1  g802(.A(G953), .B1(new_n988), .B2(G227), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n758), .A2(new_n760), .A3(new_n764), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT124), .Z(new_n991));
  NAND3_X1  g805(.A1(new_n818), .A2(new_n737), .A3(new_n796), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n976), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n980), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n984), .B(new_n989), .C1(new_n994), .C2(G953), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n987), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(KEYINPUT125), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT125), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n987), .A2(new_n995), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n997), .A2(new_n999), .ZN(G72));
  AOI211_X1 g814(.A(new_n273), .B(new_n667), .C1(new_n892), .C2(new_n903), .ZN(new_n1001));
  XNOR2_X1  g815(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n600), .A2(new_n295), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1002), .B(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n962), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1004), .B1(new_n982), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(new_n667), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT127), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n980), .A2(new_n991), .A3(new_n993), .A4(new_n962), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(new_n1004), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(new_n273), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1009), .B1(new_n1012), .B2(new_n926), .ZN(new_n1013));
  AOI211_X1 g827(.A(KEYINPUT127), .B(new_n925), .C1(new_n1011), .C2(new_n273), .ZN(new_n1014));
  OAI211_X1 g828(.A(new_n1005), .B(new_n1008), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1015), .ZN(G57));
endmodule


