//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988;
  INV_X1    g000(.A(G210), .ZN(new_n187));
  NOR3_X1   g001(.A1(new_n187), .A2(G237), .A3(G953), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT27), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT26), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(G101), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT28), .ZN(new_n192));
  XNOR2_X1  g006(.A(G116), .B(G119), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT2), .B(G113), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n193), .B(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(G146), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(G143), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT0), .B(G128), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT11), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(G137), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(G137), .ZN(new_n207));
  INV_X1    g021(.A(G137), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(KEYINPUT11), .A3(G134), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n206), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G131), .ZN(new_n211));
  INV_X1    g025(.A(G131), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n206), .A2(new_n209), .A3(new_n212), .A4(new_n207), .ZN(new_n213));
  NAND2_X1  g027(.A1(KEYINPUT0), .A2(G128), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n199), .A2(KEYINPUT64), .A3(G143), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT64), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n217), .B1(new_n197), .B2(G146), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n215), .B(new_n216), .C1(new_n218), .C2(new_n198), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT65), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT64), .B1(new_n199), .B2(G143), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n199), .A2(G143), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n223), .A2(new_n224), .A3(new_n215), .A4(new_n216), .ZN(new_n225));
  AOI221_X4 g039(.A(new_n203), .B1(new_n211), .B2(new_n213), .C1(new_n220), .C2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT1), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n223), .A2(new_n227), .A3(G128), .A4(new_n216), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT1), .B1(new_n197), .B2(G146), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G128), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n230), .B1(new_n198), .B2(new_n200), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n207), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n205), .A2(G137), .ZN(new_n234));
  OAI21_X1  g048(.A(G131), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n235), .A2(new_n213), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n232), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n196), .B1(new_n226), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n220), .A2(new_n225), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n211), .A2(new_n213), .ZN(new_n241));
  INV_X1    g055(.A(new_n203), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(new_n195), .A3(new_n237), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n192), .B1(new_n239), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n192), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n191), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT31), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n243), .A2(new_n195), .A3(new_n237), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT30), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n203), .B1(new_n220), .B2(new_n225), .ZN(new_n252));
  AOI221_X4 g066(.A(new_n251), .B1(new_n232), .B2(new_n236), .C1(new_n252), .C2(new_n241), .ZN(new_n253));
  AOI21_X1  g067(.A(KEYINPUT30), .B1(new_n243), .B2(new_n237), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n250), .B1(new_n255), .B2(new_n196), .ZN(new_n256));
  INV_X1    g070(.A(G101), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n190), .B(new_n257), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n248), .A2(new_n249), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NOR3_X1   g073(.A1(new_n253), .A2(new_n254), .A3(new_n195), .ZN(new_n260));
  NOR4_X1   g074(.A1(new_n260), .A2(KEYINPUT31), .A3(new_n191), .A4(new_n250), .ZN(new_n261));
  OAI21_X1  g075(.A(KEYINPUT66), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(G472), .A2(G902), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT66), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n256), .A2(new_n249), .A3(new_n258), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n195), .B1(new_n243), .B2(new_n237), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT28), .B1(new_n250), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n246), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT31), .B1(new_n268), .B2(new_n191), .ZN(new_n269));
  AOI211_X1 g083(.A(new_n250), .B(new_n191), .C1(new_n255), .C2(new_n196), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n264), .B(new_n265), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n262), .A2(new_n263), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT32), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n262), .A2(new_n271), .A3(KEYINPUT32), .A4(new_n263), .ZN(new_n275));
  INV_X1    g089(.A(G902), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n268), .A2(new_n191), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT29), .ZN(new_n278));
  OR2_X1    g092(.A1(new_n277), .A2(KEYINPUT29), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n256), .A2(new_n258), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n276), .B(new_n278), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G472), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n274), .A2(new_n275), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G217), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n284), .B1(G234), .B2(new_n276), .ZN(new_n285));
  INV_X1    g099(.A(G128), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT67), .B1(new_n286), .B2(G119), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT67), .ZN(new_n288));
  INV_X1    g102(.A(G119), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n289), .A3(G128), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n289), .A2(G128), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  XOR2_X1   g108(.A(KEYINPUT24), .B(G110), .Z(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n294), .A2(KEYINPUT69), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT69), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n292), .B1(new_n287), .B2(new_n290), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n298), .B1(new_n299), .B2(new_n295), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT23), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n292), .A2(new_n301), .ZN(new_n302));
  NOR3_X1   g116(.A1(new_n289), .A2(KEYINPUT23), .A3(G128), .ZN(new_n303));
  OAI22_X1  g117(.A1(new_n302), .A2(new_n303), .B1(G119), .B2(new_n286), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n297), .B(new_n300), .C1(G110), .C2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G140), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G125), .ZN(new_n307));
  INV_X1    g121(.A(G125), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G140), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT16), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT68), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n312), .B1(new_n307), .B2(KEYINPUT16), .ZN(new_n313));
  OR3_X1    g127(.A1(new_n307), .A2(new_n312), .A3(KEYINPUT16), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n311), .A2(G146), .A3(new_n313), .A4(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n310), .A2(new_n199), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n305), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT70), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n311), .A2(new_n313), .A3(new_n314), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n199), .ZN(new_n321));
  AOI22_X1  g135(.A1(new_n321), .A2(new_n315), .B1(new_n295), .B2(new_n299), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n304), .A2(G110), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n305), .A2(KEYINPUT70), .A3(new_n315), .A4(new_n316), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n319), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT72), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n319), .A2(new_n324), .A3(KEYINPUT72), .A4(new_n325), .ZN(new_n329));
  INV_X1    g143(.A(G953), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(G221), .A3(G234), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(KEYINPUT71), .ZN(new_n332));
  XOR2_X1   g146(.A(new_n332), .B(KEYINPUT22), .Z(new_n333));
  XNOR2_X1  g147(.A(new_n333), .B(new_n208), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n328), .A2(new_n329), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n326), .A2(new_n327), .A3(new_n334), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(KEYINPUT25), .B1(new_n338), .B2(new_n276), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT25), .ZN(new_n340));
  AOI211_X1 g154(.A(new_n340), .B(G902), .C1(new_n336), .C2(new_n337), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n285), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n285), .A2(G902), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT9), .B(G234), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(KEYINPUT73), .ZN(new_n347));
  OAI21_X1  g161(.A(G221), .B1(new_n347), .B2(G902), .ZN(new_n348));
  INV_X1    g162(.A(G469), .ZN(new_n349));
  INV_X1    g163(.A(G104), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT3), .B1(new_n350), .B2(G107), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT3), .ZN(new_n352));
  INV_X1    g166(.A(G107), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n352), .A2(new_n353), .A3(G104), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n350), .A2(G107), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n351), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT4), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n357), .A3(G101), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n351), .A2(new_n354), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT74), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n360), .A2(new_n361), .A3(new_n257), .A4(new_n355), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n351), .A2(new_n354), .A3(new_n257), .A4(new_n355), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT74), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n357), .B1(new_n356), .B2(G101), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n359), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n353), .A2(G104), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n257), .B1(new_n355), .B2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n369), .B1(new_n362), .B2(new_n364), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n371), .B1(new_n228), .B2(new_n231), .ZN(new_n372));
  AOI22_X1  g186(.A1(new_n367), .A2(new_n252), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n369), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n363), .A2(KEYINPUT74), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n363), .A2(KEYINPUT74), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI211_X1 g191(.A(G128), .B(new_n216), .C1(new_n218), .C2(new_n198), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n229), .A2(KEYINPUT75), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT75), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n222), .A2(new_n381), .A3(KEYINPUT1), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n380), .A2(G128), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n223), .A2(new_n216), .ZN(new_n384));
  AOI22_X1  g198(.A1(new_n379), .A2(new_n227), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n371), .B1(new_n377), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n373), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n241), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n366), .B1(new_n375), .B2(new_n376), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(new_n252), .A3(new_n358), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n370), .A2(new_n372), .ZN(new_n391));
  INV_X1    g205(.A(new_n241), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n386), .A2(new_n390), .A3(new_n391), .A4(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(G110), .B(G140), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n330), .A2(G227), .ZN(new_n395));
  XOR2_X1   g209(.A(new_n394), .B(new_n395), .Z(new_n396));
  NAND3_X1  g210(.A1(new_n388), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n396), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT12), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n377), .A2(new_n385), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n370), .A2(new_n232), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n399), .B(new_n241), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n393), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n383), .A2(new_n384), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n228), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n370), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n406), .B1(new_n232), .B2(new_n370), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n399), .B1(new_n407), .B2(new_n241), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n398), .B1(new_n403), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n397), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n349), .B1(new_n410), .B2(new_n276), .ZN(new_n411));
  XNOR2_X1  g225(.A(KEYINPUT76), .B(G469), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n392), .B1(new_n373), .B2(new_n386), .ZN(new_n413));
  INV_X1    g227(.A(new_n393), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n398), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n241), .B1(new_n400), .B2(new_n401), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT12), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n417), .A2(new_n393), .A3(new_n402), .A4(new_n396), .ZN(new_n418));
  AOI211_X1 g232(.A(G902), .B(new_n412), .C1(new_n415), .C2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n348), .B1(new_n411), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  XOR2_X1   g235(.A(G113), .B(G122), .Z(new_n422));
  XNOR2_X1  g236(.A(new_n422), .B(KEYINPUT85), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n423), .B(new_n350), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n307), .A2(new_n309), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT80), .B1(new_n425), .B2(G146), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(G146), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n425), .A2(KEYINPUT80), .A3(G146), .ZN(new_n429));
  NOR2_X1   g243(.A1(G237), .A2(G953), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G214), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n197), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n430), .A2(G143), .A3(G214), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n212), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AOI22_X1  g248(.A1(new_n428), .A2(new_n429), .B1(new_n434), .B2(KEYINPUT18), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT18), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n432), .B(new_n433), .C1(new_n436), .C2(new_n212), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT81), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n437), .A2(new_n438), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n435), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n434), .A2(KEYINPUT17), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT86), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n442), .B(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n433), .ZN(new_n445));
  AOI21_X1  g259(.A(G143), .B1(new_n430), .B2(G214), .ZN(new_n446));
  OAI21_X1  g260(.A(G131), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n432), .A2(new_n212), .A3(new_n433), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n321), .B(new_n315), .C1(new_n449), .C2(KEYINPUT17), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n424), .B(new_n441), .C1(new_n444), .C2(new_n450), .ZN(new_n451));
  NOR3_X1   g265(.A1(new_n445), .A2(new_n446), .A3(G131), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT82), .B1(new_n452), .B2(new_n434), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT19), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n310), .A2(KEYINPUT83), .A3(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT83), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n456), .B1(new_n425), .B2(KEYINPUT19), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n425), .A2(KEYINPUT19), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n455), .A2(new_n457), .A3(new_n199), .A4(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT82), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n447), .A2(new_n448), .A3(new_n460), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n453), .A2(new_n315), .A3(new_n459), .A4(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n441), .A2(new_n462), .A3(KEYINPUT84), .ZN(new_n463));
  INV_X1    g277(.A(new_n424), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(KEYINPUT84), .B1(new_n441), .B2(new_n462), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n451), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT20), .ZN(new_n468));
  NOR2_X1   g282(.A1(G475), .A2(G902), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n469), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n467), .A2(KEYINPUT87), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT87), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n473), .B(new_n451), .C1(new_n465), .C2(new_n466), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n471), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n470), .B1(new_n475), .B2(new_n468), .ZN(new_n476));
  INV_X1    g290(.A(G122), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(G116), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT88), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n478), .B(new_n479), .ZN(new_n480));
  OR2_X1    g294(.A1(new_n477), .A2(G116), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  OR2_X1    g297(.A1(new_n353), .A2(KEYINPUT14), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n353), .B1(new_n480), .B2(new_n481), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n480), .A2(KEYINPUT14), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(G128), .B(G143), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(new_n205), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n485), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(KEYINPUT13), .B1(new_n286), .B2(G143), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n492), .A2(new_n205), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(new_n489), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n480), .A2(new_n353), .A3(new_n481), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n494), .B1(new_n496), .B2(new_n486), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n491), .A2(new_n497), .ZN(new_n498));
  NOR3_X1   g312(.A1(new_n347), .A2(new_n284), .A3(G953), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n491), .A2(new_n497), .A3(new_n499), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n276), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT15), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(G478), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n504), .B(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n441), .B1(new_n444), .B2(new_n450), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n464), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n451), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n276), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n511), .A2(G475), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n476), .A2(new_n507), .A3(new_n513), .ZN(new_n514));
  XOR2_X1   g328(.A(G110), .B(G122), .Z(new_n515));
  AOI211_X1 g329(.A(new_n195), .B(new_n359), .C1(new_n365), .C2(new_n366), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT5), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n517), .A2(new_n289), .A3(G116), .ZN(new_n518));
  INV_X1    g332(.A(new_n193), .ZN(new_n519));
  OAI211_X1 g333(.A(G113), .B(new_n518), .C1(new_n519), .C2(new_n517), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n520), .B1(new_n519), .B2(new_n194), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n377), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n515), .B1(new_n516), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(KEYINPUT77), .B1(new_n523), .B2(KEYINPUT6), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n367), .A2(new_n196), .ZN(new_n525));
  OR2_X1    g339(.A1(new_n377), .A2(new_n521), .ZN(new_n526));
  INV_X1    g340(.A(new_n515), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n523), .A2(new_n528), .A3(KEYINPUT6), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n228), .A2(new_n231), .A3(new_n308), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n531), .B1(new_n252), .B2(new_n308), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT78), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT78), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n534), .B1(new_n252), .B2(new_n308), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(G224), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(G953), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n538), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n533), .A2(new_n540), .A3(new_n535), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n523), .A2(new_n528), .A3(KEYINPUT77), .A4(KEYINPUT6), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n530), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n533), .A2(KEYINPUT7), .A3(new_n540), .A4(new_n535), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT7), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n532), .B1(new_n546), .B2(new_n538), .ZN(new_n547));
  XOR2_X1   g361(.A(new_n515), .B(KEYINPUT8), .Z(new_n548));
  AND2_X1   g362(.A1(new_n377), .A2(new_n521), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n548), .B1(new_n549), .B2(new_n522), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n545), .A2(new_n528), .A3(new_n547), .A4(new_n550), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n551), .A2(new_n276), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n544), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(G210), .B1(G237), .B2(G902), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT79), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n556), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n544), .A2(new_n552), .A3(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(G214), .B1(G237), .B2(G902), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  XOR2_X1   g375(.A(KEYINPUT21), .B(G898), .Z(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(G234), .A2(G237), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n564), .A2(G902), .A3(G953), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n330), .A2(G952), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n567), .A2(new_n564), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n561), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n557), .A2(new_n559), .A3(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n514), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n283), .A2(new_n345), .A3(new_n421), .A4(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(G101), .ZN(G3));
  INV_X1    g388(.A(new_n345), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n262), .A2(new_n276), .A3(new_n271), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(G472), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n272), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n575), .A2(new_n420), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(G478), .B1(new_n503), .B2(new_n276), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT90), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n483), .A2(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n582));
  INV_X1    g396(.A(new_n486), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n495), .ZN(new_n584));
  AOI22_X1  g398(.A1(new_n582), .A2(new_n490), .B1(new_n584), .B2(new_n494), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n581), .B1(new_n585), .B2(new_n499), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n503), .A2(KEYINPUT33), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT33), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n501), .B(new_n502), .C1(new_n581), .C2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(G902), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n580), .B1(new_n590), .B2(G478), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n470), .ZN(new_n593));
  INV_X1    g407(.A(new_n474), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n441), .A2(new_n462), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT84), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n597), .A2(new_n464), .A3(new_n463), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n473), .B1(new_n598), .B2(new_n451), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n469), .B1(new_n594), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n593), .B1(new_n600), .B2(KEYINPUT20), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n592), .B1(new_n601), .B2(new_n512), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n553), .A2(KEYINPUT89), .A3(new_n554), .ZN(new_n603));
  OR2_X1    g417(.A1(new_n554), .A2(KEYINPUT89), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n554), .A2(KEYINPUT89), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n544), .A2(new_n552), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n603), .A2(new_n570), .A3(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n579), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT34), .B(G104), .Z(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G6));
  INV_X1    g425(.A(new_n507), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n472), .A2(new_n474), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n468), .B1(new_n613), .B2(new_n469), .ZN(new_n614));
  AOI211_X1 g428(.A(KEYINPUT20), .B(new_n471), .C1(new_n472), .C2(new_n474), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n612), .B(new_n513), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n616), .A2(new_n607), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n579), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT35), .B(G107), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G9));
  AND2_X1   g434(.A1(new_n262), .A2(new_n271), .ZN(new_n621));
  AOI22_X1  g435(.A1(new_n621), .A2(new_n263), .B1(new_n576), .B2(G472), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n335), .A2(KEYINPUT36), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(new_n326), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n343), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n420), .B1(new_n342), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n622), .A2(new_n572), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT91), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT37), .B(G110), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G12));
  NAND2_X1  g444(.A1(new_n603), .A2(new_n606), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n631), .A2(new_n561), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n283), .A2(new_n626), .A3(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT92), .ZN(new_n634));
  INV_X1    g448(.A(G900), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n568), .B1(new_n565), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n634), .B1(new_n616), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n600), .A2(KEYINPUT20), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n475), .A2(new_n468), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n507), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n636), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n640), .A2(KEYINPUT92), .A3(new_n513), .A4(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n633), .A2(new_n644), .A3(KEYINPUT93), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT93), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n283), .A2(new_n626), .A3(new_n632), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n646), .B1(new_n647), .B2(new_n643), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G128), .ZN(G30));
  AND3_X1   g464(.A1(new_n544), .A2(new_n552), .A3(new_n558), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n558), .B1(new_n544), .B2(new_n552), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(new_n653), .B(KEYINPUT38), .Z(new_n654));
  NOR2_X1   g468(.A1(new_n256), .A2(new_n191), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n239), .A2(new_n244), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n276), .B1(new_n656), .B2(new_n258), .ZN(new_n657));
  OAI21_X1  g471(.A(G472), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n274), .A2(new_n275), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n342), .A2(new_n625), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n476), .A2(new_n513), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n663), .A2(new_n612), .A3(new_n560), .ZN(new_n664));
  OR4_X1    g478(.A1(KEYINPUT94), .A2(new_n654), .A3(new_n662), .A4(new_n664), .ZN(new_n665));
  OR2_X1    g479(.A1(new_n654), .A2(new_n664), .ZN(new_n666));
  OAI21_X1  g480(.A(KEYINPUT94), .B1(new_n666), .B2(new_n662), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n636), .B(KEYINPUT39), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n421), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n670), .B(KEYINPUT40), .Z(new_n671));
  NAND3_X1  g485(.A1(new_n665), .A2(new_n667), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G143), .ZN(G45));
  AOI211_X1 g487(.A(new_n636), .B(new_n591), .C1(new_n476), .C2(new_n513), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n283), .A2(new_n626), .A3(new_n632), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G146), .ZN(G48));
  AOI21_X1  g490(.A(G902), .B1(new_n415), .B2(new_n418), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n677), .A2(new_n349), .ZN(new_n678));
  INV_X1    g492(.A(new_n412), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n678), .A2(new_n348), .A3(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n283), .A2(new_n608), .A3(new_n345), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT41), .B(G113), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G15));
  NAND4_X1  g499(.A1(new_n283), .A2(new_n617), .A3(new_n345), .A4(new_n682), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G116), .ZN(G18));
  INV_X1    g501(.A(new_n607), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n514), .A2(new_n681), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n283), .A2(new_n688), .A3(new_n660), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G119), .ZN(G21));
  OAI21_X1  g505(.A(new_n612), .B1(new_n601), .B2(new_n512), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n692), .A2(new_n607), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n265), .B1(new_n269), .B2(new_n270), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n694), .A2(new_n263), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n695), .B1(new_n576), .B2(G472), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n693), .A2(new_n345), .A3(new_n682), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G122), .ZN(G24));
  NOR3_X1   g512(.A1(new_n631), .A2(new_n681), .A3(new_n561), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n699), .A2(new_n660), .A3(new_n674), .A4(new_n696), .ZN(new_n700));
  XOR2_X1   g514(.A(KEYINPUT95), .B(G125), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G27));
  INV_X1    g516(.A(KEYINPUT97), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n349), .A2(new_n276), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n704), .B1(new_n677), .B2(new_n679), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n409), .A2(KEYINPUT96), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT96), .ZN(new_n707));
  OAI211_X1 g521(.A(new_n707), .B(new_n398), .C1(new_n403), .C2(new_n408), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n706), .A2(G469), .A3(new_n397), .A4(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n703), .B1(new_n710), .B2(new_n348), .ZN(new_n711));
  INV_X1    g525(.A(new_n348), .ZN(new_n712));
  AOI211_X1 g526(.A(KEYINPUT97), .B(new_n712), .C1(new_n705), .C2(new_n709), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n560), .B1(new_n651), .B2(new_n652), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n711), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n715), .A2(new_n283), .A3(new_n345), .A4(new_n674), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT42), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n283), .A2(new_n345), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n719), .A2(KEYINPUT42), .A3(new_n674), .A4(new_n715), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G131), .ZN(G33));
  AOI21_X1  g536(.A(KEYINPUT98), .B1(new_n637), .B2(new_n642), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n283), .A2(new_n345), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n710), .A2(new_n348), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT97), .ZN(new_n726));
  INV_X1    g540(.A(new_n714), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n710), .A2(new_n703), .A3(new_n348), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n723), .A2(new_n724), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n644), .A2(KEYINPUT98), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G134), .ZN(G36));
  NAND4_X1  g547(.A1(new_n706), .A2(KEYINPUT45), .A3(new_n397), .A4(new_n708), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT45), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n410), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n734), .A2(G469), .A3(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n704), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(KEYINPUT46), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n680), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n348), .ZN(new_n742));
  OAI21_X1  g556(.A(KEYINPUT99), .B1(new_n742), .B2(new_n668), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT99), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n741), .A2(new_n744), .A3(new_n348), .A4(new_n669), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT101), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n592), .A2(new_n476), .A3(new_n747), .A4(new_n513), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT100), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT43), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n663), .A2(new_n592), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT101), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n749), .B(KEYINPUT43), .C1(new_n663), .C2(new_n591), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n752), .A2(new_n578), .A3(new_n754), .A4(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT44), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n756), .A2(new_n757), .A3(new_n661), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n746), .A2(new_n758), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n756), .A2(new_n661), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n714), .B1(new_n760), .B2(new_n757), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G137), .ZN(G39));
  NOR2_X1   g577(.A1(new_n283), .A2(new_n345), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n742), .A2(KEYINPUT47), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT47), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n741), .A2(new_n766), .A3(new_n348), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n602), .A2(new_n636), .A3(new_n714), .ZN(new_n768));
  AND4_X1   g582(.A1(new_n764), .A2(new_n765), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(new_n306), .ZN(G42));
  NOR2_X1   g584(.A1(G952), .A2(G953), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n752), .A2(new_n755), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n772), .A2(new_n754), .ZN(new_n773));
  INV_X1    g587(.A(new_n696), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n575), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n773), .A2(new_n568), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n765), .A2(new_n767), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n678), .A2(new_n680), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT103), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n779), .A2(KEYINPUT108), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(KEYINPUT108), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(new_n712), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n776), .B1(new_n777), .B2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n659), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n714), .A2(new_n681), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n784), .A2(new_n345), .A3(new_n568), .A4(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT112), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n753), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n787), .A2(KEYINPUT113), .A3(new_n753), .ZN(new_n791));
  AOI22_X1  g605(.A1(new_n783), .A2(new_n727), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n773), .A2(new_n568), .A3(new_n785), .ZN(new_n793));
  OR3_X1    g607(.A1(new_n793), .A2(new_n661), .A3(new_n774), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(KEYINPUT111), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n773), .A2(new_n568), .A3(new_n775), .A4(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT111), .B1(new_n795), .B2(KEYINPUT110), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n654), .A2(new_n561), .A3(new_n682), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT109), .ZN(new_n801));
  OR3_X1    g615(.A1(new_n797), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n799), .B1(new_n797), .B2(new_n801), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n792), .A2(new_n794), .A3(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n699), .ZN(new_n808));
  OAI21_X1  g622(.A(KEYINPUT114), .B1(new_n793), .B2(new_n724), .ZN(new_n809));
  OAI221_X1 g623(.A(new_n567), .B1(new_n808), .B2(new_n776), .C1(new_n809), .C2(KEYINPUT48), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n793), .A2(KEYINPUT114), .A3(new_n724), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT48), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n810), .B1(new_n813), .B2(new_n809), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n792), .A2(KEYINPUT51), .A3(new_n804), .A4(new_n794), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n807), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n675), .A2(new_n700), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n664), .A2(new_n631), .A3(new_n636), .ZN(new_n818));
  INV_X1    g632(.A(new_n725), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n818), .A2(new_n661), .A3(new_n659), .A4(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT93), .B1(new_n633), .B2(new_n644), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n647), .A2(new_n643), .A3(new_n646), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n817), .B(new_n820), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n649), .A2(KEYINPUT52), .A3(new_n817), .A4(new_n820), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AND4_X1   g641(.A1(new_n683), .A2(new_n686), .A3(new_n690), .A4(new_n697), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n614), .A2(new_n615), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n714), .A2(new_n829), .A3(new_n512), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n612), .A2(new_n636), .ZN(new_n831));
  AND4_X1   g645(.A1(new_n283), .A2(new_n830), .A3(new_n626), .A4(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n674), .A2(new_n696), .A3(new_n660), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n833), .A2(new_n729), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n476), .A2(new_n612), .A3(new_n513), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n836), .A2(new_n571), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n622), .A2(new_n345), .A3(new_n837), .A4(new_n421), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n573), .A2(new_n838), .A3(new_n627), .ZN(new_n839));
  INV_X1    g653(.A(new_n571), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT104), .B1(new_n663), .B2(new_n592), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT104), .ZN(new_n842));
  AOI211_X1 g656(.A(new_n842), .B(new_n591), .C1(new_n476), .C2(new_n513), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n840), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT105), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT105), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n846), .B(new_n840), .C1(new_n841), .C2(new_n843), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n845), .A2(new_n579), .A3(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n828), .A2(new_n835), .A3(new_n839), .A4(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n721), .A2(new_n732), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT106), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n848), .A2(new_n835), .A3(new_n839), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n718), .A2(new_n720), .B1(new_n730), .B2(new_n731), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT106), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n852), .A2(new_n853), .A3(new_n854), .A4(new_n828), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n827), .A2(new_n851), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n827), .A2(new_n851), .A3(new_n855), .A4(KEYINPUT53), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT54), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n849), .A2(new_n850), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n827), .A2(KEYINPUT53), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n858), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n861), .A2(KEYINPUT107), .A3(new_n865), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n865), .A2(KEYINPUT107), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n816), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n602), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n787), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n771), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT49), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n779), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n654), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n779), .A2(new_n872), .ZN(new_n875));
  NOR4_X1   g689(.A1(new_n874), .A2(new_n663), .A3(new_n875), .A4(new_n591), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n345), .A2(new_n348), .A3(new_n560), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n877), .B(KEYINPUT102), .Z(new_n878));
  NAND3_X1  g692(.A1(new_n876), .A2(new_n784), .A3(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT115), .B1(new_n871), .B2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT115), .ZN(new_n882));
  INV_X1    g696(.A(new_n870), .ZN(new_n883));
  AOI211_X1 g697(.A(new_n883), .B(new_n816), .C1(new_n866), .C2(new_n867), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n882), .B(new_n879), .C1(new_n884), .C2(new_n771), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n881), .A2(new_n885), .ZN(G75));
  NAND2_X1  g700(.A1(new_n530), .A2(new_n543), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT116), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  AOI211_X1 g703(.A(new_n187), .B(new_n276), .C1(new_n858), .C2(new_n864), .ZN(new_n890));
  OAI21_X1  g704(.A(KEYINPUT55), .B1(new_n890), .B2(KEYINPUT56), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n858), .A2(new_n864), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n892), .A2(G210), .A3(G902), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT55), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT56), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n542), .B(KEYINPUT117), .Z(new_n897));
  AND3_X1   g711(.A1(new_n891), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n897), .B1(new_n891), .B2(new_n896), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n889), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n330), .A2(G952), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n897), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n890), .A2(KEYINPUT55), .A3(KEYINPUT56), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n894), .B1(new_n893), .B2(new_n895), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n891), .A2(new_n896), .A3(new_n897), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n906), .A2(new_n888), .A3(new_n907), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n900), .A2(new_n902), .A3(new_n908), .ZN(G51));
  NAND2_X1  g723(.A1(new_n415), .A2(new_n418), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n892), .A2(KEYINPUT54), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT118), .ZN(new_n912));
  INV_X1    g726(.A(new_n865), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n704), .B(KEYINPUT57), .Z(new_n915));
  OAI21_X1  g729(.A(new_n910), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n892), .A2(G902), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n917), .A2(new_n737), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n901), .B1(new_n916), .B2(new_n918), .ZN(G54));
  NAND4_X1  g733(.A1(new_n892), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(new_n613), .Z(new_n921));
  NOR2_X1   g735(.A1(new_n921), .A2(new_n901), .ZN(G60));
  NAND2_X1  g736(.A1(new_n587), .A2(new_n589), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT119), .Z(new_n924));
  XNOR2_X1  g738(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n925));
  NAND2_X1  g739(.A1(G478), .A2(G902), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n914), .A2(new_n928), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n866), .A2(new_n867), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n924), .B1(new_n930), .B2(new_n927), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n929), .A2(new_n931), .A3(new_n901), .ZN(G63));
  NAND2_X1  g746(.A1(G217), .A2(G902), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT60), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n934), .B1(new_n858), .B2(new_n864), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n901), .B1(new_n935), .B2(new_n624), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n936), .B1(new_n338), .B2(new_n935), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(KEYINPUT121), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT61), .ZN(G66));
  OAI21_X1  g753(.A(G953), .B1(new_n563), .B2(new_n537), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n828), .A2(new_n839), .A3(new_n848), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n940), .B1(new_n942), .B2(G953), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n888), .B1(G898), .B2(new_n330), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(G69));
  NAND3_X1  g759(.A1(new_n455), .A2(new_n458), .A3(new_n457), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT122), .Z(new_n947));
  XOR2_X1   g761(.A(new_n255), .B(new_n947), .Z(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n769), .B1(new_n759), .B2(new_n761), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n649), .A2(new_n817), .ZN(new_n951));
  OR4_X1    g765(.A1(new_n724), .A2(new_n746), .A3(new_n631), .A4(new_n664), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n950), .A2(new_n951), .A3(new_n853), .A4(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n949), .B1(new_n953), .B2(new_n330), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n954), .B1(G227), .B2(new_n330), .ZN(new_n955));
  OAI21_X1  g769(.A(G900), .B1(new_n948), .B2(G227), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(G953), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n841), .A2(new_n843), .ZN(new_n958));
  AOI211_X1 g772(.A(new_n670), .B(new_n724), .C1(new_n836), .C2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n727), .ZN(new_n960));
  AOI21_X1  g774(.A(KEYINPUT62), .B1(new_n672), .B2(new_n951), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n672), .A2(new_n951), .A3(KEYINPUT62), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n950), .B(new_n960), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n963), .A2(new_n330), .A3(new_n949), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n955), .A2(new_n957), .A3(new_n964), .ZN(G72));
  INV_X1    g779(.A(KEYINPUT126), .ZN(new_n966));
  NAND2_X1  g780(.A1(G472), .A2(G902), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT63), .Z(new_n968));
  OAI21_X1  g782(.A(new_n968), .B1(new_n963), .B2(new_n941), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n655), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(KEYINPUT123), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT123), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n969), .A2(new_n972), .A3(new_n655), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n968), .B1(new_n953), .B2(new_n941), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n256), .A2(new_n191), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT124), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n655), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n860), .A2(new_n979), .A3(new_n968), .A4(new_n976), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n980), .A2(KEYINPUT125), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(KEYINPUT125), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n974), .B(new_n978), .C1(new_n981), .C2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n966), .B1(new_n984), .B2(new_n901), .ZN(new_n985));
  INV_X1    g799(.A(new_n981), .ZN(new_n986));
  AOI22_X1  g800(.A1(new_n986), .A2(new_n982), .B1(new_n975), .B2(new_n977), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n987), .A2(KEYINPUT126), .A3(new_n902), .A4(new_n974), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n985), .A2(new_n988), .ZN(G57));
endmodule


