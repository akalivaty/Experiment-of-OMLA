

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U552 ( .A1(n779), .A2(n778), .ZN(n794) );
  AND2_X1 U553 ( .A1(n519), .A2(n537), .ZN(n750) );
  OR2_X1 U554 ( .A1(n744), .A2(n743), .ZN(n741) );
  AND2_X1 U555 ( .A1(n518), .A2(n525), .ZN(G160) );
  NOR2_X1 U556 ( .A1(n732), .A2(n731), .ZN(n734) );
  OR2_X1 U557 ( .A1(n730), .A2(n1017), .ZN(n731) );
  XNOR2_X1 U558 ( .A(n755), .B(KEYINPUT100), .ZN(n763) );
  XNOR2_X1 U559 ( .A(n551), .B(KEYINPUT68), .ZN(n552) );
  NAND2_X1 U560 ( .A1(n549), .A2(n548), .ZN(n526) );
  XNOR2_X1 U561 ( .A(n545), .B(KEYINPUT23), .ZN(n546) );
  OR2_X1 U562 ( .A1(n735), .A2(n736), .ZN(n738) );
  INV_X1 U563 ( .A(KEYINPUT64), .ZN(n733) );
  XNOR2_X1 U564 ( .A(n538), .B(n749), .ZN(n537) );
  INV_X1 U565 ( .A(n842), .ZN(n536) );
  OR2_X1 U566 ( .A1(n768), .A2(n767), .ZN(n769) );
  INV_X1 U567 ( .A(KEYINPUT65), .ZN(n542) );
  NAND2_X1 U568 ( .A1(n550), .A2(G2104), .ZN(n540) );
  INV_X1 U569 ( .A(KEYINPUT40), .ZN(n535) );
  NAND2_X1 U570 ( .A1(n534), .A2(n532), .ZN(n531) );
  NAND2_X1 U571 ( .A1(n842), .A2(n533), .ZN(n532) );
  NAND2_X1 U572 ( .A1(n536), .A2(n535), .ZN(n534) );
  NAND2_X1 U573 ( .A1(n828), .A2(n535), .ZN(n533) );
  NAND2_X2 U574 ( .A1(n544), .A2(n543), .ZN(n886) );
  NAND2_X1 U575 ( .A1(n541), .A2(n550), .ZN(n543) );
  NAND2_X1 U576 ( .A1(n540), .A2(KEYINPUT65), .ZN(n544) );
  AND2_X1 U577 ( .A1(n542), .A2(G2104), .ZN(n541) );
  NOR2_X2 U578 ( .A1(G2104), .A2(n550), .ZN(n891) );
  NOR2_X1 U579 ( .A1(n661), .A2(n557), .ZN(n669) );
  XOR2_X1 U580 ( .A(KEYINPUT1), .B(n556), .Z(n666) );
  NOR2_X1 U581 ( .A1(G651), .A2(n661), .ZN(n673) );
  XNOR2_X1 U582 ( .A(n526), .B(KEYINPUT67), .ZN(n525) );
  AND2_X1 U583 ( .A1(n793), .A2(n524), .ZN(n517) );
  AND2_X1 U584 ( .A1(n555), .A2(n554), .ZN(n518) );
  XNOR2_X1 U585 ( .A(KEYINPUT28), .B(n728), .ZN(n519) );
  AND2_X1 U586 ( .A1(n793), .A2(n531), .ZN(n520) );
  OR2_X1 U587 ( .A1(G299), .A2(n748), .ZN(n521) );
  NAND2_X1 U588 ( .A1(n829), .A2(KEYINPUT40), .ZN(n522) );
  NOR2_X1 U589 ( .A1(n788), .A2(n785), .ZN(n523) );
  AND2_X1 U590 ( .A1(n842), .A2(n535), .ZN(n524) );
  NAND2_X1 U591 ( .A1(G160), .A2(G40), .ZN(n707) );
  NAND2_X1 U592 ( .A1(n794), .A2(n517), .ZN(n529) );
  NAND2_X1 U593 ( .A1(n528), .A2(n527), .ZN(n530) );
  NAND2_X1 U594 ( .A1(n531), .A2(n522), .ZN(n527) );
  NAND2_X1 U595 ( .A1(n794), .A2(n520), .ZN(n528) );
  NAND2_X1 U596 ( .A1(n530), .A2(n529), .ZN(G329) );
  NAND2_X1 U597 ( .A1(n521), .A2(n539), .ZN(n538) );
  XNOR2_X1 U598 ( .A(n747), .B(KEYINPUT98), .ZN(n539) );
  INV_X1 U599 ( .A(KEYINPUT97), .ZN(n739) );
  INV_X1 U600 ( .A(KEYINPUT99), .ZN(n749) );
  AND2_X1 U601 ( .A1(n836), .A2(n830), .ZN(n827) );
  INV_X1 U602 ( .A(KEYINPUT17), .ZN(n551) );
  NAND2_X1 U603 ( .A1(n827), .A2(n826), .ZN(n828) );
  INV_X1 U604 ( .A(G2105), .ZN(n550) );
  INV_X1 U605 ( .A(n828), .ZN(n829) );
  XNOR2_X1 U606 ( .A(n553), .B(n552), .ZN(n577) );
  NOR2_X1 U607 ( .A1(n601), .A2(n600), .ZN(n603) );
  NAND2_X1 U608 ( .A1(n603), .A2(n602), .ZN(n1017) );
  NAND2_X1 U609 ( .A1(G101), .A2(n886), .ZN(n547) );
  INV_X1 U610 ( .A(KEYINPUT66), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n547), .B(n546), .ZN(n549) );
  NAND2_X1 U612 ( .A1(G125), .A2(n891), .ZN(n548) );
  NOR2_X1 U613 ( .A1(G2105), .A2(G2104), .ZN(n553) );
  NAND2_X1 U614 ( .A1(G137), .A2(n577), .ZN(n555) );
  AND2_X1 U615 ( .A1(G2105), .A2(G2104), .ZN(n889) );
  NAND2_X1 U616 ( .A1(n889), .A2(G113), .ZN(n554) );
  INV_X1 U617 ( .A(G651), .ZN(n557) );
  NOR2_X1 U618 ( .A1(G543), .A2(n557), .ZN(n556) );
  NAND2_X1 U619 ( .A1(G65), .A2(n666), .ZN(n559) );
  XOR2_X1 U620 ( .A(KEYINPUT0), .B(G543), .Z(n661) );
  NAND2_X1 U621 ( .A1(G78), .A2(n669), .ZN(n558) );
  NAND2_X1 U622 ( .A1(n559), .A2(n558), .ZN(n563) );
  NOR2_X1 U623 ( .A1(G651), .A2(G543), .ZN(n665) );
  NAND2_X1 U624 ( .A1(G91), .A2(n665), .ZN(n561) );
  NAND2_X1 U625 ( .A1(G53), .A2(n673), .ZN(n560) );
  NAND2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n562) );
  OR2_X1 U627 ( .A1(n563), .A2(n562), .ZN(G299) );
  AND2_X1 U628 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U629 ( .A1(G123), .A2(n891), .ZN(n564) );
  XOR2_X1 U630 ( .A(KEYINPUT18), .B(n564), .Z(n570) );
  NAND2_X1 U631 ( .A1(n886), .A2(G99), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(KEYINPUT78), .ZN(n567) );
  NAND2_X1 U633 ( .A1(G111), .A2(n889), .ZN(n566) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U635 ( .A(KEYINPUT79), .B(n568), .Z(n569) );
  NOR2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n572) );
  NAND2_X1 U637 ( .A1(G135), .A2(n577), .ZN(n571) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n957) );
  XNOR2_X1 U639 ( .A(G2096), .B(n957), .ZN(n573) );
  OR2_X1 U640 ( .A1(G2100), .A2(n573), .ZN(G156) );
  INV_X1 U641 ( .A(G120), .ZN(G236) );
  INV_X1 U642 ( .A(G108), .ZN(G238) );
  INV_X1 U643 ( .A(G132), .ZN(G219) );
  INV_X1 U644 ( .A(G82), .ZN(G220) );
  NAND2_X1 U645 ( .A1(G114), .A2(n889), .ZN(n574) );
  XNOR2_X1 U646 ( .A(n574), .B(KEYINPUT88), .ZN(n576) );
  NAND2_X1 U647 ( .A1(n886), .A2(G102), .ZN(n575) );
  NAND2_X1 U648 ( .A1(n576), .A2(n575), .ZN(n581) );
  NAND2_X1 U649 ( .A1(G126), .A2(n891), .ZN(n579) );
  NAND2_X1 U650 ( .A1(G138), .A2(n577), .ZN(n578) );
  NAND2_X1 U651 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U652 ( .A1(n581), .A2(n580), .ZN(G164) );
  NAND2_X1 U653 ( .A1(n665), .A2(G89), .ZN(n582) );
  XNOR2_X1 U654 ( .A(n582), .B(KEYINPUT4), .ZN(n584) );
  NAND2_X1 U655 ( .A1(G76), .A2(n669), .ZN(n583) );
  NAND2_X1 U656 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U657 ( .A(n585), .B(KEYINPUT5), .ZN(n590) );
  NAND2_X1 U658 ( .A1(G63), .A2(n666), .ZN(n587) );
  NAND2_X1 U659 ( .A1(G51), .A2(n673), .ZN(n586) );
  NAND2_X1 U660 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U661 ( .A(KEYINPUT6), .B(n588), .Z(n589) );
  NAND2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U663 ( .A(n591), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U664 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U665 ( .A1(G7), .A2(G661), .ZN(n592) );
  XNOR2_X1 U666 ( .A(n592), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U667 ( .A(G567), .ZN(n702) );
  NOR2_X1 U668 ( .A1(n702), .A2(G223), .ZN(n593) );
  XNOR2_X1 U669 ( .A(n593), .B(KEYINPUT11), .ZN(G234) );
  NAND2_X1 U670 ( .A1(G56), .A2(n666), .ZN(n594) );
  XOR2_X1 U671 ( .A(KEYINPUT14), .B(n594), .Z(n601) );
  NAND2_X1 U672 ( .A1(n669), .A2(G68), .ZN(n595) );
  XNOR2_X1 U673 ( .A(KEYINPUT73), .B(n595), .ZN(n598) );
  NAND2_X1 U674 ( .A1(n665), .A2(G81), .ZN(n596) );
  XOR2_X1 U675 ( .A(KEYINPUT12), .B(n596), .Z(n597) );
  NOR2_X1 U676 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U677 ( .A(n599), .B(KEYINPUT13), .ZN(n600) );
  NAND2_X1 U678 ( .A1(n673), .A2(G43), .ZN(n602) );
  INV_X1 U679 ( .A(G860), .ZN(n627) );
  OR2_X1 U680 ( .A1(n1017), .A2(n627), .ZN(G153) );
  NAND2_X1 U681 ( .A1(G64), .A2(n666), .ZN(n604) );
  XOR2_X1 U682 ( .A(KEYINPUT70), .B(n604), .Z(n610) );
  NAND2_X1 U683 ( .A1(n669), .A2(G77), .ZN(n605) );
  XOR2_X1 U684 ( .A(KEYINPUT71), .B(n605), .Z(n607) );
  NAND2_X1 U685 ( .A1(n665), .A2(G90), .ZN(n606) );
  NAND2_X1 U686 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U687 ( .A(KEYINPUT9), .B(n608), .Z(n609) );
  NOR2_X1 U688 ( .A1(n610), .A2(n609), .ZN(n612) );
  NAND2_X1 U689 ( .A1(n673), .A2(G52), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n612), .A2(n611), .ZN(G301) );
  NAND2_X1 U691 ( .A1(G301), .A2(G868), .ZN(n613) );
  XNOR2_X1 U692 ( .A(n613), .B(KEYINPUT74), .ZN(n622) );
  INV_X1 U693 ( .A(G868), .ZN(n686) );
  NAND2_X1 U694 ( .A1(G66), .A2(n666), .ZN(n615) );
  NAND2_X1 U695 ( .A1(G79), .A2(n669), .ZN(n614) );
  NAND2_X1 U696 ( .A1(n615), .A2(n614), .ZN(n619) );
  NAND2_X1 U697 ( .A1(G92), .A2(n665), .ZN(n617) );
  NAND2_X1 U698 ( .A1(G54), .A2(n673), .ZN(n616) );
  NAND2_X1 U699 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U700 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U701 ( .A(KEYINPUT15), .B(n620), .Z(n1012) );
  INV_X1 U702 ( .A(n1012), .ZN(n744) );
  NAND2_X1 U703 ( .A1(n686), .A2(n744), .ZN(n621) );
  NAND2_X1 U704 ( .A1(n622), .A2(n621), .ZN(n623) );
  XOR2_X1 U705 ( .A(KEYINPUT75), .B(n623), .Z(G284) );
  NOR2_X1 U706 ( .A1(G868), .A2(G299), .ZN(n624) );
  XNOR2_X1 U707 ( .A(n624), .B(KEYINPUT76), .ZN(n626) );
  NOR2_X1 U708 ( .A1(n686), .A2(G286), .ZN(n625) );
  NOR2_X1 U709 ( .A1(n626), .A2(n625), .ZN(G297) );
  NAND2_X1 U710 ( .A1(n627), .A2(G559), .ZN(n628) );
  NAND2_X1 U711 ( .A1(n628), .A2(n1012), .ZN(n629) );
  XNOR2_X1 U712 ( .A(n629), .B(KEYINPUT16), .ZN(n630) );
  XOR2_X1 U713 ( .A(KEYINPUT77), .B(n630), .Z(G148) );
  NOR2_X1 U714 ( .A1(G868), .A2(n1017), .ZN(n633) );
  NAND2_X1 U715 ( .A1(G868), .A2(n1012), .ZN(n631) );
  NOR2_X1 U716 ( .A1(G559), .A2(n631), .ZN(n632) );
  NOR2_X1 U717 ( .A1(n633), .A2(n632), .ZN(G282) );
  NAND2_X1 U718 ( .A1(n1012), .A2(G559), .ZN(n684) );
  XNOR2_X1 U719 ( .A(n1017), .B(n684), .ZN(n634) );
  NOR2_X1 U720 ( .A1(n634), .A2(G860), .ZN(n642) );
  NAND2_X1 U721 ( .A1(G93), .A2(n665), .ZN(n636) );
  NAND2_X1 U722 ( .A1(G80), .A2(n669), .ZN(n635) );
  NAND2_X1 U723 ( .A1(n636), .A2(n635), .ZN(n641) );
  NAND2_X1 U724 ( .A1(G55), .A2(n673), .ZN(n637) );
  XNOR2_X1 U725 ( .A(n637), .B(KEYINPUT80), .ZN(n639) );
  NAND2_X1 U726 ( .A1(n666), .A2(G67), .ZN(n638) );
  NAND2_X1 U727 ( .A1(n639), .A2(n638), .ZN(n640) );
  OR2_X1 U728 ( .A1(n641), .A2(n640), .ZN(n687) );
  XOR2_X1 U729 ( .A(n642), .B(n687), .Z(G145) );
  NAND2_X1 U730 ( .A1(G88), .A2(n665), .ZN(n644) );
  NAND2_X1 U731 ( .A1(G75), .A2(n669), .ZN(n643) );
  NAND2_X1 U732 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U733 ( .A(KEYINPUT82), .B(n645), .ZN(n649) );
  NAND2_X1 U734 ( .A1(G62), .A2(n666), .ZN(n647) );
  NAND2_X1 U735 ( .A1(G50), .A2(n673), .ZN(n646) );
  NAND2_X1 U736 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U737 ( .A1(n649), .A2(n648), .ZN(n650) );
  XOR2_X1 U738 ( .A(KEYINPUT83), .B(n650), .Z(G166) );
  NAND2_X1 U739 ( .A1(G60), .A2(n666), .ZN(n652) );
  NAND2_X1 U740 ( .A1(G47), .A2(n673), .ZN(n651) );
  NAND2_X1 U741 ( .A1(n652), .A2(n651), .ZN(n655) );
  NAND2_X1 U742 ( .A1(G85), .A2(n665), .ZN(n653) );
  XNOR2_X1 U743 ( .A(KEYINPUT69), .B(n653), .ZN(n654) );
  NOR2_X1 U744 ( .A1(n655), .A2(n654), .ZN(n657) );
  NAND2_X1 U745 ( .A1(n669), .A2(G72), .ZN(n656) );
  NAND2_X1 U746 ( .A1(n657), .A2(n656), .ZN(G290) );
  NAND2_X1 U747 ( .A1(G49), .A2(n673), .ZN(n659) );
  NAND2_X1 U748 ( .A1(G74), .A2(G651), .ZN(n658) );
  NAND2_X1 U749 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U750 ( .A1(n666), .A2(n660), .ZN(n664) );
  NAND2_X1 U751 ( .A1(G87), .A2(n661), .ZN(n662) );
  XOR2_X1 U752 ( .A(KEYINPUT81), .B(n662), .Z(n663) );
  NAND2_X1 U753 ( .A1(n664), .A2(n663), .ZN(G288) );
  NAND2_X1 U754 ( .A1(G86), .A2(n665), .ZN(n668) );
  NAND2_X1 U755 ( .A1(G61), .A2(n666), .ZN(n667) );
  NAND2_X1 U756 ( .A1(n668), .A2(n667), .ZN(n672) );
  NAND2_X1 U757 ( .A1(n669), .A2(G73), .ZN(n670) );
  XOR2_X1 U758 ( .A(KEYINPUT2), .B(n670), .Z(n671) );
  NOR2_X1 U759 ( .A1(n672), .A2(n671), .ZN(n675) );
  NAND2_X1 U760 ( .A1(n673), .A2(G48), .ZN(n674) );
  NAND2_X1 U761 ( .A1(n675), .A2(n674), .ZN(G305) );
  XNOR2_X1 U762 ( .A(G166), .B(n1017), .ZN(n683) );
  XOR2_X1 U763 ( .A(G290), .B(G288), .Z(n676) );
  XNOR2_X1 U764 ( .A(G299), .B(n676), .ZN(n677) );
  XOR2_X1 U765 ( .A(n677), .B(KEYINPUT85), .Z(n679) );
  XNOR2_X1 U766 ( .A(KEYINPUT84), .B(KEYINPUT19), .ZN(n678) );
  XNOR2_X1 U767 ( .A(n679), .B(n678), .ZN(n680) );
  XOR2_X1 U768 ( .A(n687), .B(n680), .Z(n681) );
  XNOR2_X1 U769 ( .A(n681), .B(G305), .ZN(n682) );
  XNOR2_X1 U770 ( .A(n683), .B(n682), .ZN(n912) );
  XNOR2_X1 U771 ( .A(n912), .B(n684), .ZN(n685) );
  NOR2_X1 U772 ( .A1(n686), .A2(n685), .ZN(n689) );
  NOR2_X1 U773 ( .A1(G868), .A2(n687), .ZN(n688) );
  NOR2_X1 U774 ( .A1(n689), .A2(n688), .ZN(G295) );
  NAND2_X1 U775 ( .A1(G2084), .A2(G2078), .ZN(n690) );
  XOR2_X1 U776 ( .A(KEYINPUT20), .B(n690), .Z(n691) );
  NAND2_X1 U777 ( .A1(G2090), .A2(n691), .ZN(n692) );
  XNOR2_X1 U778 ( .A(KEYINPUT21), .B(n692), .ZN(n693) );
  NAND2_X1 U779 ( .A1(n693), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U780 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U781 ( .A(KEYINPUT72), .B(G57), .Z(G237) );
  NOR2_X1 U782 ( .A1(G220), .A2(G219), .ZN(n694) );
  XNOR2_X1 U783 ( .A(KEYINPUT22), .B(n694), .ZN(n695) );
  NAND2_X1 U784 ( .A1(n695), .A2(G96), .ZN(n696) );
  NOR2_X1 U785 ( .A1(G218), .A2(n696), .ZN(n697) );
  XNOR2_X1 U786 ( .A(KEYINPUT86), .B(n697), .ZN(n849) );
  INV_X1 U787 ( .A(n849), .ZN(n698) );
  NAND2_X1 U788 ( .A1(n698), .A2(G2106), .ZN(n699) );
  XNOR2_X1 U789 ( .A(n699), .B(KEYINPUT87), .ZN(n704) );
  NOR2_X1 U790 ( .A1(G237), .A2(G236), .ZN(n700) );
  NAND2_X1 U791 ( .A1(G69), .A2(n700), .ZN(n701) );
  NOR2_X1 U792 ( .A1(G238), .A2(n701), .ZN(n850) );
  NOR2_X1 U793 ( .A1(n702), .A2(n850), .ZN(n703) );
  NOR2_X1 U794 ( .A1(n704), .A2(n703), .ZN(G319) );
  INV_X1 U795 ( .A(G319), .ZN(n706) );
  NAND2_X1 U796 ( .A1(G483), .A2(G661), .ZN(n705) );
  NOR2_X1 U797 ( .A1(n706), .A2(n705), .ZN(n846) );
  NAND2_X1 U798 ( .A1(n846), .A2(G36), .ZN(G176) );
  INV_X1 U799 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U800 ( .A(KEYINPUT89), .B(G166), .ZN(G303) );
  XNOR2_X1 U801 ( .A(n707), .B(KEYINPUT90), .ZN(n796) );
  INV_X1 U802 ( .A(n796), .ZN(n708) );
  NOR2_X1 U803 ( .A1(G164), .A2(G1384), .ZN(n795) );
  NAND2_X2 U804 ( .A1(n708), .A2(n795), .ZN(n736) );
  NAND2_X1 U805 ( .A1(G8), .A2(n736), .ZN(n788) );
  NOR2_X1 U806 ( .A1(G1966), .A2(n788), .ZN(n765) );
  NOR2_X1 U807 ( .A1(G2084), .A2(n736), .ZN(n764) );
  NOR2_X1 U808 ( .A1(n765), .A2(n764), .ZN(n709) );
  XOR2_X1 U809 ( .A(KEYINPUT101), .B(n709), .Z(n710) );
  NAND2_X1 U810 ( .A1(G8), .A2(n710), .ZN(n711) );
  XNOR2_X1 U811 ( .A(KEYINPUT30), .B(n711), .ZN(n712) );
  NOR2_X1 U812 ( .A1(G168), .A2(n712), .ZN(n716) );
  INV_X1 U813 ( .A(G1961), .ZN(n988) );
  NAND2_X1 U814 ( .A1(n736), .A2(n988), .ZN(n714) );
  INV_X1 U815 ( .A(n736), .ZN(n724) );
  XNOR2_X1 U816 ( .A(G2078), .B(KEYINPUT25), .ZN(n937) );
  NAND2_X1 U817 ( .A1(n724), .A2(n937), .ZN(n713) );
  NAND2_X1 U818 ( .A1(n714), .A2(n713), .ZN(n751) );
  NOR2_X1 U819 ( .A1(G171), .A2(n751), .ZN(n715) );
  NOR2_X1 U820 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U821 ( .A(KEYINPUT31), .B(n717), .Z(n762) );
  INV_X1 U822 ( .A(G8), .ZN(n723) );
  NOR2_X1 U823 ( .A1(G1971), .A2(n788), .ZN(n719) );
  NOR2_X1 U824 ( .A1(G2090), .A2(n736), .ZN(n718) );
  NOR2_X1 U825 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U826 ( .A(n720), .B(KEYINPUT102), .ZN(n721) );
  NAND2_X1 U827 ( .A1(n721), .A2(G303), .ZN(n722) );
  OR2_X1 U828 ( .A1(n723), .A2(n722), .ZN(n757) );
  AND2_X1 U829 ( .A1(n762), .A2(n757), .ZN(n756) );
  NAND2_X1 U830 ( .A1(n724), .A2(G2072), .ZN(n725) );
  XOR2_X1 U831 ( .A(KEYINPUT27), .B(n725), .Z(n727) );
  NAND2_X1 U832 ( .A1(G1956), .A2(n736), .ZN(n726) );
  NAND2_X1 U833 ( .A1(n727), .A2(n726), .ZN(n748) );
  NAND2_X1 U834 ( .A1(G299), .A2(n748), .ZN(n728) );
  INV_X1 U835 ( .A(G1996), .ZN(n938) );
  NOR2_X1 U836 ( .A1(n736), .A2(n938), .ZN(n729) );
  XNOR2_X1 U837 ( .A(n729), .B(KEYINPUT26), .ZN(n732) );
  AND2_X1 U838 ( .A1(n736), .A2(G1341), .ZN(n730) );
  XNOR2_X1 U839 ( .A(n734), .B(n733), .ZN(n742) );
  INV_X1 U840 ( .A(G2067), .ZN(n735) );
  NAND2_X1 U841 ( .A1(G1348), .A2(n736), .ZN(n737) );
  NAND2_X1 U842 ( .A1(n738), .A2(n737), .ZN(n740) );
  XNOR2_X1 U843 ( .A(n740), .B(n739), .ZN(n743) );
  NAND2_X1 U844 ( .A1(n742), .A2(n741), .ZN(n746) );
  NAND2_X1 U845 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U846 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U847 ( .A(n750), .B(KEYINPUT29), .ZN(n754) );
  AND2_X1 U848 ( .A1(n751), .A2(G171), .ZN(n752) );
  XOR2_X1 U849 ( .A(KEYINPUT96), .B(n752), .Z(n753) );
  NAND2_X1 U850 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U851 ( .A1(n756), .A2(n763), .ZN(n760) );
  INV_X1 U852 ( .A(n757), .ZN(n758) );
  OR2_X1 U853 ( .A1(n758), .A2(G286), .ZN(n759) );
  NAND2_X1 U854 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U855 ( .A(n761), .B(KEYINPUT32), .ZN(n770) );
  AND2_X1 U856 ( .A1(n763), .A2(n762), .ZN(n768) );
  AND2_X1 U857 ( .A1(G8), .A2(n764), .ZN(n766) );
  OR2_X1 U858 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U859 ( .A1(n770), .A2(n769), .ZN(n784) );
  NOR2_X1 U860 ( .A1(G2090), .A2(G303), .ZN(n771) );
  NAND2_X1 U861 ( .A1(G8), .A2(n771), .ZN(n772) );
  NAND2_X1 U862 ( .A1(n784), .A2(n772), .ZN(n773) );
  NAND2_X1 U863 ( .A1(n773), .A2(n788), .ZN(n774) );
  XNOR2_X1 U864 ( .A(n774), .B(KEYINPUT103), .ZN(n779) );
  NOR2_X1 U865 ( .A1(G1981), .A2(G305), .ZN(n775) );
  XNOR2_X1 U866 ( .A(n775), .B(KEYINPUT24), .ZN(n776) );
  XNOR2_X1 U867 ( .A(n776), .B(KEYINPUT95), .ZN(n777) );
  NOR2_X1 U868 ( .A1(n788), .A2(n777), .ZN(n778) );
  NOR2_X1 U869 ( .A1(G1971), .A2(G303), .ZN(n780) );
  NOR2_X1 U870 ( .A1(G1976), .A2(G288), .ZN(n1022) );
  NOR2_X1 U871 ( .A1(n780), .A2(n1022), .ZN(n782) );
  INV_X1 U872 ( .A(KEYINPUT33), .ZN(n781) );
  AND2_X1 U873 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U874 ( .A1(n784), .A2(n783), .ZN(n787) );
  NAND2_X1 U875 ( .A1(G1976), .A2(G288), .ZN(n1025) );
  INV_X1 U876 ( .A(n1025), .ZN(n785) );
  OR2_X1 U877 ( .A1(KEYINPUT33), .A2(n523), .ZN(n786) );
  NAND2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n791) );
  NAND2_X1 U879 ( .A1(n1022), .A2(KEYINPUT33), .ZN(n789) );
  NOR2_X1 U880 ( .A1(n789), .A2(n788), .ZN(n790) );
  NOR2_X1 U881 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U882 ( .A(G1981), .B(G305), .Z(n1031) );
  NAND2_X1 U883 ( .A1(n792), .A2(n1031), .ZN(n793) );
  NOR2_X1 U884 ( .A1(n796), .A2(n795), .ZN(n840) );
  XNOR2_X1 U885 ( .A(G2067), .B(KEYINPUT37), .ZN(n838) );
  NAND2_X1 U886 ( .A1(G104), .A2(n886), .ZN(n798) );
  NAND2_X1 U887 ( .A1(G140), .A2(n577), .ZN(n797) );
  NAND2_X1 U888 ( .A1(n798), .A2(n797), .ZN(n800) );
  XOR2_X1 U889 ( .A(KEYINPUT91), .B(KEYINPUT34), .Z(n799) );
  XNOR2_X1 U890 ( .A(n800), .B(n799), .ZN(n805) );
  NAND2_X1 U891 ( .A1(G128), .A2(n891), .ZN(n802) );
  NAND2_X1 U892 ( .A1(G116), .A2(n889), .ZN(n801) );
  NAND2_X1 U893 ( .A1(n802), .A2(n801), .ZN(n803) );
  XOR2_X1 U894 ( .A(KEYINPUT35), .B(n803), .Z(n804) );
  NOR2_X1 U895 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U896 ( .A(KEYINPUT36), .B(n806), .ZN(n897) );
  NOR2_X1 U897 ( .A1(n838), .A2(n897), .ZN(n956) );
  NAND2_X1 U898 ( .A1(n840), .A2(n956), .ZN(n836) );
  NAND2_X1 U899 ( .A1(G95), .A2(n886), .ZN(n808) );
  NAND2_X1 U900 ( .A1(G131), .A2(n577), .ZN(n807) );
  NAND2_X1 U901 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U902 ( .A(n809), .B(KEYINPUT93), .ZN(n811) );
  NAND2_X1 U903 ( .A1(G107), .A2(n889), .ZN(n810) );
  NAND2_X1 U904 ( .A1(n811), .A2(n810), .ZN(n814) );
  NAND2_X1 U905 ( .A1(n891), .A2(G119), .ZN(n812) );
  XOR2_X1 U906 ( .A(KEYINPUT92), .B(n812), .Z(n813) );
  OR2_X1 U907 ( .A1(n814), .A2(n813), .ZN(n904) );
  AND2_X1 U908 ( .A1(n904), .A2(G1991), .ZN(n824) );
  NAND2_X1 U909 ( .A1(G105), .A2(n886), .ZN(n815) );
  XNOR2_X1 U910 ( .A(n815), .B(KEYINPUT38), .ZN(n822) );
  NAND2_X1 U911 ( .A1(G117), .A2(n889), .ZN(n817) );
  NAND2_X1 U912 ( .A1(G141), .A2(n577), .ZN(n816) );
  NAND2_X1 U913 ( .A1(n817), .A2(n816), .ZN(n820) );
  NAND2_X1 U914 ( .A1(n891), .A2(G129), .ZN(n818) );
  XOR2_X1 U915 ( .A(KEYINPUT94), .B(n818), .Z(n819) );
  NOR2_X1 U916 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U917 ( .A1(n822), .A2(n821), .ZN(n898) );
  AND2_X1 U918 ( .A1(n898), .A2(G1996), .ZN(n823) );
  NOR2_X1 U919 ( .A1(n824), .A2(n823), .ZN(n969) );
  INV_X1 U920 ( .A(n969), .ZN(n825) );
  NAND2_X1 U921 ( .A1(n825), .A2(n840), .ZN(n830) );
  XNOR2_X1 U922 ( .A(G1986), .B(G290), .ZN(n1016) );
  NAND2_X1 U923 ( .A1(n1016), .A2(n840), .ZN(n826) );
  NOR2_X1 U924 ( .A1(G1996), .A2(n898), .ZN(n964) );
  INV_X1 U925 ( .A(n830), .ZN(n833) );
  NOR2_X1 U926 ( .A1(G1986), .A2(G290), .ZN(n831) );
  NOR2_X1 U927 ( .A1(G1991), .A2(n904), .ZN(n955) );
  NOR2_X1 U928 ( .A1(n831), .A2(n955), .ZN(n832) );
  NOR2_X1 U929 ( .A1(n833), .A2(n832), .ZN(n834) );
  NOR2_X1 U930 ( .A1(n964), .A2(n834), .ZN(n835) );
  XNOR2_X1 U931 ( .A(n835), .B(KEYINPUT39), .ZN(n837) );
  NAND2_X1 U932 ( .A1(n837), .A2(n836), .ZN(n839) );
  NAND2_X1 U933 ( .A1(n838), .A2(n897), .ZN(n971) );
  NAND2_X1 U934 ( .A1(n839), .A2(n971), .ZN(n841) );
  NAND2_X1 U935 ( .A1(n841), .A2(n840), .ZN(n842) );
  INV_X1 U936 ( .A(G223), .ZN(n843) );
  NAND2_X1 U937 ( .A1(G2106), .A2(n843), .ZN(G217) );
  AND2_X1 U938 ( .A1(G15), .A2(G2), .ZN(n844) );
  NAND2_X1 U939 ( .A1(G661), .A2(n844), .ZN(G259) );
  NAND2_X1 U940 ( .A1(G3), .A2(G1), .ZN(n845) );
  XNOR2_X1 U941 ( .A(KEYINPUT104), .B(n845), .ZN(n847) );
  NAND2_X1 U942 ( .A1(n847), .A2(n846), .ZN(n848) );
  XOR2_X1 U943 ( .A(KEYINPUT105), .B(n848), .Z(G188) );
  XOR2_X1 U944 ( .A(G69), .B(KEYINPUT106), .Z(G235) );
  INV_X1 U946 ( .A(G96), .ZN(G221) );
  NAND2_X1 U947 ( .A1(n850), .A2(n849), .ZN(G261) );
  INV_X1 U948 ( .A(G261), .ZN(G325) );
  XOR2_X1 U949 ( .A(KEYINPUT42), .B(G2090), .Z(n852) );
  XNOR2_X1 U950 ( .A(G2078), .B(G2072), .ZN(n851) );
  XNOR2_X1 U951 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U952 ( .A(n853), .B(G2100), .Z(n855) );
  XNOR2_X1 U953 ( .A(G2067), .B(G2084), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U955 ( .A(G2096), .B(KEYINPUT43), .Z(n857) );
  XNOR2_X1 U956 ( .A(KEYINPUT107), .B(G2678), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U958 ( .A(n859), .B(n858), .Z(G227) );
  XNOR2_X1 U959 ( .A(G1996), .B(KEYINPUT41), .ZN(n869) );
  XOR2_X1 U960 ( .A(G1956), .B(G1961), .Z(n861) );
  XNOR2_X1 U961 ( .A(G1991), .B(G1981), .ZN(n860) );
  XNOR2_X1 U962 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U963 ( .A(G1966), .B(G1971), .Z(n863) );
  XNOR2_X1 U964 ( .A(G1986), .B(G1976), .ZN(n862) );
  XNOR2_X1 U965 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U966 ( .A(n865), .B(n864), .Z(n867) );
  XNOR2_X1 U967 ( .A(KEYINPUT108), .B(G2474), .ZN(n866) );
  XNOR2_X1 U968 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U969 ( .A(n869), .B(n868), .ZN(G229) );
  NAND2_X1 U970 ( .A1(G100), .A2(n886), .ZN(n871) );
  NAND2_X1 U971 ( .A1(G112), .A2(n889), .ZN(n870) );
  NAND2_X1 U972 ( .A1(n871), .A2(n870), .ZN(n877) );
  NAND2_X1 U973 ( .A1(n891), .A2(G124), .ZN(n872) );
  XNOR2_X1 U974 ( .A(n872), .B(KEYINPUT44), .ZN(n874) );
  NAND2_X1 U975 ( .A1(G136), .A2(n577), .ZN(n873) );
  NAND2_X1 U976 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U977 ( .A(KEYINPUT109), .B(n875), .Z(n876) );
  NOR2_X1 U978 ( .A1(n877), .A2(n876), .ZN(G162) );
  NAND2_X1 U979 ( .A1(G130), .A2(n891), .ZN(n879) );
  NAND2_X1 U980 ( .A1(G118), .A2(n889), .ZN(n878) );
  NAND2_X1 U981 ( .A1(n879), .A2(n878), .ZN(n884) );
  NAND2_X1 U982 ( .A1(G106), .A2(n886), .ZN(n881) );
  NAND2_X1 U983 ( .A1(G142), .A2(n577), .ZN(n880) );
  NAND2_X1 U984 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U985 ( .A(KEYINPUT45), .B(n882), .Z(n883) );
  NOR2_X1 U986 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U987 ( .A(G162), .B(n885), .ZN(n908) );
  NAND2_X1 U988 ( .A1(G103), .A2(n886), .ZN(n888) );
  NAND2_X1 U989 ( .A1(G139), .A2(n577), .ZN(n887) );
  NAND2_X1 U990 ( .A1(n888), .A2(n887), .ZN(n896) );
  NAND2_X1 U991 ( .A1(n889), .A2(G115), .ZN(n890) );
  XNOR2_X1 U992 ( .A(n890), .B(KEYINPUT110), .ZN(n893) );
  NAND2_X1 U993 ( .A1(G127), .A2(n891), .ZN(n892) );
  NAND2_X1 U994 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U995 ( .A(KEYINPUT47), .B(n894), .Z(n895) );
  NOR2_X1 U996 ( .A1(n896), .A2(n895), .ZN(n973) );
  XNOR2_X1 U997 ( .A(n973), .B(n897), .ZN(n899) );
  XNOR2_X1 U998 ( .A(n899), .B(n898), .ZN(n903) );
  XOR2_X1 U999 ( .A(KEYINPUT46), .B(KEYINPUT111), .Z(n901) );
  XNOR2_X1 U1000 ( .A(KEYINPUT112), .B(KEYINPUT48), .ZN(n900) );
  XNOR2_X1 U1001 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U1002 ( .A(n903), .B(n902), .Z(n906) );
  XOR2_X1 U1003 ( .A(G164), .B(n904), .Z(n905) );
  XNOR2_X1 U1004 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(n908), .B(n907), .ZN(n910) );
  XOR2_X1 U1006 ( .A(n957), .B(G160), .Z(n909) );
  XNOR2_X1 U1007 ( .A(n910), .B(n909), .ZN(n911) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n911), .ZN(G395) );
  XOR2_X1 U1009 ( .A(n912), .B(G286), .Z(n914) );
  XNOR2_X1 U1010 ( .A(G171), .B(n1012), .ZN(n913) );
  XNOR2_X1 U1011 ( .A(n914), .B(n913), .ZN(n915) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n915), .ZN(G397) );
  XOR2_X1 U1013 ( .A(G2451), .B(G2430), .Z(n917) );
  XNOR2_X1 U1014 ( .A(G2438), .B(G2443), .ZN(n916) );
  XNOR2_X1 U1015 ( .A(n917), .B(n916), .ZN(n923) );
  XOR2_X1 U1016 ( .A(G2435), .B(G2454), .Z(n919) );
  XNOR2_X1 U1017 ( .A(G1341), .B(G1348), .ZN(n918) );
  XNOR2_X1 U1018 ( .A(n919), .B(n918), .ZN(n921) );
  XOR2_X1 U1019 ( .A(G2446), .B(G2427), .Z(n920) );
  XNOR2_X1 U1020 ( .A(n921), .B(n920), .ZN(n922) );
  XOR2_X1 U1021 ( .A(n923), .B(n922), .Z(n924) );
  NAND2_X1 U1022 ( .A1(G14), .A2(n924), .ZN(n932) );
  NAND2_X1 U1023 ( .A1(G319), .A2(n932), .ZN(n929) );
  XNOR2_X1 U1024 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n926) );
  NOR2_X1 U1025 ( .A1(G227), .A2(G229), .ZN(n925) );
  XNOR2_X1 U1026 ( .A(n926), .B(n925), .ZN(n927) );
  XOR2_X1 U1027 ( .A(KEYINPUT49), .B(n927), .Z(n928) );
  NOR2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n931) );
  NOR2_X1 U1029 ( .A1(G395), .A2(G397), .ZN(n930) );
  NAND2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(G225) );
  INV_X1 U1031 ( .A(G225), .ZN(G308) );
  INV_X1 U1032 ( .A(n932), .ZN(G401) );
  XNOR2_X1 U1033 ( .A(KEYINPUT119), .B(G2090), .ZN(n933) );
  XNOR2_X1 U1034 ( .A(n933), .B(G35), .ZN(n951) );
  XOR2_X1 U1035 ( .A(G25), .B(G1991), .Z(n934) );
  NAND2_X1 U1036 ( .A1(n934), .A2(G28), .ZN(n944) );
  XNOR2_X1 U1037 ( .A(G2067), .B(G26), .ZN(n936) );
  XNOR2_X1 U1038 ( .A(G33), .B(G2072), .ZN(n935) );
  NOR2_X1 U1039 ( .A1(n936), .A2(n935), .ZN(n942) );
  XOR2_X1 U1040 ( .A(n937), .B(G27), .Z(n940) );
  XOR2_X1 U1041 ( .A(n938), .B(G32), .Z(n939) );
  NOR2_X1 U1042 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1043 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1044 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1045 ( .A(n945), .B(KEYINPUT120), .ZN(n946) );
  XNOR2_X1 U1046 ( .A(n946), .B(KEYINPUT53), .ZN(n949) );
  XNOR2_X1 U1047 ( .A(G2084), .B(G34), .ZN(n947) );
  XNOR2_X1 U1048 ( .A(KEYINPUT54), .B(n947), .ZN(n948) );
  NOR2_X1 U1049 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1050 ( .A1(n951), .A2(n950), .ZN(n954) );
  NOR2_X1 U1051 ( .A1(G29), .A2(KEYINPUT55), .ZN(n952) );
  NAND2_X1 U1052 ( .A1(n954), .A2(n952), .ZN(n953) );
  NAND2_X1 U1053 ( .A1(G11), .A2(n953), .ZN(n987) );
  INV_X1 U1054 ( .A(KEYINPUT55), .ZN(n981) );
  OR2_X1 U1055 ( .A1(n981), .A2(n954), .ZN(n985) );
  NOR2_X1 U1056 ( .A1(n956), .A2(n955), .ZN(n958) );
  NAND2_X1 U1057 ( .A1(n958), .A2(n957), .ZN(n961) );
  XNOR2_X1 U1058 ( .A(G2084), .B(G160), .ZN(n959) );
  XNOR2_X1 U1059 ( .A(KEYINPUT115), .B(n959), .ZN(n960) );
  NOR2_X1 U1060 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1061 ( .A(KEYINPUT116), .B(n962), .Z(n967) );
  XOR2_X1 U1062 ( .A(G2090), .B(G162), .Z(n963) );
  NOR2_X1 U1063 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1064 ( .A(KEYINPUT51), .B(n965), .ZN(n966) );
  NOR2_X1 U1065 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1067 ( .A(n970), .B(KEYINPUT117), .ZN(n972) );
  NAND2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n979) );
  XOR2_X1 U1069 ( .A(G164), .B(G2078), .Z(n976) );
  XOR2_X1 U1070 ( .A(n973), .B(KEYINPUT118), .Z(n974) );
  XNOR2_X1 U1071 ( .A(G2072), .B(n974), .ZN(n975) );
  NOR2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1073 ( .A(KEYINPUT50), .B(n977), .Z(n978) );
  NOR2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(n980), .B(KEYINPUT52), .ZN(n982) );
  NAND2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(G29), .A2(n983), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n1043) );
  XNOR2_X1 U1080 ( .A(G5), .B(n988), .ZN(n1007) );
  XNOR2_X1 U1081 ( .A(KEYINPUT59), .B(G1348), .ZN(n989) );
  XNOR2_X1 U1082 ( .A(n989), .B(G4), .ZN(n996) );
  XNOR2_X1 U1083 ( .A(G1956), .B(G20), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(G1981), .B(G6), .ZN(n991) );
  XNOR2_X1 U1085 ( .A(G19), .B(G1341), .ZN(n990) );
  NOR2_X1 U1086 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1087 ( .A(KEYINPUT125), .B(n992), .ZN(n993) );
  NOR2_X1 U1088 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1090 ( .A(KEYINPUT60), .B(n997), .ZN(n1005) );
  XNOR2_X1 U1091 ( .A(G1986), .B(G24), .ZN(n999) );
  XNOR2_X1 U1092 ( .A(G23), .B(G1976), .ZN(n998) );
  NOR2_X1 U1093 ( .A1(n999), .A2(n998), .ZN(n1002) );
  XOR2_X1 U1094 ( .A(G1971), .B(G22), .Z(n1000) );
  XNOR2_X1 U1095 ( .A(KEYINPUT126), .B(n1000), .ZN(n1001) );
  NAND2_X1 U1096 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1097 ( .A(KEYINPUT58), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1098 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1099 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  XNOR2_X1 U1100 ( .A(G21), .B(G1966), .ZN(n1008) );
  NOR2_X1 U1101 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1102 ( .A(KEYINPUT61), .B(n1010), .Z(n1011) );
  NOR2_X1 U1103 ( .A1(G16), .A2(n1011), .ZN(n1040) );
  XOR2_X1 U1104 ( .A(G16), .B(KEYINPUT56), .Z(n1038) );
  XOR2_X1 U1105 ( .A(G299), .B(G1956), .Z(n1014) );
  XNOR2_X1 U1106 ( .A(n1012), .B(G1348), .ZN(n1013) );
  NAND2_X1 U1107 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1108 ( .A1(n1016), .A2(n1015), .ZN(n1021) );
  XNOR2_X1 U1109 ( .A(G301), .B(G1961), .ZN(n1019) );
  XNOR2_X1 U1110 ( .A(n1017), .B(G1341), .ZN(n1018) );
  NOR2_X1 U1111 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1112 ( .A1(n1021), .A2(n1020), .ZN(n1029) );
  XOR2_X1 U1113 ( .A(n1022), .B(KEYINPUT121), .Z(n1024) );
  XNOR2_X1 U1114 ( .A(G303), .B(G1971), .ZN(n1023) );
  NOR2_X1 U1115 ( .A1(n1024), .A2(n1023), .ZN(n1026) );
  NAND2_X1 U1116 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1117 ( .A(KEYINPUT122), .B(n1027), .ZN(n1028) );
  NOR2_X1 U1118 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1119 ( .A(KEYINPUT123), .B(n1030), .ZN(n1035) );
  XNOR2_X1 U1120 ( .A(G1966), .B(G168), .ZN(n1032) );
  NAND2_X1 U1121 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XOR2_X1 U1122 ( .A(KEYINPUT57), .B(n1033), .Z(n1034) );
  NOR2_X1 U1123 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XNOR2_X1 U1124 ( .A(n1036), .B(KEYINPUT124), .ZN(n1037) );
  NOR2_X1 U1125 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NOR2_X1 U1126 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XOR2_X1 U1127 ( .A(KEYINPUT127), .B(n1041), .Z(n1042) );
  NAND2_X1 U1128 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
  XOR2_X1 U1129 ( .A(KEYINPUT62), .B(n1044), .Z(G311) );
  INV_X1 U1130 ( .A(G311), .ZN(G150) );
endmodule

