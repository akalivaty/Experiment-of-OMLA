

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753;

  XNOR2_X1 U377 ( .A(n396), .B(KEYINPUT32), .ZN(n752) );
  AND2_X1 U378 ( .A1(n613), .A2(n569), .ZN(n570) );
  XNOR2_X1 U379 ( .A(n391), .B(n433), .ZN(n463) );
  XNOR2_X1 U380 ( .A(n466), .B(n467), .ZN(n721) );
  BUF_X1 U381 ( .A(G143), .Z(n354) );
  AND2_X2 U382 ( .A1(n627), .A2(n730), .ZN(n374) );
  NOR2_X2 U383 ( .A1(n659), .A2(n571), .ZN(n574) );
  XOR2_X2 U384 ( .A(n567), .B(KEYINPUT38), .Z(n672) );
  AND2_X2 U385 ( .A1(n546), .A2(n606), .ZN(n543) );
  XNOR2_X2 U386 ( .A(KEYINPUT86), .B(KEYINPUT74), .ZN(n388) );
  INV_X2 U387 ( .A(G953), .ZN(n745) );
  INV_X1 U388 ( .A(n623), .ZN(n686) );
  XNOR2_X2 U389 ( .A(n490), .B(n489), .ZN(n544) );
  XNOR2_X1 U390 ( .A(n484), .B(n483), .ZN(n522) );
  XOR2_X2 U391 ( .A(G113), .B(G104), .Z(n465) );
  XOR2_X2 U392 ( .A(G122), .B(G107), .Z(n464) );
  AND2_X1 U393 ( .A1(n418), .A2(n553), .ZN(n417) );
  XNOR2_X1 U394 ( .A(n376), .B(KEYINPUT35), .ZN(n750) );
  XNOR2_X1 U395 ( .A(n570), .B(KEYINPUT39), .ZN(n571) );
  XNOR2_X1 U396 ( .A(n372), .B(n535), .ZN(n704) );
  OR2_X1 U397 ( .A1(n606), .A2(n534), .ZN(n372) );
  NOR2_X1 U398 ( .A1(n529), .A2(n530), .ZN(n655) );
  XNOR2_X1 U399 ( .A(n390), .B(n389), .ZN(n590) );
  XNOR2_X1 U400 ( .A(n544), .B(n415), .ZN(n579) );
  XNOR2_X1 U401 ( .A(n426), .B(n425), .ZN(n631) );
  XNOR2_X1 U402 ( .A(n463), .B(n392), .ZN(n710) );
  XNOR2_X1 U403 ( .A(n513), .B(n427), .ZN(n735) );
  XNOR2_X1 U404 ( .A(KEYINPUT36), .B(KEYINPUT83), .ZN(n608) );
  INV_X2 U405 ( .A(G143), .ZN(n370) );
  BUF_X1 U406 ( .A(n642), .Z(n355) );
  XNOR2_X1 U407 ( .A(n446), .B(G125), .ZN(n468) );
  INV_X1 U408 ( .A(G146), .ZN(n446) );
  XNOR2_X1 U409 ( .A(n588), .B(n587), .ZN(n600) );
  XNOR2_X1 U410 ( .A(G137), .B(G134), .ZN(n500) );
  AND2_X1 U411 ( .A1(n579), .A2(n413), .ZN(n580) );
  AND2_X1 U412 ( .A1(n578), .A2(n414), .ZN(n413) );
  INV_X1 U413 ( .A(n602), .ZN(n414) );
  XNOR2_X1 U414 ( .A(n452), .B(n423), .ZN(n539) );
  XNOR2_X1 U415 ( .A(n424), .B(G475), .ZN(n423) );
  INV_X1 U416 ( .A(KEYINPUT13), .ZN(n424) );
  XNOR2_X1 U417 ( .A(n379), .B(G469), .ZN(n582) );
  OR2_X1 U418 ( .A1(n636), .A2(G902), .ZN(n379) );
  XNOR2_X1 U419 ( .A(n736), .B(n492), .ZN(n391) );
  NOR2_X1 U420 ( .A1(G953), .A2(G237), .ZN(n451) );
  XNOR2_X1 U421 ( .A(n468), .B(n447), .ZN(n513) );
  AND2_X1 U422 ( .A1(n612), .A2(n568), .ZN(n569) );
  XNOR2_X1 U423 ( .A(n395), .B(n394), .ZN(n552) );
  INV_X1 U424 ( .A(KEYINPUT82), .ZN(n394) );
  NAND2_X1 U425 ( .A1(n538), .A2(n539), .ZN(n575) );
  NOR2_X1 U426 ( .A1(G902), .A2(n488), .ZN(n490) );
  XNOR2_X1 U427 ( .A(n383), .B(n520), .ZN(n578) );
  XNOR2_X1 U428 ( .A(n519), .B(n518), .ZN(n520) );
  INV_X1 U429 ( .A(KEYINPUT25), .ZN(n518) );
  XNOR2_X1 U430 ( .A(G131), .B(KEYINPUT5), .ZN(n435) );
  XNOR2_X1 U431 ( .A(n500), .B(n434), .ZN(n412) );
  XNOR2_X1 U432 ( .A(G146), .B(G113), .ZN(n434) );
  AND2_X1 U433 ( .A1(n381), .A2(n398), .ZN(n402) );
  NAND2_X1 U434 ( .A1(n403), .A2(n401), .ZN(n400) );
  XNOR2_X1 U435 ( .A(n385), .B(n384), .ZN(n512) );
  INV_X1 U436 ( .A(KEYINPUT8), .ZN(n384) );
  NAND2_X1 U437 ( .A1(n745), .A2(G234), .ZN(n385) );
  XNOR2_X1 U438 ( .A(G128), .B(G119), .ZN(n506) );
  XNOR2_X1 U439 ( .A(G140), .B(KEYINPUT23), .ZN(n508) );
  XNOR2_X1 U440 ( .A(n450), .B(n358), .ZN(n425) );
  XNOR2_X1 U441 ( .A(n449), .B(n735), .ZN(n426) );
  XNOR2_X1 U442 ( .A(n503), .B(n502), .ZN(n636) );
  XNOR2_X1 U443 ( .A(n373), .B(n471), .ZN(n393) );
  NOR2_X1 U444 ( .A1(n562), .A2(n561), .ZN(n380) );
  NAND2_X1 U445 ( .A1(n375), .A2(n356), .ZN(n422) );
  INV_X1 U446 ( .A(KEYINPUT47), .ZN(n408) );
  OR2_X1 U447 ( .A1(G237), .A2(G902), .ZN(n475) );
  INV_X1 U448 ( .A(G101), .ZN(n492) );
  AND2_X1 U449 ( .A1(n600), .A2(n407), .ZN(n401) );
  NOR2_X1 U450 ( .A1(n621), .A2(n668), .ZN(n397) );
  NAND2_X1 U451 ( .A1(n406), .A2(n399), .ZN(n398) );
  NOR2_X1 U452 ( .A1(n668), .A2(n621), .ZN(n399) );
  XNOR2_X1 U453 ( .A(KEYINPUT4), .B(KEYINPUT66), .ZN(n430) );
  NOR2_X1 U454 ( .A1(n552), .A2(n549), .ZN(n550) );
  XNOR2_X1 U455 ( .A(G902), .B(KEYINPUT15), .ZN(n628) );
  INV_X1 U456 ( .A(n494), .ZN(n427) );
  XNOR2_X1 U457 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n444) );
  XOR2_X1 U458 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n445) );
  XOR2_X1 U459 ( .A(G107), .B(KEYINPUT73), .Z(n498) );
  XOR2_X1 U460 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n470) );
  XNOR2_X1 U461 ( .A(n387), .B(n468), .ZN(n373) );
  XNOR2_X1 U462 ( .A(n388), .B(KEYINPUT85), .ZN(n387) );
  XNOR2_X1 U463 ( .A(KEYINPUT3), .B(KEYINPUT68), .ZN(n431) );
  XOR2_X1 U464 ( .A(G116), .B(G119), .Z(n432) );
  XOR2_X1 U465 ( .A(G110), .B(KEYINPUT16), .Z(n467) );
  XNOR2_X1 U466 ( .A(G116), .B(G134), .ZN(n455) );
  INV_X1 U467 ( .A(n628), .ZN(n472) );
  NAND2_X1 U468 ( .A1(n730), .A2(n386), .ZN(n375) );
  BUF_X1 U469 ( .A(n522), .Z(n526) );
  NOR2_X1 U470 ( .A1(n584), .A2(n583), .ZN(n589) );
  INV_X1 U471 ( .A(KEYINPUT102), .ZN(n415) );
  INV_X1 U472 ( .A(KEYINPUT22), .ZN(n486) );
  XNOR2_X1 U473 ( .A(n582), .B(n378), .ZN(n623) );
  INV_X1 U474 ( .A(KEYINPUT1), .ZN(n378) );
  XNOR2_X1 U475 ( .A(n524), .B(KEYINPUT92), .ZN(n562) );
  XNOR2_X1 U476 ( .A(n437), .B(n412), .ZN(n439) );
  XNOR2_X1 U477 ( .A(n515), .B(n516), .ZN(n716) );
  XNOR2_X1 U478 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U479 ( .A(n636), .B(n428), .ZN(n637) );
  XNOR2_X1 U480 ( .A(n375), .B(n670), .ZN(n702) );
  XNOR2_X1 U481 ( .A(n572), .B(KEYINPUT108), .ZN(n573) );
  INV_X1 U482 ( .A(KEYINPUT56), .ZN(n364) );
  INV_X1 U483 ( .A(n668), .ZN(n407) );
  AND2_X1 U484 ( .A1(n472), .A2(KEYINPUT2), .ZN(n356) );
  NOR2_X1 U485 ( .A1(n578), .A2(n523), .ZN(n357) );
  AND2_X1 U486 ( .A1(G214), .A2(n451), .ZN(n358) );
  XOR2_X1 U487 ( .A(n488), .B(KEYINPUT62), .Z(n359) );
  XNOR2_X1 U488 ( .A(n620), .B(KEYINPUT48), .ZN(n621) );
  XOR2_X1 U489 ( .A(n710), .B(n711), .Z(n360) );
  AND2_X1 U490 ( .A1(n472), .A2(n670), .ZN(n361) );
  AND2_X1 U491 ( .A1(n596), .A2(n408), .ZN(n362) );
  NOR2_X1 U492 ( .A1(G952), .A2(n745), .ZN(n720) );
  INV_X1 U493 ( .A(n720), .ZN(n368) );
  XNOR2_X1 U494 ( .A(n393), .B(n721), .ZN(n392) );
  XNOR2_X1 U495 ( .A(n474), .B(n473), .ZN(n566) );
  NOR2_X1 U496 ( .A1(n472), .A2(n710), .ZN(n474) );
  NAND2_X1 U497 ( .A1(n429), .A2(G475), .ZN(n633) );
  XNOR2_X1 U498 ( .A(n363), .B(n635), .ZN(G60) );
  NAND2_X1 U499 ( .A1(n634), .A2(n368), .ZN(n363) );
  XNOR2_X1 U500 ( .A(n365), .B(n364), .ZN(G51) );
  NAND2_X1 U501 ( .A1(n366), .A2(n368), .ZN(n365) );
  XNOR2_X1 U502 ( .A(n712), .B(n360), .ZN(n366) );
  NAND2_X1 U503 ( .A1(n374), .A2(n361), .ZN(n371) );
  XNOR2_X1 U504 ( .A(n367), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U505 ( .A1(n369), .A2(n368), .ZN(n367) );
  XNOR2_X1 U506 ( .A(n629), .B(n359), .ZN(n369) );
  NAND2_X2 U507 ( .A1(n371), .A2(n422), .ZN(n429) );
  XNOR2_X1 U508 ( .A(n543), .B(KEYINPUT79), .ZN(n504) );
  XNOR2_X2 U509 ( .A(n459), .B(n430), .ZN(n736) );
  XNOR2_X2 U510 ( .A(n370), .B(G128), .ZN(n459) );
  NAND2_X1 U511 ( .A1(n382), .A2(n397), .ZN(n381) );
  NAND2_X2 U512 ( .A1(n626), .A2(n669), .ZN(n743) );
  XNOR2_X1 U513 ( .A(n421), .B(KEYINPUT81), .ZN(n420) );
  NAND2_X1 U514 ( .A1(n420), .A2(n417), .ZN(n416) );
  NAND2_X1 U515 ( .A1(n522), .A2(n485), .ZN(n487) );
  NAND2_X1 U516 ( .A1(n541), .A2(n540), .ZN(n421) );
  NAND2_X1 U517 ( .A1(n750), .A2(KEYINPUT44), .ZN(n540) );
  NAND2_X1 U518 ( .A1(n377), .A2(n616), .ZN(n376) );
  XNOR2_X1 U519 ( .A(n537), .B(KEYINPUT34), .ZN(n377) );
  XNOR2_X1 U520 ( .A(n380), .B(KEYINPUT72), .ZN(n613) );
  INV_X1 U521 ( .A(n600), .ZN(n382) );
  NOR2_X1 U522 ( .A1(n716), .A2(G902), .ZN(n383) );
  INV_X1 U523 ( .A(n743), .ZN(n386) );
  XNOR2_X2 U524 ( .A(n416), .B(KEYINPUT45), .ZN(n730) );
  INV_X1 U525 ( .A(n567), .ZN(n607) );
  NAND2_X1 U526 ( .A1(n590), .A2(n482), .ZN(n484) );
  INV_X1 U527 ( .A(KEYINPUT19), .ZN(n389) );
  NOR2_X2 U528 ( .A1(n566), .A2(n671), .ZN(n390) );
  NAND2_X1 U529 ( .A1(n752), .A2(n650), .ZN(n395) );
  NAND2_X1 U530 ( .A1(n543), .A2(n542), .ZN(n396) );
  NAND2_X1 U531 ( .A1(n619), .A2(n621), .ZN(n404) );
  INV_X1 U532 ( .A(n599), .ZN(n405) );
  NAND2_X1 U533 ( .A1(n402), .A2(n400), .ZN(n626) );
  NOR2_X1 U534 ( .A1(n405), .A2(n404), .ZN(n403) );
  NAND2_X1 U535 ( .A1(n599), .A2(n619), .ZN(n406) );
  NAND2_X1 U536 ( .A1(n409), .A2(n362), .ZN(n597) );
  NAND2_X1 U537 ( .A1(n411), .A2(n410), .ZN(n409) );
  INV_X1 U538 ( .A(KEYINPUT65), .ZN(n410) );
  NAND2_X1 U539 ( .A1(n592), .A2(n595), .ZN(n411) );
  XNOR2_X1 U540 ( .A(n550), .B(n419), .ZN(n418) );
  INV_X1 U541 ( .A(KEYINPUT64), .ZN(n419) );
  XNOR2_X1 U542 ( .A(n492), .B(G146), .ZN(n493) );
  XNOR2_X1 U543 ( .A(n487), .B(n486), .ZN(n546) );
  XNOR2_X1 U544 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n428) );
  INV_X1 U545 ( .A(KEYINPUT67), .ZN(n620) );
  XNOR2_X1 U546 ( .A(n448), .B(n354), .ZN(n449) );
  INV_X1 U547 ( .A(n722), .ZN(n433) );
  INV_X1 U548 ( .A(KEYINPUT10), .ZN(n447) );
  INV_X1 U549 ( .A(KEYINPUT0), .ZN(n483) );
  XNOR2_X1 U550 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U551 ( .A(n609), .B(n608), .ZN(n610) );
  XNOR2_X1 U552 ( .A(n432), .B(n431), .ZN(n722) );
  XOR2_X1 U553 ( .A(KEYINPUT93), .B(KEYINPUT70), .Z(n436) );
  XNOR2_X1 U554 ( .A(n436), .B(n435), .ZN(n437) );
  NAND2_X1 U555 ( .A1(n451), .A2(G210), .ZN(n438) );
  XNOR2_X1 U556 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U557 ( .A(n463), .B(n440), .ZN(n488) );
  XOR2_X1 U558 ( .A(KEYINPUT90), .B(KEYINPUT21), .Z(n443) );
  NAND2_X1 U559 ( .A1(G234), .A2(n628), .ZN(n441) );
  XNOR2_X1 U560 ( .A(KEYINPUT20), .B(n441), .ZN(n517) );
  NAND2_X1 U561 ( .A1(n517), .A2(G221), .ZN(n442) );
  XNOR2_X1 U562 ( .A(n443), .B(n442), .ZN(n683) );
  XNOR2_X1 U563 ( .A(n683), .B(KEYINPUT91), .ZN(n523) );
  XNOR2_X1 U564 ( .A(n445), .B(n444), .ZN(n450) );
  XOR2_X1 U565 ( .A(G131), .B(G140), .Z(n494) );
  XOR2_X1 U566 ( .A(G122), .B(n465), .Z(n448) );
  NOR2_X1 U567 ( .A1(G902), .A2(n631), .ZN(n452) );
  XOR2_X1 U568 ( .A(KEYINPUT7), .B(KEYINPUT98), .Z(n454) );
  NAND2_X1 U569 ( .A1(G217), .A2(n512), .ZN(n453) );
  XNOR2_X1 U570 ( .A(n454), .B(n453), .ZN(n458) );
  XOR2_X1 U571 ( .A(KEYINPUT9), .B(KEYINPUT99), .Z(n456) );
  XNOR2_X1 U572 ( .A(n456), .B(n455), .ZN(n457) );
  XOR2_X1 U573 ( .A(n458), .B(n457), .Z(n461) );
  XNOR2_X1 U574 ( .A(n459), .B(n464), .ZN(n460) );
  XNOR2_X1 U575 ( .A(n461), .B(n460), .ZN(n714) );
  NOR2_X1 U576 ( .A1(n714), .A2(G902), .ZN(n462) );
  XOR2_X1 U577 ( .A(n462), .B(G478), .Z(n530) );
  INV_X1 U578 ( .A(n530), .ZN(n538) );
  NOR2_X1 U579 ( .A1(n523), .A2(n575), .ZN(n485) );
  XNOR2_X1 U580 ( .A(n465), .B(n464), .ZN(n466) );
  NAND2_X1 U581 ( .A1(G224), .A2(n745), .ZN(n469) );
  XNOR2_X1 U582 ( .A(n470), .B(n469), .ZN(n471) );
  AND2_X1 U583 ( .A1(G210), .A2(n475), .ZN(n473) );
  NAND2_X1 U584 ( .A1(n475), .A2(G214), .ZN(n476) );
  XNOR2_X1 U585 ( .A(KEYINPUT87), .B(n476), .ZN(n671) );
  INV_X1 U586 ( .A(n671), .ZN(n563) );
  NAND2_X1 U587 ( .A1(G234), .A2(G237), .ZN(n477) );
  XNOR2_X1 U588 ( .A(n477), .B(KEYINPUT14), .ZN(n478) );
  AND2_X1 U589 ( .A1(G952), .A2(n478), .ZN(n699) );
  NAND2_X1 U590 ( .A1(n699), .A2(n745), .ZN(n557) );
  NOR2_X1 U591 ( .A1(G898), .A2(n745), .ZN(n726) );
  NAND2_X1 U592 ( .A1(G902), .A2(n478), .ZN(n554) );
  INV_X1 U593 ( .A(n554), .ZN(n479) );
  NAND2_X1 U594 ( .A1(n726), .A2(n479), .ZN(n480) );
  NAND2_X1 U595 ( .A1(n557), .A2(n480), .ZN(n481) );
  XNOR2_X1 U596 ( .A(KEYINPUT88), .B(n481), .ZN(n482) );
  XNOR2_X1 U597 ( .A(G472), .B(KEYINPUT94), .ZN(n489) );
  XNOR2_X1 U598 ( .A(n544), .B(KEYINPUT100), .ZN(n491) );
  XOR2_X1 U599 ( .A(n491), .B(KEYINPUT6), .Z(n606) );
  XNOR2_X1 U600 ( .A(n736), .B(n493), .ZN(n496) );
  XOR2_X1 U601 ( .A(G110), .B(n494), .Z(n495) );
  XNOR2_X1 U602 ( .A(n496), .B(n495), .ZN(n503) );
  NAND2_X1 U603 ( .A1(G227), .A2(n745), .ZN(n497) );
  XNOR2_X1 U604 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U605 ( .A(G104), .B(n499), .ZN(n501) );
  XNOR2_X1 U606 ( .A(KEYINPUT89), .B(n500), .ZN(n738) );
  XNOR2_X1 U607 ( .A(n501), .B(n738), .ZN(n502) );
  NOR2_X2 U608 ( .A1(n504), .A2(n686), .ZN(n505) );
  XNOR2_X1 U609 ( .A(n505), .B(KEYINPUT80), .ZN(n521) );
  XOR2_X1 U610 ( .A(G110), .B(G137), .Z(n507) );
  XNOR2_X1 U611 ( .A(n507), .B(n506), .ZN(n511) );
  XOR2_X1 U612 ( .A(KEYINPUT77), .B(KEYINPUT24), .Z(n509) );
  XNOR2_X1 U613 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U614 ( .A(n511), .B(n510), .Z(n516) );
  NAND2_X1 U615 ( .A1(G221), .A2(n512), .ZN(n514) );
  NAND2_X1 U616 ( .A1(n517), .A2(G217), .ZN(n519) );
  INV_X1 U617 ( .A(n578), .ZN(n682) );
  NAND2_X1 U618 ( .A1(n521), .A2(n682), .ZN(n642) );
  INV_X1 U619 ( .A(n526), .ZN(n536) );
  NAND2_X1 U620 ( .A1(n582), .A2(n357), .ZN(n524) );
  NOR2_X1 U621 ( .A1(n536), .A2(n562), .ZN(n525) );
  NAND2_X1 U622 ( .A1(n544), .A2(n525), .ZN(n644) );
  NAND2_X1 U623 ( .A1(n686), .A2(n357), .ZN(n534) );
  NOR2_X1 U624 ( .A1(n544), .A2(n534), .ZN(n691) );
  NAND2_X1 U625 ( .A1(n691), .A2(n526), .ZN(n527) );
  XOR2_X1 U626 ( .A(KEYINPUT31), .B(n527), .Z(n663) );
  NAND2_X1 U627 ( .A1(n644), .A2(n663), .ZN(n531) );
  INV_X1 U628 ( .A(KEYINPUT97), .ZN(n528) );
  XNOR2_X1 U629 ( .A(n528), .B(n539), .ZN(n529) );
  INV_X1 U630 ( .A(n655), .ZN(n659) );
  NAND2_X1 U631 ( .A1(n530), .A2(n529), .ZN(n664) );
  NAND2_X1 U632 ( .A1(n659), .A2(n664), .ZN(n675) );
  NAND2_X1 U633 ( .A1(n531), .A2(n675), .ZN(n532) );
  NAND2_X1 U634 ( .A1(n642), .A2(n532), .ZN(n533) );
  XNOR2_X1 U635 ( .A(n533), .B(KEYINPUT101), .ZN(n541) );
  XOR2_X1 U636 ( .A(KEYINPUT84), .B(KEYINPUT33), .Z(n535) );
  NOR2_X1 U637 ( .A1(n536), .A2(n704), .ZN(n537) );
  NOR2_X1 U638 ( .A1(n539), .A2(n538), .ZN(n616) );
  NOR2_X1 U639 ( .A1(n682), .A2(n623), .ZN(n542) );
  INV_X1 U640 ( .A(n579), .ZN(n545) );
  NAND2_X1 U641 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U642 ( .A1(n682), .A2(n547), .ZN(n548) );
  NAND2_X1 U643 ( .A1(n623), .A2(n548), .ZN(n650) );
  INV_X1 U644 ( .A(KEYINPUT44), .ZN(n549) );
  NOR2_X1 U645 ( .A1(n750), .A2(KEYINPUT44), .ZN(n551) );
  NAND2_X1 U646 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U647 ( .A1(G900), .A2(n554), .ZN(n555) );
  NAND2_X1 U648 ( .A1(G953), .A2(n555), .ZN(n556) );
  XNOR2_X1 U649 ( .A(KEYINPUT103), .B(n556), .ZN(n559) );
  INV_X1 U650 ( .A(n557), .ZN(n558) );
  NOR2_X1 U651 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U652 ( .A(n560), .B(KEYINPUT76), .Z(n577) );
  INV_X1 U653 ( .A(n577), .ZN(n561) );
  XOR2_X1 U654 ( .A(KEYINPUT104), .B(KEYINPUT30), .Z(n565) );
  NAND2_X1 U655 ( .A1(n579), .A2(n563), .ZN(n564) );
  XNOR2_X1 U656 ( .A(n565), .B(n564), .ZN(n612) );
  BUF_X1 U657 ( .A(n566), .Z(n567) );
  INV_X1 U658 ( .A(n672), .ZN(n568) );
  NOR2_X1 U659 ( .A1(n664), .A2(n571), .ZN(n668) );
  INV_X1 U660 ( .A(KEYINPUT40), .ZN(n572) );
  XNOR2_X1 U661 ( .A(n574), .B(n573), .ZN(n749) );
  XOR2_X1 U662 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n586) );
  NOR2_X1 U663 ( .A1(n671), .A2(n672), .ZN(n676) );
  INV_X1 U664 ( .A(n575), .ZN(n673) );
  NAND2_X1 U665 ( .A1(n676), .A2(n673), .ZN(n576) );
  XOR2_X1 U666 ( .A(n576), .B(KEYINPUT41), .Z(n703) );
  INV_X1 U667 ( .A(n703), .ZN(n693) );
  XNOR2_X1 U668 ( .A(KEYINPUT107), .B(KEYINPUT28), .ZN(n581) );
  NAND2_X1 U669 ( .A1(n683), .A2(n577), .ZN(n602) );
  XNOR2_X1 U670 ( .A(n581), .B(n580), .ZN(n584) );
  XOR2_X1 U671 ( .A(KEYINPUT106), .B(n582), .Z(n583) );
  NAND2_X1 U672 ( .A1(n693), .A2(n589), .ZN(n585) );
  XNOR2_X1 U673 ( .A(n586), .B(n585), .ZN(n753) );
  NAND2_X1 U674 ( .A1(n749), .A2(n753), .ZN(n588) );
  XOR2_X1 U675 ( .A(KEYINPUT78), .B(KEYINPUT46), .Z(n587) );
  INV_X1 U676 ( .A(KEYINPUT69), .ZN(n595) );
  XOR2_X1 U677 ( .A(KEYINPUT65), .B(n595), .Z(n593) );
  NAND2_X1 U678 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U679 ( .A(KEYINPUT75), .B(n591), .ZN(n656) );
  NAND2_X1 U680 ( .A1(n656), .A2(n675), .ZN(n601) );
  INV_X1 U681 ( .A(n601), .ZN(n592) );
  NAND2_X1 U682 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U683 ( .A1(KEYINPUT47), .A2(n594), .ZN(n598) );
  NAND2_X1 U684 ( .A1(KEYINPUT65), .A2(n595), .ZN(n596) );
  AND2_X1 U685 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U686 ( .A1(KEYINPUT69), .A2(n601), .ZN(n611) );
  NOR2_X1 U687 ( .A1(n671), .A2(n602), .ZN(n604) );
  NOR2_X1 U688 ( .A1(n682), .A2(n659), .ZN(n603) );
  NAND2_X1 U689 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U690 ( .A1(n606), .A2(n605), .ZN(n622) );
  NAND2_X1 U691 ( .A1(n622), .A2(n607), .ZN(n609) );
  NAND2_X1 U692 ( .A1(n610), .A2(n686), .ZN(n667) );
  NAND2_X1 U693 ( .A1(n611), .A2(n667), .ZN(n618) );
  NAND2_X1 U694 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U695 ( .A1(n567), .A2(n614), .ZN(n615) );
  NAND2_X1 U696 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U697 ( .A(KEYINPUT105), .B(n617), .ZN(n751) );
  NOR2_X1 U698 ( .A1(n618), .A2(n751), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U700 ( .A(n624), .B(KEYINPUT43), .ZN(n625) );
  NAND2_X1 U701 ( .A1(n625), .A2(n567), .ZN(n669) );
  XNOR2_X1 U702 ( .A(n743), .B(KEYINPUT71), .ZN(n627) );
  INV_X1 U703 ( .A(KEYINPUT2), .ZN(n670) );
  NAND2_X1 U704 ( .A1(n429), .A2(G472), .ZN(n629) );
  INV_X1 U705 ( .A(KEYINPUT60), .ZN(n635) );
  XOR2_X1 U706 ( .A(KEYINPUT121), .B(KEYINPUT59), .Z(n630) );
  XNOR2_X1 U707 ( .A(n633), .B(n632), .ZN(n634) );
  NAND2_X1 U708 ( .A1(n429), .A2(G469), .ZN(n638) );
  XNOR2_X1 U709 ( .A(n638), .B(n637), .ZN(n639) );
  NAND2_X1 U710 ( .A1(n639), .A2(n368), .ZN(n641) );
  INV_X1 U711 ( .A(KEYINPUT120), .ZN(n640) );
  XNOR2_X1 U712 ( .A(n641), .B(n640), .ZN(G54) );
  XNOR2_X1 U713 ( .A(n355), .B(G101), .ZN(G3) );
  NOR2_X1 U714 ( .A1(n659), .A2(n644), .ZN(n643) );
  XOR2_X1 U715 ( .A(G104), .B(n643), .Z(G6) );
  NOR2_X1 U716 ( .A1(n664), .A2(n644), .ZN(n649) );
  XOR2_X1 U717 ( .A(KEYINPUT27), .B(KEYINPUT111), .Z(n646) );
  XNOR2_X1 U718 ( .A(G107), .B(KEYINPUT110), .ZN(n645) );
  XNOR2_X1 U719 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U720 ( .A(KEYINPUT26), .B(n647), .ZN(n648) );
  XNOR2_X1 U721 ( .A(n649), .B(n648), .ZN(G9) );
  XNOR2_X1 U722 ( .A(G110), .B(KEYINPUT112), .ZN(n651) );
  XNOR2_X1 U723 ( .A(n651), .B(n650), .ZN(G12) );
  XOR2_X1 U724 ( .A(G128), .B(KEYINPUT29), .Z(n654) );
  INV_X1 U725 ( .A(n664), .ZN(n652) );
  NAND2_X1 U726 ( .A1(n656), .A2(n652), .ZN(n653) );
  XNOR2_X1 U727 ( .A(n654), .B(n653), .ZN(G30) );
  XOR2_X1 U728 ( .A(G146), .B(KEYINPUT113), .Z(n658) );
  NAND2_X1 U729 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U730 ( .A(n658), .B(n657), .ZN(G48) );
  NOR2_X1 U731 ( .A1(n659), .A2(n663), .ZN(n661) );
  XNOR2_X1 U732 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n660) );
  XNOR2_X1 U733 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U734 ( .A(G113), .B(n662), .ZN(G15) );
  NOR2_X1 U735 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U736 ( .A(G116), .B(n665), .Z(G18) );
  XOR2_X1 U737 ( .A(G125), .B(KEYINPUT37), .Z(n666) );
  XNOR2_X1 U738 ( .A(n667), .B(n666), .ZN(G27) );
  XOR2_X1 U739 ( .A(G134), .B(n668), .Z(G36) );
  XNOR2_X1 U740 ( .A(G140), .B(n669), .ZN(G42) );
  NAND2_X1 U741 ( .A1(n672), .A2(n671), .ZN(n674) );
  NAND2_X1 U742 ( .A1(n674), .A2(n673), .ZN(n679) );
  NAND2_X1 U743 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U744 ( .A(KEYINPUT117), .B(n677), .Z(n678) );
  NAND2_X1 U745 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U746 ( .A(KEYINPUT118), .B(n680), .Z(n681) );
  NOR2_X1 U747 ( .A1(n704), .A2(n681), .ZN(n697) );
  NOR2_X1 U748 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U749 ( .A(n684), .B(KEYINPUT49), .ZN(n685) );
  NAND2_X1 U750 ( .A1(n544), .A2(n685), .ZN(n689) );
  NOR2_X1 U751 ( .A1(n357), .A2(n686), .ZN(n687) );
  XNOR2_X1 U752 ( .A(n687), .B(KEYINPUT50), .ZN(n688) );
  NOR2_X1 U753 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U754 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U755 ( .A(KEYINPUT51), .B(n692), .ZN(n694) );
  NAND2_X1 U756 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U757 ( .A(KEYINPUT116), .B(n695), .Z(n696) );
  NOR2_X1 U758 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U759 ( .A(KEYINPUT52), .B(n698), .Z(n700) );
  NAND2_X1 U760 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U761 ( .A1(n702), .A2(n701), .ZN(n708) );
  NOR2_X1 U762 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U763 ( .A(n705), .B(KEYINPUT119), .ZN(n706) );
  NAND2_X1 U764 ( .A1(n745), .A2(n706), .ZN(n707) );
  NOR2_X1 U765 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U766 ( .A(n709), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U767 ( .A1(n429), .A2(G210), .ZN(n712) );
  XOR2_X1 U768 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n711) );
  NAND2_X1 U769 ( .A1(G478), .A2(n429), .ZN(n713) );
  XNOR2_X1 U770 ( .A(n714), .B(n713), .ZN(n715) );
  NOR2_X1 U771 ( .A1(n720), .A2(n715), .ZN(G63) );
  XNOR2_X1 U772 ( .A(n716), .B(KEYINPUT122), .ZN(n718) );
  NAND2_X1 U773 ( .A1(G217), .A2(n429), .ZN(n717) );
  XNOR2_X1 U774 ( .A(n718), .B(n717), .ZN(n719) );
  NOR2_X1 U775 ( .A1(n720), .A2(n719), .ZN(G66) );
  XNOR2_X1 U776 ( .A(n722), .B(n721), .ZN(n723) );
  XNOR2_X1 U777 ( .A(n723), .B(KEYINPUT124), .ZN(n724) );
  XNOR2_X1 U778 ( .A(n724), .B(G101), .ZN(n725) );
  NOR2_X1 U779 ( .A1(n726), .A2(n725), .ZN(n734) );
  XOR2_X1 U780 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n728) );
  NAND2_X1 U781 ( .A1(G224), .A2(G953), .ZN(n727) );
  XNOR2_X1 U782 ( .A(n728), .B(n727), .ZN(n729) );
  NAND2_X1 U783 ( .A1(n729), .A2(G898), .ZN(n732) );
  NAND2_X1 U784 ( .A1(n730), .A2(n745), .ZN(n731) );
  NAND2_X1 U785 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U786 ( .A(n734), .B(n733), .ZN(G69) );
  XOR2_X1 U787 ( .A(n736), .B(n735), .Z(n737) );
  XNOR2_X1 U788 ( .A(n738), .B(n737), .ZN(n744) );
  XNOR2_X1 U789 ( .A(G227), .B(n744), .ZN(n739) );
  NAND2_X1 U790 ( .A1(n739), .A2(G900), .ZN(n740) );
  XOR2_X1 U791 ( .A(KEYINPUT125), .B(n740), .Z(n741) );
  NAND2_X1 U792 ( .A1(G953), .A2(n741), .ZN(n742) );
  XNOR2_X1 U793 ( .A(n742), .B(KEYINPUT126), .ZN(n748) );
  XNOR2_X1 U794 ( .A(n744), .B(n743), .ZN(n746) );
  NAND2_X1 U795 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U796 ( .A1(n748), .A2(n747), .ZN(G72) );
  XNOR2_X1 U797 ( .A(n749), .B(G131), .ZN(G33) );
  XOR2_X1 U798 ( .A(n750), .B(G122), .Z(G24) );
  XOR2_X1 U799 ( .A(n354), .B(n751), .Z(G45) );
  XNOR2_X1 U800 ( .A(G119), .B(n752), .ZN(G21) );
  XNOR2_X1 U801 ( .A(G137), .B(n753), .ZN(G39) );
endmodule

