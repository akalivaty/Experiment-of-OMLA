//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 0 0 1 0 0 0 1 0 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 1 0 1 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n955, new_n956, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1008, new_n1009, new_n1010, new_n1011, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1018, new_n1019, new_n1020;
  INV_X1    g000(.A(KEYINPUT15), .ZN(new_n202));
  OR2_X1    g001(.A1(G43gat), .A2(G50gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(G43gat), .A2(G50gat), .ZN(new_n204));
  AOI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G29gat), .ZN(new_n206));
  INV_X1    g005(.A(G36gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT14), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT14), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n209), .B1(G29gat), .B2(G36gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n210), .A3(KEYINPUT89), .ZN(new_n211));
  NAND2_X1  g010(.A1(G29gat), .A2(G36gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT89), .B1(new_n208), .B2(new_n210), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n205), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n205), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n208), .A2(new_n210), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n203), .A2(new_n202), .A3(new_n204), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n216), .A2(new_n217), .A3(new_n212), .A4(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT17), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G8gat), .ZN(new_n223));
  INV_X1    g022(.A(G15gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G22gat), .ZN(new_n225));
  INV_X1    g024(.A(G22gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G15gat), .ZN(new_n227));
  AOI21_X1  g026(.A(G1gat), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G1gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT16), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n231), .A2(new_n225), .A3(new_n227), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n223), .B1(new_n229), .B2(new_n232), .ZN(new_n233));
  AND3_X1   g032(.A1(new_n231), .A2(new_n225), .A3(new_n227), .ZN(new_n234));
  NOR3_X1   g033(.A1(new_n234), .A2(new_n228), .A3(G8gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n215), .A2(KEYINPUT17), .A3(new_n219), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n222), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT90), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT91), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(new_n233), .B2(new_n235), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n229), .A2(new_n232), .A3(new_n223), .ZN(new_n242));
  OAI21_X1  g041(.A(G8gat), .B1(new_n234), .B2(new_n228), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n242), .A2(new_n243), .A3(KEYINPUT91), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n241), .A2(new_n220), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT90), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n222), .A2(new_n246), .A3(new_n236), .A4(new_n237), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT18), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n248), .B1(G229gat), .B2(G233gat), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n239), .A2(new_n245), .A3(new_n247), .A4(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT92), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n247), .A2(new_n245), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n253), .A2(KEYINPUT92), .A3(new_n239), .A4(new_n249), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G229gat), .A2(G233gat), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n239), .A2(new_n245), .A3(new_n247), .A4(new_n256), .ZN(new_n257));
  XOR2_X1   g056(.A(new_n256), .B(KEYINPUT13), .Z(new_n258));
  AND3_X1   g057(.A1(new_n241), .A2(new_n220), .A3(new_n244), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n220), .B1(new_n241), .B2(new_n244), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT93), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI211_X1 g062(.A(KEYINPUT93), .B(new_n258), .C1(new_n259), .C2(new_n260), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n257), .A2(new_n248), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G113gat), .B(G141gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(G169gat), .B(G197gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  XOR2_X1   g067(.A(KEYINPUT88), .B(KEYINPUT11), .Z(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT12), .ZN(new_n271));
  AND3_X1   g070(.A1(new_n255), .A2(new_n265), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n271), .B1(new_n255), .B2(new_n265), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AND2_X1   g073(.A1(G232gat), .A2(G233gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n275), .A2(KEYINPUT41), .ZN(new_n276));
  XNOR2_X1  g075(.A(G134gat), .B(G162gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT101), .ZN(new_n279));
  AND3_X1   g078(.A1(KEYINPUT99), .A2(G85gat), .A3(G92gat), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT99), .B1(G85gat), .B2(G92gat), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT7), .ZN(new_n282));
  OAI22_X1  g081(.A1(new_n280), .A2(new_n281), .B1(KEYINPUT98), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G85gat), .A2(G92gat), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT99), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n282), .A2(KEYINPUT98), .ZN(new_n287));
  NAND3_X1  g086(.A1(KEYINPUT99), .A2(G85gat), .A3(G92gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G99gat), .A2(G106gat), .ZN(new_n290));
  INV_X1    g089(.A(G85gat), .ZN(new_n291));
  INV_X1    g090(.A(G92gat), .ZN(new_n292));
  AOI22_X1  g091(.A1(KEYINPUT8), .A2(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n283), .A2(new_n289), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n290), .ZN(new_n295));
  NOR2_X1   g094(.A1(G99gat), .A2(G106gat), .ZN(new_n296));
  OAI21_X1  g095(.A(KEYINPUT100), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OR2_X1    g096(.A1(G99gat), .A2(G106gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT100), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n299), .A3(new_n290), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n294), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n294), .A2(new_n301), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n279), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n297), .A2(new_n300), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n305), .A2(new_n289), .A3(new_n283), .A4(new_n293), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n294), .A2(new_n301), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n306), .A2(KEYINPUT101), .A3(new_n307), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n222), .A2(new_n304), .A3(new_n237), .A4(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n306), .A2(new_n307), .ZN(new_n310));
  AOI22_X1  g109(.A1(new_n310), .A2(new_n220), .B1(KEYINPUT41), .B2(new_n275), .ZN(new_n311));
  XNOR2_X1  g110(.A(G190gat), .B(G218gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n309), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n312), .B1(new_n309), .B2(new_n311), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n278), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n309), .A2(new_n311), .ZN(new_n317));
  INV_X1    g116(.A(new_n312), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n278), .B(KEYINPUT97), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n319), .A2(new_n313), .A3(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n316), .A2(new_n321), .A3(KEYINPUT102), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT102), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n319), .A2(new_n323), .A3(new_n313), .A4(new_n320), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  AND2_X1   g124(.A1(G71gat), .A2(G78gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(G71gat), .A2(G78gat), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT94), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G71gat), .ZN(new_n329));
  INV_X1    g128(.A(G78gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT94), .ZN(new_n332));
  NAND2_X1  g131(.A1(G71gat), .A2(G78gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G57gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G64gat), .ZN(new_n336));
  INV_X1    g135(.A(G64gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(G57gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n333), .A2(new_n340), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n328), .A2(new_n334), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT96), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n343), .B1(new_n326), .B2(new_n327), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n331), .A2(KEYINPUT96), .A3(new_n333), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n344), .A2(new_n345), .A3(new_n341), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT95), .B1(new_n335), .B2(G64gat), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT95), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n348), .A2(new_n337), .A3(G57gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n347), .A2(new_n349), .A3(new_n336), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n342), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n351), .B1(new_n302), .B2(new_n303), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT10), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n328), .A2(new_n334), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n341), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n350), .A2(new_n341), .A3(new_n345), .A4(new_n344), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n306), .A2(new_n358), .A3(new_n307), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n352), .A2(new_n353), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n310), .A2(KEYINPUT10), .A3(new_n351), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(G230gat), .A2(G233gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(G120gat), .B(G148gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(G176gat), .B(G204gat), .ZN(new_n366));
  XOR2_X1   g165(.A(new_n365), .B(new_n366), .Z(new_n367));
  AND2_X1   g166(.A1(new_n352), .A2(new_n359), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n364), .B(new_n367), .C1(new_n368), .C2(new_n363), .ZN(new_n369));
  INV_X1    g168(.A(new_n367), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n368), .A2(new_n363), .ZN(new_n371));
  INV_X1    g170(.A(new_n363), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n372), .B1(new_n360), .B2(new_n361), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n370), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n377));
  INV_X1    g176(.A(G155gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G183gat), .B(G211gat), .ZN(new_n380));
  XOR2_X1   g179(.A(new_n379), .B(new_n380), .Z(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT21), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n358), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n384), .A2(G231gat), .A3(G233gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(G231gat), .A2(G233gat), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n358), .A2(new_n383), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(G127gat), .ZN(new_n389));
  INV_X1    g188(.A(G127gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n385), .A2(new_n390), .A3(new_n387), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n241), .A2(new_n244), .B1(new_n351), .B2(KEYINPUT21), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n389), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n393), .B1(new_n389), .B2(new_n391), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n382), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n396), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n398), .A2(new_n394), .A3(new_n381), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n325), .A2(new_n376), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(G134gat), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n402), .A2(G127gat), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n390), .A2(G134gat), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT68), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(G120gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(G113gat), .ZN(new_n407));
  INV_X1    g206(.A(G113gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(G120gat), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT1), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n390), .A2(G134gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n402), .A2(G127gat), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT68), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n405), .A2(new_n410), .A3(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n411), .A2(new_n412), .A3(KEYINPUT67), .ZN(new_n416));
  OR3_X1    g215(.A1(new_n402), .A2(KEYINPUT67), .A3(G127gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(G113gat), .B(G120gat), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n416), .B(new_n417), .C1(KEYINPUT1), .C2(new_n418), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(G183gat), .A2(G190gat), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT24), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(G183gat), .ZN(new_n424));
  INV_X1    g223(.A(G190gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n423), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT64), .ZN(new_n429));
  NOR2_X1   g228(.A1(G169gat), .A2(G176gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT23), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT23), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n432), .B1(G169gat), .B2(G176gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(G169gat), .A2(G176gat), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n431), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT64), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n423), .A2(new_n426), .A3(new_n436), .A4(new_n427), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n429), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT25), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT65), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n421), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n422), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n421), .A2(new_n440), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n426), .B(new_n427), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n431), .A2(new_n433), .A3(new_n434), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n445), .A2(new_n439), .ZN(new_n446));
  AOI22_X1  g245(.A1(new_n438), .A2(new_n439), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n430), .A2(KEYINPUT26), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n421), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT26), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n451), .A2(new_n430), .ZN(new_n452));
  OR2_X1    g251(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT28), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT27), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(G183gat), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT66), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n425), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n424), .A2(KEYINPUT27), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT66), .B1(new_n456), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n454), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n456), .A2(new_n459), .A3(KEYINPUT28), .A4(new_n425), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n453), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n420), .B1(new_n447), .B2(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n449), .A2(new_n452), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n456), .A2(new_n459), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT66), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(G190gat), .B1(new_n456), .B2(KEYINPUT66), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT28), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n462), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n465), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n415), .A2(new_n419), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n445), .B1(KEYINPUT64), .B2(new_n428), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT25), .B1(new_n474), .B2(new_n437), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n446), .A2(new_n444), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n472), .B(new_n473), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(G227gat), .A2(G233gat), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n464), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  XOR2_X1   g279(.A(G71gat), .B(G99gat), .Z(new_n481));
  XNOR2_X1  g280(.A(G15gat), .B(G43gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n481), .B(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(KEYINPUT69), .B(KEYINPUT33), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n480), .A2(KEYINPUT32), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT70), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT70), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n480), .A2(new_n489), .A3(KEYINPUT32), .A4(new_n486), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n479), .B1(new_n464), .B2(new_n477), .ZN(new_n492));
  NAND2_X1  g291(.A1(KEYINPUT71), .A2(KEYINPUT34), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(KEYINPUT71), .A2(KEYINPUT34), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  AOI211_X1 g296(.A(new_n479), .B(new_n494), .C1(new_n464), .C2(new_n477), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT72), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n480), .A2(KEYINPUT32), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n480), .A2(new_n484), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n500), .A2(new_n501), .A3(new_n483), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n491), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  OR3_X1    g302(.A1(new_n497), .A2(new_n498), .A3(KEYINPUT72), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n504), .A2(new_n491), .A3(new_n499), .A4(new_n502), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n506), .A2(KEYINPUT73), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT36), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT36), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n506), .A2(KEYINPUT73), .A3(new_n510), .A4(new_n507), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(G8gat), .B(G36gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(G64gat), .B(G92gat), .ZN(new_n514));
  XOR2_X1   g313(.A(new_n513), .B(new_n514), .Z(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(G226gat), .A2(G233gat), .ZN(new_n517));
  XOR2_X1   g316(.A(new_n517), .B(KEYINPUT74), .Z(new_n518));
  OAI21_X1  g317(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT29), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n438), .A2(new_n439), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n446), .A2(new_n444), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n461), .A2(new_n462), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n522), .A2(new_n523), .B1(new_n524), .B2(new_n465), .ZN(new_n525));
  XOR2_X1   g324(.A(new_n518), .B(KEYINPUT75), .Z(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G197gat), .B(G204gat), .ZN(new_n529));
  AND2_X1   g328(.A1(G211gat), .A2(G218gat), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n529), .B1(KEYINPUT22), .B2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G211gat), .B(G218gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NOR3_X1   g332(.A1(new_n521), .A2(new_n528), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n533), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n527), .B1(new_n525), .B2(KEYINPUT29), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n518), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n516), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n536), .A2(new_n537), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(new_n533), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n519), .A2(new_n526), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n525), .A2(KEYINPUT29), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n535), .B(new_n542), .C1(new_n543), .C2(new_n518), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n541), .A2(new_n544), .A3(new_n515), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n539), .A2(new_n545), .A3(KEYINPUT30), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT30), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n541), .A2(new_n547), .A3(new_n544), .A4(new_n515), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(G225gat), .A2(G233gat), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT79), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n473), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G155gat), .A2(G162gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT2), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT78), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n554), .A2(KEYINPUT78), .A3(KEYINPUT2), .ZN(new_n558));
  XNOR2_X1  g357(.A(G155gat), .B(G162gat), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(G148gat), .ZN(new_n561));
  NOR3_X1   g360(.A1(new_n561), .A2(KEYINPUT77), .A3(G141gat), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(G141gat), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT77), .ZN(new_n565));
  INV_X1    g364(.A(G141gat), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n565), .B1(new_n566), .B2(G148gat), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n562), .B1(new_n564), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n561), .A2(G141gat), .ZN(new_n569));
  AOI21_X1  g368(.A(KEYINPUT2), .B1(new_n564), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(G162gat), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n378), .A2(new_n571), .A3(KEYINPUT76), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT76), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n573), .B1(G155gat), .B2(G162gat), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n572), .A2(new_n574), .A3(new_n554), .ZN(new_n575));
  OAI22_X1  g374(.A1(new_n560), .A2(new_n568), .B1(new_n570), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n415), .A2(new_n419), .A3(KEYINPUT79), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n553), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n578), .A2(KEYINPUT81), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT81), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n553), .A2(new_n580), .A3(new_n576), .A4(new_n577), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n565), .A2(new_n566), .A3(G148gat), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT77), .B1(new_n561), .B2(G141gat), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n582), .B1(new_n583), .B2(new_n563), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n584), .A2(new_n557), .A3(new_n558), .A4(new_n559), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT2), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n566), .A2(G148gat), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n586), .B1(new_n563), .B2(new_n587), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n588), .A2(new_n554), .A3(new_n572), .A4(new_n574), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n585), .A2(new_n589), .A3(new_n419), .A4(new_n415), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n581), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n551), .B1(new_n579), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n576), .A2(KEYINPUT3), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT3), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n585), .A2(new_n589), .A3(new_n594), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n593), .A2(new_n553), .A3(new_n577), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(new_n550), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n420), .A2(KEYINPUT4), .A3(new_n585), .A4(new_n589), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT4), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n590), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(KEYINPUT80), .B1(new_n597), .B2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n590), .B(KEYINPUT4), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT80), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n603), .A2(new_n604), .A3(new_n550), .A4(new_n596), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n592), .A2(new_n602), .A3(KEYINPUT5), .A4(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(G1gat), .B(G29gat), .Z(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G57gat), .B(G85gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n603), .A2(KEYINPUT83), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT83), .B1(new_n598), .B2(new_n600), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n597), .A2(KEYINPUT5), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AND3_X1   g416(.A1(new_n606), .A2(new_n611), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n611), .B1(new_n606), .B2(new_n617), .ZN(new_n619));
  NOR3_X1   g418(.A1(new_n618), .A2(new_n619), .A3(KEYINPUT6), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n606), .A2(new_n617), .ZN(new_n621));
  INV_X1    g420(.A(new_n611), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n621), .A2(KEYINPUT6), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n549), .B1(new_n620), .B2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(KEYINPUT31), .B(G50gat), .ZN(new_n626));
  INV_X1    g425(.A(G228gat), .ZN(new_n627));
  INV_X1    g426(.A(G233gat), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n595), .A2(new_n520), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(KEYINPUT84), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT84), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n595), .A2(new_n633), .A3(new_n520), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n632), .A2(new_n533), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n594), .B1(new_n533), .B2(KEYINPUT29), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n576), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n630), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n631), .A2(new_n533), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n637), .A2(new_n630), .A3(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n626), .B1(new_n638), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n634), .A2(new_n533), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n633), .B1(new_n595), .B2(new_n520), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n637), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n629), .ZN(new_n646));
  INV_X1    g445(.A(new_n626), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n646), .A2(new_n640), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(G78gat), .B(G106gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(G22gat), .ZN(new_n650));
  AND3_X1   g449(.A1(new_n642), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n650), .B1(new_n642), .B2(new_n648), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n625), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n623), .A2(KEYINPUT86), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT86), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n619), .A2(new_n657), .A3(KEYINPUT6), .ZN(new_n658));
  OAI21_X1  g457(.A(KEYINPUT37), .B1(new_n534), .B2(new_n538), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n516), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT37), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n541), .A2(new_n661), .A3(new_n544), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(KEYINPUT85), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT85), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n541), .A2(new_n664), .A3(new_n661), .A4(new_n544), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n660), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT38), .ZN(new_n667));
  OAI211_X1 g466(.A(new_n656), .B(new_n658), .C1(new_n666), .C2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n621), .A2(new_n622), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT6), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n606), .A2(new_n611), .A3(new_n617), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n663), .A2(new_n665), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n661), .B1(new_n540), .B2(new_n535), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n533), .B(new_n542), .C1(new_n543), .C2(new_n518), .ZN(new_n675));
  AOI211_X1 g474(.A(KEYINPUT38), .B(new_n515), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n672), .A2(new_n677), .A3(new_n545), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n668), .A2(new_n678), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n598), .A2(new_n600), .A3(KEYINPUT83), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n596), .B1(new_n680), .B2(new_n613), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT39), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n681), .A2(new_n682), .A3(new_n551), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n683), .A2(new_n611), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n681), .A2(new_n551), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n578), .A2(KEYINPUT81), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n686), .A2(new_n590), .A3(new_n581), .ZN(new_n687));
  OAI21_X1  g486(.A(KEYINPUT39), .B1(new_n687), .B2(new_n551), .ZN(new_n688));
  OAI211_X1 g487(.A(new_n684), .B(KEYINPUT40), .C1(new_n685), .C2(new_n688), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n611), .B(new_n683), .C1(new_n685), .C2(new_n688), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT40), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n689), .A2(new_n692), .A3(new_n669), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n653), .B1(new_n693), .B2(new_n549), .ZN(new_n694));
  OAI211_X1 g493(.A(new_n512), .B(new_n655), .C1(new_n679), .C2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n507), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n492), .A2(new_n493), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n697), .B1(new_n492), .B2(new_n496), .ZN(new_n698));
  AOI211_X1 g497(.A(KEYINPUT72), .B(new_n698), .C1(new_n491), .C2(new_n502), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n653), .B1(new_n696), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(KEYINPUT35), .B1(new_n625), .B2(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT35), .B1(new_n546), .B2(new_n548), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n653), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n672), .A2(new_n656), .A3(new_n658), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n506), .A2(KEYINPUT87), .A3(new_n507), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT87), .B1(new_n506), .B2(new_n507), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n703), .B(new_n704), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n701), .A2(new_n707), .ZN(new_n708));
  AOI211_X1 g507(.A(new_n274), .B(new_n401), .C1(new_n695), .C2(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n620), .A2(new_n624), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT103), .B(G1gat), .Z(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1324gat));
  INV_X1    g512(.A(new_n549), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n709), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g514(.A(KEYINPUT16), .B(G8gat), .Z(new_n716));
  AND2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n715), .A2(new_n223), .ZN(new_n718));
  OAI21_X1  g517(.A(KEYINPUT42), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(KEYINPUT42), .B2(new_n717), .ZN(G1325gat));
  NOR2_X1   g519(.A1(new_n705), .A2(new_n706), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n709), .A2(new_n224), .A3(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n512), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n709), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n723), .B1(new_n725), .B2(new_n224), .ZN(G1326gat));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n654), .ZN(new_n727));
  XNOR2_X1  g526(.A(KEYINPUT43), .B(G22gat), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1327gat));
  NAND2_X1  g528(.A1(new_n695), .A2(new_n708), .ZN(new_n730));
  INV_X1    g529(.A(new_n325), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n274), .A2(new_n400), .A3(new_n375), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n735), .A2(new_n206), .A3(new_n710), .ZN(new_n736));
  XOR2_X1   g535(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT107), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n740));
  NAND2_X1  g539(.A1(new_n731), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT106), .B1(new_n730), .B2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n744), .B1(new_n730), .B2(new_n731), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT106), .ZN(new_n746));
  AOI211_X1 g545(.A(new_n746), .B(new_n741), .C1(new_n695), .C2(new_n708), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n743), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n739), .B1(new_n748), .B2(new_n734), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n730), .A2(new_n742), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n746), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n732), .A2(KEYINPUT44), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n730), .A2(KEYINPUT106), .A3(new_n742), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n751), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n754), .A2(KEYINPUT107), .A3(new_n733), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n749), .A2(new_n710), .A3(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n738), .B1(new_n756), .B2(new_n206), .ZN(G1328gat));
  NAND3_X1  g556(.A1(new_n749), .A2(new_n714), .A3(new_n755), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(KEYINPUT108), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT108), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n749), .A2(new_n755), .A3(new_n760), .A4(new_n714), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n759), .A2(G36gat), .A3(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n735), .A2(new_n207), .A3(new_n714), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n763), .B(KEYINPUT46), .Z(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(G1329gat));
  NOR4_X1   g564(.A1(new_n732), .A2(G43gat), .A3(new_n721), .A4(new_n734), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n749), .A2(new_n724), .A3(new_n755), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n766), .B1(new_n767), .B2(G43gat), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n754), .A2(new_n724), .A3(new_n733), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n769), .A2(G43gat), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT47), .ZN(new_n771));
  OR2_X1    g570(.A1(new_n766), .A2(new_n771), .ZN(new_n772));
  OAI22_X1  g571(.A1(new_n768), .A2(KEYINPUT47), .B1(new_n770), .B2(new_n772), .ZN(G1330gat));
  NAND3_X1  g572(.A1(new_n749), .A2(new_n654), .A3(new_n755), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n653), .A2(G50gat), .ZN(new_n775));
  AOI22_X1  g574(.A1(new_n774), .A2(G50gat), .B1(new_n735), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n735), .A2(new_n775), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT48), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n754), .A2(new_n654), .A3(new_n733), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n778), .B1(new_n779), .B2(G50gat), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT109), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI211_X1 g581(.A(KEYINPUT109), .B(new_n778), .C1(new_n779), .C2(G50gat), .ZN(new_n783));
  OAI22_X1  g582(.A1(new_n776), .A2(KEYINPUT48), .B1(new_n782), .B2(new_n783), .ZN(G1331gat));
  INV_X1    g583(.A(new_n400), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n731), .A2(new_n785), .A3(new_n376), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n730), .A2(new_n274), .A3(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n710), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(new_n335), .ZN(G1332gat));
  NOR2_X1   g589(.A1(new_n787), .A2(new_n549), .ZN(new_n791));
  NOR2_X1   g590(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n792));
  AND2_X1   g591(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n794), .B1(new_n791), .B2(new_n792), .ZN(G1333gat));
  INV_X1    g594(.A(new_n787), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT87), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n797), .B1(new_n696), .B2(new_n699), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n506), .A2(KEYINPUT87), .A3(new_n507), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n798), .A2(KEYINPUT110), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT110), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n801), .B1(new_n705), .B2(new_n706), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n796), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n724), .A2(G71gat), .ZN(new_n804));
  OAI22_X1  g603(.A1(new_n803), .A2(G71gat), .B1(new_n787), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g605(.A1(new_n787), .A2(new_n653), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(new_n330), .ZN(G1335gat));
  INV_X1    g607(.A(KEYINPUT111), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n732), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n255), .A2(new_n265), .ZN(new_n811));
  INV_X1    g610(.A(new_n271), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n255), .A2(new_n265), .A3(new_n271), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n815), .A2(new_n400), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n325), .B1(new_n695), .B2(new_n708), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n817), .B1(new_n818), .B2(KEYINPUT111), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n810), .A2(new_n819), .A3(KEYINPUT51), .ZN(new_n820));
  AOI21_X1  g619(.A(KEYINPUT51), .B1(new_n810), .B2(new_n819), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n822), .A2(new_n291), .A3(new_n710), .A4(new_n375), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n817), .A2(new_n376), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n754), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(G85gat), .B1(new_n825), .B2(new_n788), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n823), .A2(new_n826), .ZN(G1336gat));
  INV_X1    g626(.A(KEYINPUT52), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n714), .A2(new_n292), .A3(new_n375), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(KEYINPUT113), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n830), .B1(new_n820), .B2(new_n821), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT112), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n828), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(G92gat), .B1(new_n825), .B2(new_n549), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n831), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n834), .B(new_n831), .C1(new_n832), .C2(new_n828), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(G1337gat));
  NOR3_X1   g637(.A1(new_n721), .A2(G99gat), .A3(new_n376), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n822), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(G99gat), .B1(new_n825), .B2(new_n512), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(G1338gat));
  OAI21_X1  g641(.A(G106gat), .B1(new_n825), .B2(new_n653), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n653), .A2(G106gat), .A3(new_n376), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n844), .B1(new_n820), .B2(new_n821), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g645(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n846), .B(new_n847), .ZN(G1339gat));
  INV_X1    g647(.A(KEYINPUT55), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n360), .A2(new_n361), .A3(new_n372), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT54), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n850), .A2(new_n373), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n362), .A2(new_n851), .A3(new_n363), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n370), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n849), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n360), .A2(new_n361), .A3(new_n372), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n364), .A2(KEYINPUT54), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n367), .B1(new_n373), .B2(new_n851), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(KEYINPUT55), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n855), .A2(new_n369), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n860), .B1(new_n813), .B2(new_n814), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n256), .B1(new_n253), .B2(new_n239), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n259), .A2(new_n260), .A3(new_n258), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n270), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n814), .A2(new_n375), .A3(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n325), .B1(new_n861), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n814), .A2(new_n864), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n868), .A2(new_n860), .A3(new_n325), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n400), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  AND3_X1   g670(.A1(new_n325), .A2(new_n376), .A3(new_n400), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT115), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n872), .A2(new_n873), .A3(new_n274), .ZN(new_n874));
  OAI21_X1  g673(.A(KEYINPUT115), .B1(new_n815), .B2(new_n401), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n871), .A2(new_n876), .A3(KEYINPUT116), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT116), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n859), .A2(new_n369), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n879), .B(new_n855), .C1(new_n272), .C2(new_n273), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n731), .B1(new_n880), .B2(new_n865), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n785), .B1(new_n881), .B2(new_n869), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n874), .A2(new_n875), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n878), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n877), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n788), .A2(new_n714), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n885), .A2(new_n653), .A3(new_n722), .A4(new_n886), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n887), .A2(new_n408), .A3(new_n274), .ZN(new_n888));
  OAI21_X1  g687(.A(KEYINPUT116), .B1(new_n871), .B2(new_n876), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n882), .A2(new_n878), .A3(new_n883), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OR3_X1    g690(.A1(new_n891), .A2(new_n788), .A3(new_n700), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n892), .A2(KEYINPUT117), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n714), .B1(new_n892), .B2(KEYINPUT117), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n815), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n888), .B1(new_n897), .B2(new_n408), .ZN(G1340gat));
  NOR3_X1   g697(.A1(new_n887), .A2(new_n406), .A3(new_n376), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n896), .A2(new_n375), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(new_n406), .ZN(G1341gat));
  NOR3_X1   g700(.A1(new_n887), .A2(new_n390), .A3(new_n785), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT118), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n902), .B(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n896), .A2(new_n400), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n904), .B1(new_n905), .B2(new_n390), .ZN(G1342gat));
  NOR2_X1   g705(.A1(new_n325), .A2(G134gat), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  OR3_X1    g707(.A1(new_n895), .A2(KEYINPUT56), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(G134gat), .B1(new_n887), .B2(new_n325), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT56), .B1(new_n895), .B2(new_n908), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(G1343gat));
  NAND2_X1  g711(.A1(new_n886), .A2(new_n512), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT57), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n914), .B1(new_n891), .B2(new_n653), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT119), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n916), .B1(new_n852), .B2(new_n854), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n857), .A2(KEYINPUT119), .A3(new_n858), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n917), .A2(new_n918), .A3(new_n849), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(new_n879), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n865), .B1(new_n274), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(new_n325), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n400), .B1(new_n922), .B2(new_n870), .ZN(new_n923));
  OAI211_X1 g722(.A(KEYINPUT57), .B(new_n654), .C1(new_n923), .C2(new_n876), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n913), .B1(new_n915), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(new_n815), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(G141gat), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT120), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n724), .A2(new_n714), .A3(new_n653), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n885), .A2(new_n710), .A3(new_n930), .ZN(new_n931));
  OR3_X1    g730(.A1(new_n931), .A2(G141gat), .A3(new_n274), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n927), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n929), .A2(new_n933), .A3(KEYINPUT58), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT58), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n927), .B(new_n932), .C1(new_n928), .C2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(G1344gat));
  INV_X1    g736(.A(KEYINPUT59), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n376), .B1(new_n913), .B2(KEYINPUT121), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n815), .A2(new_n401), .ZN(new_n940));
  OR2_X1    g739(.A1(new_n923), .A2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT122), .ZN(new_n942));
  OR2_X1    g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n653), .B1(new_n941), .B2(new_n942), .ZN(new_n944));
  AOI21_X1  g743(.A(KEYINPUT57), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n891), .A2(new_n914), .A3(new_n653), .ZN(new_n946));
  OAI221_X1 g745(.A(new_n939), .B1(KEYINPUT121), .B2(new_n913), .C1(new_n945), .C2(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n938), .B1(new_n947), .B2(G148gat), .ZN(new_n948));
  AOI211_X1 g747(.A(KEYINPUT59), .B(new_n561), .C1(new_n925), .C2(new_n375), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n375), .A2(new_n561), .ZN(new_n950));
  OAI22_X1  g749(.A1(new_n948), .A2(new_n949), .B1(new_n931), .B2(new_n950), .ZN(G1345gat));
  AND2_X1   g750(.A1(new_n925), .A2(new_n400), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n400), .A2(new_n378), .ZN(new_n953));
  OAI22_X1  g752(.A1(new_n952), .A2(new_n378), .B1(new_n931), .B2(new_n953), .ZN(G1346gat));
  OR2_X1    g753(.A1(new_n931), .A2(new_n325), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n325), .A2(new_n571), .ZN(new_n956));
  AOI22_X1  g755(.A1(new_n955), .A2(new_n571), .B1(new_n925), .B2(new_n956), .ZN(G1347gat));
  OAI211_X1 g756(.A(new_n714), .B(new_n653), .C1(new_n696), .C2(new_n699), .ZN(new_n958));
  XOR2_X1   g757(.A(new_n958), .B(KEYINPUT123), .Z(new_n959));
  NAND4_X1  g758(.A1(new_n889), .A2(new_n890), .A3(new_n788), .A4(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(G169gat), .B1(new_n961), .B2(new_n815), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n710), .A2(new_n549), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n802), .A2(new_n800), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(KEYINPUT124), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT124), .ZN(new_n966));
  NAND4_X1  g765(.A1(new_n802), .A2(new_n800), .A3(new_n963), .A4(new_n966), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n968), .A2(new_n653), .A3(new_n889), .A4(new_n890), .ZN(new_n969));
  INV_X1    g768(.A(G169gat), .ZN(new_n970));
  NOR3_X1   g769(.A1(new_n969), .A2(new_n970), .A3(new_n274), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n962), .A2(new_n971), .ZN(G1348gat));
  OR3_X1    g771(.A1(new_n960), .A2(G176gat), .A3(new_n376), .ZN(new_n973));
  OAI21_X1  g772(.A(G176gat), .B1(new_n969), .B2(new_n376), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(G1349gat));
  OAI21_X1  g774(.A(G183gat), .B1(new_n969), .B2(new_n785), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n400), .A2(new_n456), .A3(new_n459), .ZN(new_n977));
  OR2_X1    g776(.A1(new_n960), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n976), .A2(new_n978), .A3(KEYINPUT126), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT125), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT60), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n960), .A2(new_n977), .ZN(new_n983));
  NAND4_X1  g782(.A1(new_n885), .A2(new_n653), .A3(new_n400), .A4(new_n968), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n983), .B1(new_n984), .B2(G183gat), .ZN(new_n985));
  AOI21_X1  g784(.A(KEYINPUT125), .B1(new_n985), .B2(KEYINPUT126), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n976), .A2(new_n978), .A3(KEYINPUT125), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n987), .A2(KEYINPUT60), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n982), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n989), .A2(KEYINPUT127), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT127), .ZN(new_n991));
  OAI211_X1 g790(.A(new_n991), .B(new_n982), .C1(new_n986), .C2(new_n988), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n990), .A2(new_n992), .ZN(G1350gat));
  OAI21_X1  g792(.A(G190gat), .B1(new_n969), .B2(new_n325), .ZN(new_n994));
  XNOR2_X1  g793(.A(new_n994), .B(KEYINPUT61), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n961), .A2(new_n425), .A3(new_n731), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(G1351gat));
  NOR2_X1   g796(.A1(new_n891), .A2(new_n710), .ZN(new_n998));
  NOR3_X1   g797(.A1(new_n724), .A2(new_n549), .A3(new_n653), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g799(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g800(.A(G197gat), .B1(new_n1001), .B2(new_n815), .ZN(new_n1002));
  OR2_X1    g801(.A1(new_n945), .A2(new_n946), .ZN(new_n1003));
  AND2_X1   g802(.A1(new_n512), .A2(new_n963), .ZN(new_n1004));
  AND2_X1   g803(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AND2_X1   g804(.A1(new_n815), .A2(G197gat), .ZN(new_n1006));
  AOI21_X1  g805(.A(new_n1002), .B1(new_n1005), .B2(new_n1006), .ZN(G1352gat));
  NAND3_X1  g806(.A1(new_n1003), .A2(new_n375), .A3(new_n1004), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1008), .A2(G204gat), .ZN(new_n1009));
  NOR3_X1   g808(.A1(new_n1000), .A2(G204gat), .A3(new_n376), .ZN(new_n1010));
  XNOR2_X1  g809(.A(new_n1010), .B(KEYINPUT62), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1009), .A2(new_n1011), .ZN(G1353gat));
  OR3_X1    g811(.A1(new_n1000), .A2(G211gat), .A3(new_n785), .ZN(new_n1013));
  OAI211_X1 g812(.A(new_n400), .B(new_n1004), .C1(new_n945), .C2(new_n946), .ZN(new_n1014));
  AND3_X1   g813(.A1(new_n1014), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1015));
  AOI21_X1  g814(.A(KEYINPUT63), .B1(new_n1014), .B2(G211gat), .ZN(new_n1016));
  OAI21_X1  g815(.A(new_n1013), .B1(new_n1015), .B2(new_n1016), .ZN(G1354gat));
  NAND3_X1  g816(.A1(new_n1003), .A2(new_n731), .A3(new_n1004), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n1018), .A2(G218gat), .ZN(new_n1019));
  OR2_X1    g818(.A1(new_n325), .A2(G218gat), .ZN(new_n1020));
  OAI21_X1  g819(.A(new_n1019), .B1(new_n1000), .B2(new_n1020), .ZN(G1355gat));
endmodule


