//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 1 1 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 0 0 0 1 0 1 1 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n835,
    new_n836, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944;
  INV_X1    g000(.A(KEYINPUT15), .ZN(new_n202));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(G29gat), .A2(G36gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT14), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n205), .B1(KEYINPUT91), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(KEYINPUT91), .B(KEYINPUT14), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n207), .B1(new_n208), .B2(new_n205), .ZN(new_n209));
  NAND2_X1  g008(.A1(G29gat), .A2(G36gat), .ZN(new_n210));
  AOI211_X1 g009(.A(new_n202), .B(new_n204), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  XOR2_X1   g010(.A(new_n209), .B(KEYINPUT93), .Z(new_n212));
  NAND3_X1  g011(.A1(new_n204), .A2(KEYINPUT92), .A3(new_n202), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT92), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT15), .B1(new_n203), .B2(new_n214), .ZN(new_n215));
  AND3_X1   g014(.A1(new_n213), .A2(new_n210), .A3(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n211), .B1(new_n212), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT17), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n217), .B(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G15gat), .B(G22gat), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n220), .A2(G1gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT16), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n220), .B1(new_n222), .B2(G1gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT94), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n221), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G8gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n224), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n221), .B(new_n223), .C1(new_n225), .C2(G8gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n219), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G229gat), .A2(G233gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n230), .B(KEYINPUT95), .ZN(new_n233));
  OR2_X1    g032(.A1(new_n233), .A2(new_n217), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n231), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT18), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n237), .A2(KEYINPUT96), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT96), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n239), .B1(new_n235), .B2(new_n236), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n233), .B(new_n217), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n232), .B(KEYINPUT13), .Z(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n231), .A2(new_n234), .A3(KEYINPUT18), .A4(new_n232), .ZN(new_n244));
  XNOR2_X1  g043(.A(G113gat), .B(G141gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(G197gat), .ZN(new_n246));
  XOR2_X1   g045(.A(KEYINPUT11), .B(G169gat), .Z(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(new_n248), .B(KEYINPUT12), .Z(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n243), .A2(new_n244), .A3(new_n250), .ZN(new_n251));
  NOR3_X1   g050(.A1(new_n238), .A2(new_n240), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n243), .A2(new_n244), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n250), .B1(new_n254), .B2(new_n237), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G78gat), .B(G106gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT31), .B(G50gat), .ZN(new_n258));
  XOR2_X1   g057(.A(new_n257), .B(new_n258), .Z(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(G228gat), .ZN(new_n261));
  INV_X1    g060(.A(G233gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G211gat), .B(G218gat), .ZN(new_n264));
  XOR2_X1   g063(.A(new_n264), .B(KEYINPUT74), .Z(new_n265));
  INV_X1    g064(.A(G197gat), .ZN(new_n266));
  INV_X1    g065(.A(G204gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G197gat), .A2(G204gat), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT22), .ZN(new_n270));
  NAND2_X1  g069(.A1(G211gat), .A2(G218gat), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n268), .A2(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n265), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n264), .B(KEYINPUT74), .ZN(new_n274));
  INV_X1    g073(.A(new_n272), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT29), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT3), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(G148gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(G141gat), .ZN(new_n281));
  INV_X1    g080(.A(G141gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(G148gat), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n281), .A2(new_n283), .B1(KEYINPUT78), .B2(KEYINPUT2), .ZN(new_n284));
  NAND2_X1  g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT78), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(G155gat), .ZN(new_n288));
  INV_X1    g087(.A(G162gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(KEYINPUT78), .A2(G155gat), .A3(G162gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n287), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n284), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT79), .B1(new_n282), .B2(G148gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT79), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n295), .A2(new_n280), .A3(G141gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n294), .A2(new_n296), .A3(new_n283), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n285), .B1(new_n290), .B2(KEYINPUT2), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT80), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n297), .A2(new_n298), .A3(KEYINPUT80), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n293), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OR2_X1    g102(.A1(new_n279), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT3), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n277), .B1(new_n306), .B2(new_n278), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n263), .B1(new_n304), .B2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n279), .A2(new_n303), .ZN(new_n310));
  INV_X1    g109(.A(new_n263), .ZN(new_n311));
  NOR3_X1   g110(.A1(new_n310), .A2(new_n311), .A3(new_n307), .ZN(new_n312));
  OAI21_X1  g111(.A(G22gat), .B1(new_n309), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n304), .A2(new_n263), .A3(new_n308), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n311), .B1(new_n310), .B2(new_n307), .ZN(new_n315));
  INV_X1    g114(.A(G22gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n260), .B1(new_n313), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n313), .A2(KEYINPUT85), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(new_n260), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n317), .A2(KEYINPUT86), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT86), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n314), .A2(new_n315), .A3(new_n323), .A4(new_n316), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT85), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n325), .B(G22gat), .C1(new_n309), .C2(new_n312), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n322), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n319), .B1(new_n321), .B2(new_n327), .ZN(new_n328));
  XOR2_X1   g127(.A(G1gat), .B(G29gat), .Z(new_n329));
  XNOR2_X1  g128(.A(G57gat), .B(G85gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n329), .B(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT1), .ZN(new_n335));
  INV_X1    g134(.A(G113gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n336), .A2(G120gat), .ZN(new_n337));
  INV_X1    g136(.A(G120gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n338), .A2(G113gat), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n335), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(KEYINPUT65), .A2(G134gat), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(KEYINPUT65), .A2(G134gat), .ZN(new_n343));
  INV_X1    g142(.A(G127gat), .ZN(new_n344));
  NOR3_X1   g143(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(G134gat), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT66), .B1(new_n346), .B2(G127gat), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT66), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n348), .A2(new_n344), .A3(G134gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n340), .B1(new_n345), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT67), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT67), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n340), .B(new_n353), .C1(new_n345), .C2(new_n350), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  XOR2_X1   g154(.A(G127gat), .B(G134gat), .Z(new_n356));
  OR2_X1    g155(.A1(new_n340), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n303), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT4), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n354), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT65), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(new_n346), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n363), .A2(G127gat), .A3(new_n341), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n364), .A2(new_n347), .A3(new_n349), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n353), .B1(new_n365), .B2(new_n340), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n357), .B1(new_n361), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT68), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT68), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n355), .A2(new_n369), .A3(new_n357), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n368), .A2(new_n303), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n360), .B1(new_n371), .B2(new_n359), .ZN(new_n372));
  INV_X1    g171(.A(new_n293), .ZN(new_n373));
  INV_X1    g172(.A(new_n302), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT80), .B1(new_n297), .B2(new_n298), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT3), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n377), .A2(new_n306), .A3(new_n367), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT5), .ZN(new_n379));
  NAND2_X1  g178(.A1(G225gat), .A2(G233gat), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n334), .B1(new_n372), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n380), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n367), .A2(new_n376), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n301), .A2(new_n302), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n355), .A2(new_n357), .B1(new_n385), .B2(new_n373), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n383), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT81), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(new_n388), .A3(KEYINPUT5), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n367), .A2(new_n376), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n380), .B1(new_n390), .B2(new_n358), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT81), .B1(new_n391), .B2(new_n379), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT82), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n368), .A2(KEYINPUT4), .A3(new_n370), .A4(new_n303), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n358), .A2(new_n359), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n395), .A2(new_n380), .A3(new_n378), .A4(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n393), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n394), .B1(new_n393), .B2(new_n397), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n382), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT6), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n388), .B1(new_n387), .B2(KEYINPUT5), .ZN(new_n404));
  NOR3_X1   g203(.A1(new_n391), .A2(KEYINPUT81), .A3(new_n379), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n397), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT82), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n398), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n372), .A2(new_n381), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n333), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT84), .B1(new_n403), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n409), .B1(new_n399), .B2(new_n400), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n334), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT6), .B1(new_n408), .B2(new_n382), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT84), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n410), .A2(KEYINPUT6), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n411), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(G226gat), .A2(G233gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(KEYINPUT75), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NOR2_X1   g220(.A1(G169gat), .A2(G176gat), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT23), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(G169gat), .ZN(new_n425));
  INV_X1    g224(.A(G176gat), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT24), .ZN(new_n428));
  NAND2_X1  g227(.A1(G183gat), .A2(G190gat), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n427), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(G183gat), .ZN(new_n432));
  INV_X1    g231(.A(G190gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n434), .A2(KEYINPUT24), .A3(new_n429), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n424), .A2(new_n431), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT25), .ZN(new_n437));
  OR2_X1    g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n436), .A2(new_n437), .ZN(new_n439));
  NOR3_X1   g238(.A1(new_n427), .A2(KEYINPUT26), .A3(new_n422), .ZN(new_n440));
  AOI211_X1 g239(.A(new_n430), .B(new_n440), .C1(KEYINPUT26), .C2(new_n422), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT27), .B1(new_n432), .B2(KEYINPUT64), .ZN(new_n442));
  OR2_X1    g241(.A1(new_n432), .A2(KEYINPUT27), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n433), .B(new_n442), .C1(new_n443), .C2(KEYINPUT64), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT28), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  XOR2_X1   g245(.A(KEYINPUT27), .B(G183gat), .Z(new_n447));
  NAND2_X1  g246(.A1(new_n433), .A2(KEYINPUT28), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AOI22_X1  g248(.A1(new_n438), .A2(new_n439), .B1(new_n441), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n421), .B1(new_n450), .B2(KEYINPUT29), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT76), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n452), .B1(new_n450), .B2(new_n419), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n436), .B(new_n437), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n441), .A2(new_n449), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n419), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(KEYINPUT76), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n451), .A2(new_n453), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n277), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n419), .B1(new_n450), .B2(KEYINPUT29), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n462), .B(new_n277), .C1(new_n450), .C2(new_n421), .ZN(new_n463));
  XNOR2_X1  g262(.A(G8gat), .B(G36gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(G64gat), .B(G92gat), .ZN(new_n465));
  XOR2_X1   g264(.A(new_n464), .B(new_n465), .Z(new_n466));
  NAND3_X1  g265(.A1(new_n461), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT77), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OR2_X1    g268(.A1(new_n469), .A2(KEYINPUT30), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n461), .A2(new_n463), .ZN(new_n471));
  INV_X1    g270(.A(new_n466), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n469), .A2(KEYINPUT30), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n328), .B1(new_n418), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G15gat), .B(G43gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n476), .B(KEYINPUT69), .ZN(new_n477));
  XNOR2_X1  g276(.A(G71gat), .B(G99gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n477), .B(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  OR2_X1    g279(.A1(new_n480), .A2(KEYINPUT70), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(KEYINPUT70), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n481), .A2(KEYINPUT33), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n368), .A2(new_n370), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n456), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n450), .A2(new_n368), .A3(new_n370), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(G227gat), .A2(G233gat), .ZN(new_n488));
  OAI211_X1 g287(.A(KEYINPUT32), .B(new_n483), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n488), .B1(new_n485), .B2(new_n486), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT32), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n479), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n490), .A2(KEYINPUT33), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n489), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT72), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n485), .A2(new_n488), .A3(new_n486), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT34), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT71), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n497), .B1(new_n488), .B2(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n496), .B(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n494), .A2(KEYINPUT72), .A3(new_n500), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n502), .A2(KEYINPUT36), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT36), .ZN(new_n505));
  OR3_X1    g304(.A1(new_n494), .A2(KEYINPUT73), .A3(new_n500), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n494), .A2(new_n500), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT73), .B1(new_n494), .B2(new_n500), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n504), .B1(new_n505), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT87), .B1(new_n475), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT87), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n502), .A2(KEYINPUT36), .A3(new_n503), .ZN(new_n513));
  INV_X1    g312(.A(new_n509), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n513), .B1(new_n514), .B2(KEYINPUT36), .ZN(new_n515));
  INV_X1    g314(.A(new_n474), .ZN(new_n516));
  AOI22_X1  g315(.A1(new_n407), .A2(new_n398), .B1(new_n372), .B2(new_n381), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n401), .B(new_n402), .C1(new_n517), .C2(new_n333), .ZN(new_n518));
  AOI22_X1  g317(.A1(new_n518), .A2(KEYINPUT84), .B1(KEYINPUT6), .B2(new_n410), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n516), .B1(new_n519), .B2(new_n416), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n512), .B(new_n515), .C1(new_n520), .C2(new_n328), .ZN(new_n521));
  INV_X1    g320(.A(new_n328), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n410), .B1(new_n470), .B2(new_n473), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n380), .B1(new_n372), .B2(new_n378), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n390), .A2(new_n358), .A3(new_n380), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT39), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT39), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n334), .B1(new_n524), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT40), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n522), .B1(new_n523), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n518), .A2(KEYINPUT88), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT88), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n413), .A2(new_n414), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n533), .A2(new_n417), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT37), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n459), .A2(new_n460), .ZN(new_n538));
  OR2_X1    g337(.A1(new_n538), .A2(KEYINPUT89), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n462), .B1(new_n450), .B2(new_n421), .ZN(new_n540));
  AOI22_X1  g339(.A1(new_n538), .A2(KEYINPUT89), .B1(new_n460), .B2(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n537), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT38), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n543), .B(new_n472), .C1(new_n471), .C2(KEYINPUT37), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n472), .B1(new_n471), .B2(KEYINPUT37), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n545), .B1(KEYINPUT37), .B2(new_n471), .ZN(new_n546));
  OAI221_X1 g345(.A(new_n467), .B1(new_n542), .B2(new_n544), .C1(new_n546), .C2(new_n543), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n532), .B1(new_n536), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n511), .A2(new_n521), .A3(new_n548), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n328), .A2(new_n502), .A3(new_n503), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n418), .A2(new_n474), .A3(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT90), .B(KEYINPUT35), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n474), .A2(new_n328), .A3(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n553), .A2(new_n509), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n551), .A2(KEYINPUT35), .B1(new_n554), .B2(new_n536), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n256), .B1(new_n549), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n418), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT99), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT7), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT7), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT99), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n560), .A2(new_n562), .A3(G85gat), .A4(G92gat), .ZN(new_n563));
  INV_X1    g362(.A(G85gat), .ZN(new_n564));
  INV_X1    g363(.A(G92gat), .ZN(new_n565));
  OAI211_X1 g364(.A(KEYINPUT99), .B(new_n561), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G99gat), .A2(G106gat), .ZN(new_n567));
  AOI22_X1  g366(.A1(KEYINPUT8), .A2(new_n567), .B1(new_n564), .B2(new_n565), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n563), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  OR2_X1    g368(.A1(G99gat), .A2(G106gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(new_n567), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n567), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n563), .A2(new_n572), .A3(new_n566), .A4(new_n568), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n571), .A2(KEYINPUT100), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n571), .A2(new_n573), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT100), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n219), .A2(new_n574), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n217), .B1(new_n574), .B2(new_n577), .ZN(new_n579));
  AND2_X1   g378(.A1(G232gat), .A2(G233gat), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n579), .B1(KEYINPUT41), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT101), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT101), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n578), .A2(new_n584), .A3(new_n581), .ZN(new_n585));
  XOR2_X1   g384(.A(G134gat), .B(G162gat), .Z(new_n586));
  AND3_X1   g385(.A1(new_n583), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n586), .B1(new_n583), .B2(new_n585), .ZN(new_n588));
  XOR2_X1   g387(.A(G190gat), .B(G218gat), .Z(new_n589));
  NOR2_X1   g388(.A1(new_n580), .A2(KEYINPUT41), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  OR3_X1    g390(.A1(new_n587), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n591), .B1(new_n587), .B2(new_n588), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G57gat), .B(G64gat), .Z(new_n596));
  INV_X1    g395(.A(KEYINPUT9), .ZN(new_n597));
  INV_X1    g396(.A(G71gat), .ZN(new_n598));
  INV_X1    g397(.A(G78gat), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G71gat), .B(G78gat), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n596), .A2(new_n602), .A3(new_n600), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT21), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G231gat), .A2(G233gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(G127gat), .B(G155gat), .Z(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G183gat), .B(G211gat), .Z(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n233), .B1(new_n607), .B2(new_n606), .ZN(new_n617));
  XNOR2_X1  g416(.A(KEYINPUT98), .B(KEYINPUT20), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n617), .B(new_n618), .Z(new_n619));
  AND2_X1   g418(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n616), .A2(new_n619), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G230gat), .A2(G233gat), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n606), .B1(KEYINPUT102), .B2(new_n573), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(new_n575), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n573), .B(new_n571), .C1(new_n606), .C2(KEYINPUT102), .ZN(new_n626));
  AOI21_X1  g425(.A(KEYINPUT10), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT10), .ZN(new_n628));
  AOI211_X1 g427(.A(new_n628), .B(new_n606), .C1(new_n577), .C2(new_n574), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n623), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n625), .A2(new_n626), .ZN(new_n631));
  INV_X1    g430(.A(new_n623), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(G120gat), .B(G148gat), .Z(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT103), .ZN(new_n636));
  XNOR2_X1  g435(.A(G176gat), .B(G204gat), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n636), .B(new_n637), .Z(new_n638));
  OR2_X1    g437(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n634), .A2(new_n638), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n595), .A2(new_n622), .A3(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n557), .A2(new_n558), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(G1gat), .ZN(G1324gat));
  INV_X1    g445(.A(KEYINPUT42), .ZN(new_n647));
  AND3_X1   g446(.A1(new_n557), .A2(new_n516), .A3(new_n644), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n648), .A2(new_n227), .ZN(new_n649));
  XOR2_X1   g448(.A(KEYINPUT16), .B(G8gat), .Z(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n647), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(KEYINPUT42), .B1(new_n648), .B2(new_n650), .ZN(new_n653));
  OR3_X1    g452(.A1(new_n652), .A2(KEYINPUT104), .A3(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(KEYINPUT104), .B1(new_n652), .B2(new_n653), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(G1325gat));
  NAND2_X1  g455(.A1(new_n557), .A2(new_n644), .ZN(new_n657));
  OAI21_X1  g456(.A(G15gat), .B1(new_n657), .B2(new_n515), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n509), .A2(G15gat), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n658), .B1(new_n657), .B2(new_n659), .ZN(G1326gat));
  NOR2_X1   g459(.A1(new_n657), .A2(new_n328), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT43), .B(G22gat), .Z(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(G1327gat));
  NOR3_X1   g462(.A1(new_n595), .A2(new_n622), .A3(new_n641), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n557), .A2(new_n664), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n665), .A2(G29gat), .A3(new_n418), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT45), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT35), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n669), .B1(new_n520), .B2(new_n550), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n554), .A2(new_n536), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT106), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n551), .A2(KEYINPUT35), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT106), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n554), .A2(new_n536), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  OAI211_X1 g475(.A(new_n548), .B(new_n515), .C1(new_n520), .C2(new_n328), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n672), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n594), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n549), .A2(new_n556), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n595), .A2(new_n680), .ZN(new_n682));
  AOI22_X1  g481(.A1(new_n679), .A2(new_n680), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n641), .B(KEYINPUT105), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n622), .A2(new_n256), .A3(new_n684), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n683), .A2(KEYINPUT107), .A3(new_n558), .A4(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT107), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n681), .A2(new_n682), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n418), .A2(new_n474), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n510), .B1(new_n689), .B2(new_n522), .ZN(new_n690));
  AOI22_X1  g489(.A1(new_n555), .A2(new_n674), .B1(new_n690), .B2(new_n548), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n595), .B1(new_n691), .B2(new_n672), .ZN(new_n692));
  OAI211_X1 g491(.A(new_n688), .B(new_n685), .C1(new_n692), .C2(KEYINPUT44), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n687), .B1(new_n693), .B2(new_n418), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n686), .A2(new_n694), .A3(G29gat), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n668), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT108), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT108), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n668), .A2(new_n695), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(new_n699), .ZN(G1328gat));
  NOR3_X1   g499(.A1(new_n665), .A2(G36gat), .A3(new_n474), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT46), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT109), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n693), .A2(new_n703), .A3(new_n474), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n703), .B1(new_n693), .B2(new_n474), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(G36gat), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n702), .B1(new_n704), .B2(new_n706), .ZN(G1329gat));
  OR3_X1    g506(.A1(new_n665), .A2(G43gat), .A3(new_n509), .ZN(new_n708));
  AOI21_X1  g507(.A(KEYINPUT47), .B1(new_n708), .B2(KEYINPUT110), .ZN(new_n709));
  OAI21_X1  g508(.A(G43gat), .B1(new_n693), .B2(new_n515), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n708), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n709), .B(new_n711), .ZN(G1330gat));
  OAI21_X1  g511(.A(G50gat), .B1(new_n693), .B2(new_n328), .ZN(new_n713));
  OR3_X1    g512(.A1(new_n665), .A2(G50gat), .A3(new_n328), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n715), .B(KEYINPUT48), .Z(G1331gat));
  NAND2_X1  g515(.A1(new_n676), .A2(new_n677), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n555), .A2(new_n674), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n595), .A2(new_n622), .A3(new_n256), .A4(new_n684), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n558), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(G57gat), .ZN(G1332gat));
  INV_X1    g522(.A(new_n721), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(new_n474), .ZN(new_n725));
  NOR2_X1   g524(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n726));
  AND2_X1   g525(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n728), .B1(new_n725), .B2(new_n726), .ZN(G1333gat));
  OAI21_X1  g528(.A(KEYINPUT111), .B1(new_n724), .B2(new_n509), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT111), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n721), .A2(new_n731), .A3(new_n514), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n730), .A2(new_n598), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n721), .A2(G71gat), .A3(new_n510), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n522), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(G78gat), .ZN(G1335gat));
  OR2_X1    g537(.A1(new_n620), .A2(new_n621), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n256), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT112), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n741), .A2(new_n641), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n688), .B(new_n742), .C1(new_n692), .C2(KEYINPUT44), .ZN(new_n743));
  OAI21_X1  g542(.A(G85gat), .B1(new_n743), .B2(new_n418), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n594), .B(new_n741), .C1(new_n717), .C2(new_n718), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT51), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n678), .A2(KEYINPUT51), .A3(new_n594), .A4(new_n741), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n558), .A2(new_n564), .A3(new_n641), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n744), .B1(new_n750), .B2(new_n751), .ZN(G1336gat));
  INV_X1    g551(.A(KEYINPUT113), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n747), .A2(new_n753), .A3(new_n748), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n745), .A2(KEYINPUT113), .A3(new_n746), .ZN(new_n755));
  INV_X1    g554(.A(new_n684), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n756), .A2(new_n474), .A3(G92gat), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n754), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(G92gat), .B1(new_n743), .B2(new_n474), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT52), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n749), .A2(new_n757), .ZN(new_n763));
  XOR2_X1   g562(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n764));
  NAND3_X1  g563(.A1(new_n759), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n761), .A2(new_n762), .A3(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n767), .B1(new_n758), .B2(new_n759), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n759), .A2(new_n763), .A3(new_n764), .ZN(new_n769));
  OAI21_X1  g568(.A(KEYINPUT115), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n766), .A2(new_n770), .ZN(G1337gat));
  NOR2_X1   g570(.A1(new_n642), .A2(G99gat), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n749), .A2(new_n514), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(G99gat), .B1(new_n743), .B2(new_n515), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT116), .ZN(G1338gat));
  NOR3_X1   g575(.A1(new_n756), .A2(G106gat), .A3(new_n328), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n754), .A2(new_n755), .A3(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(G106gat), .B1(new_n743), .B2(new_n328), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT53), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT53), .B1(new_n749), .B2(new_n777), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n779), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(G1339gat));
  INV_X1    g583(.A(new_n256), .ZN(new_n785));
  OR3_X1    g584(.A1(new_n627), .A2(new_n629), .A3(new_n623), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n786), .A2(KEYINPUT54), .A3(new_n630), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n788), .B(new_n623), .C1(new_n627), .C2(new_n629), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n789), .A2(new_n638), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n787), .A2(KEYINPUT55), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n639), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(KEYINPUT117), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n787), .A2(new_n790), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT117), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n791), .A2(new_n797), .A3(new_n639), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n793), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT118), .ZN(new_n800));
  AOI22_X1  g599(.A1(new_n792), .A2(KEYINPUT117), .B1(new_n795), .B2(new_n794), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(new_n802), .A3(new_n798), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n785), .A2(new_n800), .A3(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n252), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n241), .A2(new_n242), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n232), .B1(new_n231), .B2(new_n234), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n248), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n805), .A2(new_n641), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n594), .B1(new_n804), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n805), .A2(new_n808), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n811), .A2(new_n594), .A3(new_n800), .A4(new_n803), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n739), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n643), .A2(new_n785), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n522), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n418), .A2(new_n516), .A3(new_n509), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n819), .A2(new_n336), .A3(new_n256), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n814), .A2(new_n816), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n822), .A2(new_n418), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n823), .A2(new_n550), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n824), .A2(new_n785), .A3(new_n474), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n820), .B1(new_n825), .B2(new_n336), .ZN(G1340gat));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n474), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n338), .B1(new_n827), .B2(new_n642), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n817), .A2(G120gat), .A3(new_n684), .A4(new_n818), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(KEYINPUT119), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n828), .A2(new_n832), .A3(new_n829), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(G1341gat));
  OAI21_X1  g633(.A(G127gat), .B1(new_n819), .B2(new_n739), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n622), .A2(new_n344), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n835), .B1(new_n827), .B2(new_n836), .ZN(G1342gat));
  NAND2_X1  g636(.A1(new_n594), .A2(new_n474), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT120), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n824), .A2(new_n363), .A3(new_n341), .A4(new_n840), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n841), .A2(KEYINPUT56), .ZN(new_n842));
  OAI21_X1  g641(.A(G134gat), .B1(new_n819), .B2(new_n595), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(KEYINPUT56), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(G1343gat));
  NAND2_X1  g644(.A1(new_n821), .A2(new_n522), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(KEYINPUT122), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n522), .A2(KEYINPUT57), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT124), .ZN(new_n851));
  INV_X1    g650(.A(new_n792), .ZN(new_n852));
  XOR2_X1   g651(.A(KEYINPUT123), .B(KEYINPUT55), .Z(new_n853));
  NAND2_X1  g652(.A1(new_n794), .A2(new_n853), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n852), .B(new_n854), .C1(new_n252), .C2(new_n255), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n809), .A2(new_n851), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n851), .B1(new_n809), .B2(new_n855), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n595), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n622), .B1(new_n858), .B2(new_n812), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n850), .B1(new_n859), .B2(new_n815), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT125), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT122), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n328), .B1(new_n814), .B2(new_n816), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n863), .B1(new_n864), .B2(KEYINPUT57), .ZN(new_n865));
  OAI211_X1 g664(.A(KEYINPUT125), .B(new_n850), .C1(new_n859), .C2(new_n815), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n848), .A2(new_n862), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n510), .A2(new_n418), .A3(new_n516), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(KEYINPUT121), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n867), .A2(new_n785), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(G141gat), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n510), .A2(new_n328), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n256), .A2(G141gat), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n823), .A2(new_n474), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT126), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT58), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n871), .A2(new_n874), .A3(new_n878), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(G1344gat));
  NOR2_X1   g681(.A1(new_n280), .A2(KEYINPUT59), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n869), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n883), .B1(new_n884), .B2(new_n642), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n811), .A2(new_n594), .A3(new_n798), .A4(new_n801), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n622), .B1(new_n858), .B2(new_n886), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n847), .B(new_n522), .C1(new_n887), .C2(new_n815), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n888), .B1(new_n847), .B2(new_n864), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n869), .A2(new_n641), .ZN(new_n890));
  OAI21_X1  g689(.A(G148gat), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT59), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n885), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n823), .A2(new_n872), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n894), .A2(new_n516), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n280), .A3(new_n641), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n893), .A2(new_n896), .ZN(G1345gat));
  OAI21_X1  g696(.A(G155gat), .B1(new_n884), .B2(new_n739), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n895), .A2(new_n288), .A3(new_n622), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(G1346gat));
  OAI21_X1  g699(.A(G162gat), .B1(new_n884), .B2(new_n595), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n840), .A2(new_n289), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n894), .B2(new_n902), .ZN(G1347gat));
  NOR2_X1   g702(.A1(new_n822), .A2(new_n558), .ZN(new_n904));
  AND3_X1   g703(.A1(new_n904), .A2(new_n516), .A3(new_n550), .ZN(new_n905));
  AOI21_X1  g704(.A(G169gat), .B1(new_n905), .B2(new_n785), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n558), .A2(new_n474), .A3(new_n509), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n817), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n256), .A2(new_n425), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(G1348gat));
  NAND3_X1  g709(.A1(new_n905), .A2(new_n426), .A3(new_n641), .ZN(new_n911));
  INV_X1    g710(.A(new_n908), .ZN(new_n912));
  OAI21_X1  g711(.A(G176gat), .B1(new_n912), .B2(new_n756), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(G1349gat));
  AOI21_X1  g713(.A(new_n432), .B1(new_n908), .B2(new_n622), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n739), .A2(new_n447), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(new_n905), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(KEYINPUT127), .A2(KEYINPUT60), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n917), .B(new_n918), .ZN(G1350gat));
  AOI21_X1  g718(.A(new_n433), .B1(new_n908), .B2(new_n594), .ZN(new_n920));
  XOR2_X1   g719(.A(new_n920), .B(KEYINPUT61), .Z(new_n921));
  NAND3_X1  g720(.A1(new_n905), .A2(new_n433), .A3(new_n594), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(G1351gat));
  NAND3_X1  g722(.A1(new_n515), .A2(new_n418), .A3(new_n516), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n889), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n785), .A2(G197gat), .ZN(new_n926));
  AND4_X1   g725(.A1(new_n418), .A2(new_n821), .A3(new_n516), .A4(new_n872), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n927), .A2(new_n785), .ZN(new_n928));
  OAI22_X1  g727(.A1(new_n925), .A2(new_n926), .B1(G197gat), .B2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(G1352gat));
  NAND3_X1  g729(.A1(new_n927), .A2(new_n267), .A3(new_n641), .ZN(new_n931));
  XOR2_X1   g730(.A(new_n931), .B(KEYINPUT62), .Z(new_n932));
  OAI21_X1  g731(.A(G204gat), .B1(new_n925), .B2(new_n756), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1353gat));
  INV_X1    g733(.A(G211gat), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n927), .A2(new_n935), .A3(new_n622), .ZN(new_n936));
  OR3_X1    g735(.A1(new_n889), .A2(new_n739), .A3(new_n924), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n937), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(KEYINPUT63), .B1(new_n937), .B2(G211gat), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n936), .B1(new_n939), .B2(new_n940), .ZN(G1354gat));
  OAI21_X1  g740(.A(G218gat), .B1(new_n925), .B2(new_n595), .ZN(new_n942));
  INV_X1    g741(.A(G218gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n927), .A2(new_n943), .A3(new_n594), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n942), .A2(new_n944), .ZN(G1355gat));
endmodule


