//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 1 0 1 0 1 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1222, new_n1223, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n202), .B(KEYINPUT64), .ZN(G355));
  NAND2_X1  g0003(.A1(G1), .A2(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G13), .ZN(new_n205));
  OAI211_X1 g0005(.A(new_n205), .B(G250), .C1(G257), .C2(G264), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT0), .Z(new_n207));
  AOI22_X1  g0007(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n208));
  INV_X1    g0008(.A(G68), .ZN(new_n209));
  INV_X1    g0009(.A(G238), .ZN(new_n210));
  INV_X1    g0010(.A(G107), .ZN(new_n211));
  INV_X1    g0011(.A(G264), .ZN(new_n212));
  OAI221_X1 g0012(.A(new_n208), .B1(new_n209), .B2(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n213), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G50), .ZN(new_n215));
  INV_X1    g0015(.A(G226), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G58), .ZN(new_n220));
  INV_X1    g0020(.A(G232), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n204), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(KEYINPUT65), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g0028(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n225), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(G50), .B1(G58), .B2(G68), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n207), .B(new_n224), .C1(new_n230), .C2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n212), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  NAND2_X1  g0041(.A1(new_n211), .A2(G97), .ZN(new_n242));
  INV_X1    g0042(.A(G97), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G107), .ZN(new_n244));
  AND2_X1   g0044(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n252), .B1(G41), .B2(G45), .ZN(new_n253));
  INV_X1    g0053(.A(G274), .ZN(new_n254));
  OR2_X1    g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  OR2_X1    g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n259), .A2(G226), .A3(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n259), .A2(G232), .A3(G1698), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n261), .B(new_n262), .C1(new_n263), .C2(new_n243), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  AND3_X1   g0065(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n266));
  AOI21_X1  g0066(.A(KEYINPUT65), .B1(G1), .B2(G13), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n256), .B1(new_n264), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT13), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n265), .A2(G1), .A3(G13), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n253), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G238), .ZN(new_n275));
  AND3_X1   g0075(.A1(new_n270), .A2(new_n271), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n271), .B1(new_n270), .B2(new_n275), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G190), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n270), .A2(new_n275), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT13), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n270), .A2(new_n271), .A3(new_n275), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G200), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n252), .A2(G13), .A3(G20), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT68), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n252), .A2(KEYINPUT68), .A3(G13), .A4(G20), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n209), .ZN(new_n291));
  XNOR2_X1  g0091(.A(new_n291), .B(KEYINPUT12), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n228), .A2(new_n229), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n252), .A2(G20), .ZN(new_n296));
  AND3_X1   g0096(.A1(new_n295), .A2(new_n289), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G68), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n209), .A2(G20), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n225), .A2(G33), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n225), .A2(new_n263), .ZN(new_n302));
  OAI221_X1 g0102(.A(new_n300), .B1(new_n301), .B2(new_n217), .C1(new_n215), .C2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n294), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n304), .A2(KEYINPUT71), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(KEYINPUT71), .ZN(new_n306));
  AND3_X1   g0106(.A1(new_n305), .A2(KEYINPUT11), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(KEYINPUT11), .B1(new_n305), .B2(new_n306), .ZN(new_n308));
  NOR3_X1   g0108(.A1(new_n299), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  AND3_X1   g0109(.A1(new_n279), .A2(new_n284), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n309), .ZN(new_n311));
  OAI21_X1  g0111(.A(G169), .B1(new_n276), .B2(new_n277), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT14), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT14), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n283), .A2(new_n314), .A3(G169), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n278), .A2(G179), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n313), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n310), .B1(new_n311), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n257), .A2(new_n225), .A3(new_n258), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT7), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AND2_X1   g0121(.A1(KEYINPUT3), .A2(G33), .ZN(new_n322));
  NOR2_X1   g0122(.A1(KEYINPUT3), .A2(G33), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(KEYINPUT7), .B1(new_n324), .B2(new_n225), .ZN(new_n325));
  OAI21_X1  g0125(.A(G68), .B1(new_n321), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT72), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT16), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n220), .A2(new_n209), .ZN(new_n329));
  NOR2_X1   g0129(.A1(G58), .A2(G68), .ZN(new_n330));
  OAI21_X1  g0130(.A(G20), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n302), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G159), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n326), .A2(new_n327), .A3(new_n328), .A4(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n326), .A2(new_n328), .A3(new_n335), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n319), .A2(new_n320), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n324), .A2(KEYINPUT7), .A3(new_n225), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n209), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(KEYINPUT16), .B1(new_n340), .B2(new_n334), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  NOR3_X1   g0142(.A1(new_n326), .A2(KEYINPUT72), .A3(new_n334), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n294), .B(new_n336), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n216), .A2(G1698), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n259), .B(new_n345), .C1(G223), .C2(G1698), .ZN(new_n346));
  NAND2_X1  g0146(.A1(G33), .A2(G87), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n268), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n255), .B1(new_n273), .B2(new_n221), .ZN(new_n349));
  OR2_X1    g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G190), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT8), .B(G58), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n289), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(new_n297), .B2(new_n353), .ZN(new_n355));
  AND3_X1   g0155(.A1(new_n344), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT17), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(KEYINPUT74), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n350), .A2(G200), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n357), .A2(KEYINPUT74), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n356), .A2(new_n359), .A3(new_n360), .A4(new_n361), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n344), .A2(new_n360), .A3(new_n352), .A4(new_n355), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n363), .A2(KEYINPUT74), .A3(new_n357), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(G169), .B1(new_n348), .B2(new_n349), .ZN(new_n366));
  INV_X1    g0166(.A(G179), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n366), .B1(new_n350), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT73), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT73), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n370), .B(new_n366), .C1(new_n350), .C2(new_n367), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n344), .A2(new_n355), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n372), .A2(new_n373), .A3(KEYINPUT18), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT18), .B1(new_n372), .B2(new_n373), .ZN(new_n375));
  OR2_X1    g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT67), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n324), .B2(new_n260), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n259), .A2(KEYINPUT67), .A3(G1698), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(new_n379), .A3(G238), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n259), .A2(G232), .A3(new_n260), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n380), .B(new_n381), .C1(new_n211), .C2(new_n259), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n269), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n256), .B1(new_n274), .B2(G244), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n367), .ZN(new_n387));
  OAI22_X1  g0187(.A1(new_n353), .A2(new_n302), .B1(new_n225), .B2(new_n217), .ZN(new_n388));
  XNOR2_X1  g0188(.A(KEYINPUT15), .B(G87), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n389), .A2(new_n301), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n294), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n297), .A2(G77), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n391), .B(new_n392), .C1(G77), .C2(new_n289), .ZN(new_n393));
  INV_X1    g0193(.A(G169), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n385), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n387), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n318), .A2(new_n365), .A3(new_n376), .A4(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n255), .B1(new_n273), .B2(new_n216), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT66), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n255), .B(KEYINPUT66), .C1(new_n216), .C2(new_n273), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n378), .A2(new_n379), .A3(G223), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n259), .A2(G222), .A3(new_n260), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n403), .B(new_n404), .C1(new_n217), .C2(new_n259), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n402), .B1(new_n405), .B2(new_n269), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n407), .A2(G179), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n290), .A2(new_n215), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n295), .A2(new_n289), .A3(G50), .A4(new_n296), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n353), .A2(new_n301), .ZN(new_n411));
  NOR3_X1   g0211(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n412));
  INV_X1    g0212(.A(G150), .ZN(new_n413));
  OAI22_X1  g0213(.A1(new_n412), .A2(new_n225), .B1(new_n302), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n294), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n409), .A2(new_n410), .A3(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n406), .A2(G169), .ZN(new_n417));
  NOR3_X1   g0217(.A1(new_n408), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT9), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n409), .A2(new_n410), .A3(new_n415), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT9), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n406), .A2(G190), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT70), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n407), .A2(G200), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n423), .B2(new_n424), .ZN(new_n427));
  OAI21_X1  g0227(.A(KEYINPUT10), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n420), .A2(KEYINPUT69), .A3(new_n422), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT10), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(KEYINPUT69), .B1(new_n420), .B2(new_n422), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n433), .B(new_n426), .C1(new_n351), .C2(new_n407), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n418), .B1(new_n428), .B2(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n385), .A2(new_n351), .ZN(new_n436));
  OR2_X1    g0236(.A1(new_n436), .A2(new_n393), .ZN(new_n437));
  INV_X1    g0237(.A(G200), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n386), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n435), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(KEYINPUT75), .B1(new_n397), .B2(new_n442), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n362), .B(new_n364), .C1(new_n374), .C2(new_n375), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n317), .A2(new_n311), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n279), .A2(new_n284), .A3(new_n309), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  AOI211_X1 g0248(.A(new_n418), .B(new_n440), .C1(new_n428), .C2(new_n434), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT75), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n448), .A2(new_n449), .A3(new_n450), .A4(new_n396), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n443), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT22), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT84), .ZN(new_n454));
  AOI21_X1  g0254(.A(G20), .B1(new_n257), .B2(new_n258), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n454), .B1(new_n455), .B2(G87), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n225), .B(G87), .C1(new_n322), .C2(new_n323), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(KEYINPUT84), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n453), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n225), .A2(KEYINPUT23), .A3(G107), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G33), .A2(G116), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(G20), .ZN(new_n462));
  OAI21_X1  g0262(.A(KEYINPUT23), .B1(new_n225), .B2(G107), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT85), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT85), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n465), .B(KEYINPUT23), .C1(new_n225), .C2(G107), .ZN(new_n466));
  AOI211_X1 g0266(.A(new_n460), .B(new_n462), .C1(new_n464), .C2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n455), .A2(new_n454), .A3(G87), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n457), .A2(KEYINPUT84), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n468), .A2(new_n469), .A3(KEYINPUT22), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n459), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT86), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT86), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n459), .A2(new_n473), .A3(new_n467), .A4(new_n470), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(KEYINPUT24), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT24), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n471), .A2(KEYINPUT86), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n475), .A2(new_n294), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(G41), .ZN(new_n479));
  AND2_X1   g0279(.A1(KEYINPUT78), .A2(KEYINPUT5), .ZN(new_n480));
  NOR2_X1   g0280(.A1(KEYINPUT78), .A2(KEYINPUT5), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT79), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT79), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n484), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT5), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G41), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n487), .A2(new_n252), .A3(G45), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n483), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n489), .A2(G264), .A3(new_n272), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT87), .ZN(new_n491));
  OAI22_X1  g0291(.A1(new_n322), .A2(new_n323), .B1(G250), .B2(G1698), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n260), .A2(G257), .ZN(new_n493));
  INV_X1    g0293(.A(G294), .ZN(new_n494));
  OAI22_X1  g0294(.A1(new_n492), .A2(new_n493), .B1(new_n263), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n269), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n252), .A2(G45), .A3(G274), .ZN(new_n497));
  INV_X1    g0297(.A(new_n226), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n497), .B1(new_n498), .B2(new_n265), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n483), .A2(new_n485), .A3(new_n487), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT87), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n489), .A2(new_n503), .A3(G264), .A4(new_n272), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n491), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n438), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n502), .A2(new_n351), .A3(new_n490), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n252), .A2(G33), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n295), .A2(new_n289), .A3(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n290), .A2(KEYINPUT25), .A3(new_n211), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT25), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n289), .B2(G107), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n511), .A2(G107), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n478), .A2(new_n508), .A3(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n490), .ZN(new_n517));
  OAI21_X1  g0317(.A(G169), .B1(new_n517), .B2(new_n501), .ZN(new_n518));
  INV_X1    g0318(.A(new_n500), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(new_n367), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n491), .A2(new_n520), .A3(new_n496), .A4(new_n504), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n478), .A2(new_n515), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n516), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n510), .A2(new_n243), .ZN(new_n524));
  OAI21_X1  g0324(.A(G107), .B1(new_n321), .B2(new_n325), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n332), .A2(G77), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT6), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT76), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT76), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(KEYINPUT6), .ZN(new_n530));
  AND4_X1   g0330(.A1(new_n242), .A2(new_n244), .A3(new_n528), .A4(new_n530), .ZN(new_n531));
  XNOR2_X1  g0331(.A(KEYINPUT76), .B(KEYINPUT6), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n532), .A2(new_n242), .ZN(new_n533));
  OAI21_X1  g0333(.A(G20), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n525), .A2(new_n526), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n524), .B1(new_n535), .B2(new_n294), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n289), .A2(G97), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(G250), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n540), .B1(new_n257), .B2(new_n258), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT77), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n542), .A2(KEYINPUT4), .ZN(new_n543));
  OAI21_X1  g0343(.A(G1698), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G33), .A2(G283), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(G244), .B1(new_n322), .B2(new_n323), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n546), .B1(new_n547), .B2(new_n543), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n218), .B1(new_n257), .B2(new_n258), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n542), .B1(new_n549), .B2(new_n260), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT4), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n544), .B(new_n548), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n519), .B1(new_n552), .B2(new_n269), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n489), .A2(G257), .A3(new_n272), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n394), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n544), .A2(new_n548), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n259), .A2(G244), .A3(new_n260), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n551), .B1(new_n557), .B2(KEYINPUT77), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n269), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  AND4_X1   g0359(.A1(G179), .A2(new_n559), .A3(new_n500), .A4(new_n554), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n539), .B1(new_n555), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n301), .A2(new_n243), .ZN(new_n562));
  XNOR2_X1  g0362(.A(KEYINPUT81), .B(KEYINPUT19), .ZN(new_n563));
  OR2_X1    g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n455), .A2(G68), .ZN(new_n565));
  XNOR2_X1  g0365(.A(KEYINPUT82), .B(G87), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n566), .A2(new_n243), .A3(new_n211), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n263), .A2(new_n243), .ZN(new_n568));
  AOI21_X1  g0368(.A(G20), .B1(new_n563), .B2(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n564), .B(new_n565), .C1(new_n567), .C2(new_n569), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n570), .A2(new_n294), .B1(new_n290), .B2(new_n389), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(new_n389), .B2(new_n510), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n210), .A2(new_n260), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n218), .A2(G1698), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n573), .B(new_n574), .C1(new_n322), .C2(new_n323), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n461), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n269), .ZN(new_n577));
  INV_X1    g0377(.A(new_n499), .ZN(new_n578));
  INV_X1    g0378(.A(G45), .ZN(new_n579));
  OAI21_X1  g0379(.A(G250), .B1(new_n579), .B2(G1), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n580), .B1(new_n498), .B2(new_n265), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n577), .A2(new_n578), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(G169), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT80), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n499), .B1(new_n576), .B2(new_n269), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n586), .A2(G179), .A3(new_n582), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n584), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n585), .B1(new_n584), .B2(new_n587), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n572), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AOI211_X1 g0390(.A(new_n537), .B(new_n524), .C1(new_n535), .C2(new_n294), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n559), .A2(new_n500), .A3(new_n554), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G200), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n553), .A2(G190), .A3(new_n554), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n511), .A2(G87), .ZN(new_n596));
  AND2_X1   g0396(.A1(new_n571), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n583), .A2(G200), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n268), .B1(new_n461), .B2(new_n575), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n599), .A2(new_n499), .A3(new_n581), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(G190), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n597), .A2(new_n598), .A3(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n561), .A2(new_n590), .A3(new_n595), .A4(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT83), .ZN(new_n604));
  INV_X1    g0404(.A(G116), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(G20), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n545), .B(new_n225), .C1(G33), .C2(new_n243), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n294), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT20), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n294), .A2(KEYINPUT20), .A3(new_n606), .A4(new_n607), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n290), .A2(new_n605), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n295), .A2(new_n289), .A3(G116), .A4(new_n509), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G179), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n489), .A2(G270), .A3(new_n272), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n260), .A2(G257), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n259), .B(new_n618), .C1(new_n212), .C2(new_n260), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n619), .B(new_n269), .C1(G303), .C2(new_n259), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n617), .A2(new_n500), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n604), .B1(new_n616), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n621), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n623), .A2(KEYINPUT83), .A3(G179), .A4(new_n615), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n621), .A2(new_n615), .A3(G169), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(KEYINPUT21), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT21), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n621), .A2(new_n615), .A3(new_n628), .A4(G169), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n621), .A2(G200), .ZN(new_n631));
  INV_X1    g0431(.A(new_n615), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n631), .B(new_n632), .C1(new_n351), .C2(new_n621), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n625), .A2(new_n630), .A3(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n603), .A2(new_n634), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n452), .A2(new_n523), .A3(new_n635), .ZN(G372));
  NAND2_X1  g0436(.A1(new_n584), .A2(new_n587), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n572), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n561), .A2(new_n595), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n625), .A2(new_n630), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n640), .B1(new_n522), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n478), .A2(new_n508), .A3(new_n515), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n598), .A2(KEYINPUT88), .ZN(new_n644));
  OR3_X1    g0444(.A1(new_n600), .A2(KEYINPUT88), .A3(new_n438), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n597), .A2(new_n601), .A3(new_n644), .A4(new_n645), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n646), .A2(KEYINPUT89), .A3(new_n638), .ZN(new_n647));
  AOI21_X1  g0447(.A(KEYINPUT89), .B1(new_n646), .B2(new_n638), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n643), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n638), .B1(new_n642), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n590), .A2(new_n602), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT26), .B1(new_n651), .B2(new_n561), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT90), .B1(new_n555), .B2(new_n560), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n592), .A2(G169), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT90), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n654), .B(new_n655), .C1(new_n367), .C2(new_n592), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n591), .B1(new_n653), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n647), .B2(new_n648), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n652), .B1(new_n658), .B2(KEYINPUT26), .ZN(new_n659));
  OR2_X1    g0459(.A1(new_n650), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n452), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n368), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n662), .B1(new_n344), .B2(new_n355), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT18), .ZN(new_n664));
  INV_X1    g0464(.A(new_n365), .ZN(new_n665));
  INV_X1    g0465(.A(new_n396), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n446), .A2(new_n666), .B1(new_n317), .B2(new_n311), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n664), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n428), .A2(new_n434), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n418), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n661), .A2(new_n670), .ZN(G369));
  NAND2_X1  g0471(.A1(new_n478), .A2(new_n515), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n252), .A2(new_n225), .A3(G13), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AOI211_X1 g0478(.A(new_n522), .B(new_n516), .C1(new_n672), .C2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n521), .A2(new_n518), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n672), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n678), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n625), .A2(new_n630), .ZN(new_n685));
  OAI211_X1 g0485(.A(new_n685), .B(new_n633), .C1(new_n632), .C2(new_n682), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n641), .A2(new_n615), .A3(new_n678), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(G330), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n684), .A2(new_n689), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n643), .B(new_n682), .C1(new_n522), .C2(new_n641), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(G399));
  INV_X1    g0492(.A(new_n205), .ZN(new_n693));
  OR3_X1    g0493(.A1(new_n693), .A2(KEYINPUT91), .A3(G41), .ZN(new_n694));
  OAI21_X1  g0494(.A(KEYINPUT91), .B1(new_n693), .B2(G41), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n696), .A2(G1), .A3(new_n605), .A4(new_n567), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n231), .B2(new_n696), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT92), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT28), .ZN(new_n700));
  INV_X1    g0500(.A(new_n648), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n646), .A2(KEYINPUT89), .A3(new_n638), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n516), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n639), .B1(new_n681), .B2(new_n685), .ZN(new_n704));
  AOI22_X1  g0504(.A1(new_n703), .A2(new_n704), .B1(new_n572), .B2(new_n637), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n651), .A2(KEYINPUT26), .A3(new_n561), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n706), .B1(new_n658), .B2(KEYINPUT26), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n678), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT29), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n709), .B(new_n682), .C1(new_n650), .C2(new_n659), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(G330), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT30), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n617), .A2(new_n620), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n716), .A2(new_n553), .A3(new_n554), .A4(new_n600), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n715), .B1(new_n717), .B2(new_n521), .ZN(new_n718));
  AND4_X1   g0518(.A1(new_n496), .A2(new_n491), .A3(new_n520), .A4(new_n504), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n600), .A2(new_n617), .A3(new_n620), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n592), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n719), .A2(new_n721), .A3(KEYINPUT30), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n600), .A2(G179), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n505), .A2(new_n723), .A3(new_n592), .A4(new_n621), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n718), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n678), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(KEYINPUT31), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT31), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n725), .A2(new_n728), .A3(new_n678), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n523), .A2(new_n635), .A3(new_n682), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n714), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n713), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n700), .B1(new_n735), .B2(G1), .ZN(G364));
  NOR2_X1   g0536(.A1(G13), .A2(G33), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G20), .ZN(new_n739));
  XOR2_X1   g0539(.A(new_n739), .B(KEYINPUT95), .Z(new_n740));
  NAND3_X1  g0540(.A1(new_n686), .A2(new_n687), .A3(new_n740), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n266), .A2(new_n267), .B1(new_n225), .B2(G169), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n742), .A2(KEYINPUT93), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(KEYINPUT93), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n225), .A2(G190), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n438), .A2(G179), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n211), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G179), .A2(G200), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G159), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT32), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n225), .B1(new_n750), .B2(G190), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G97), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n367), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n746), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n367), .A2(new_n438), .ZN(new_n760));
  AND2_X1   g0560(.A1(new_n760), .A2(new_n746), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI221_X1 g0562(.A(new_n757), .B1(new_n217), .B2(new_n759), .C1(new_n762), .C2(new_n209), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n225), .A2(new_n351), .ZN(new_n764));
  AND2_X1   g0564(.A1(new_n764), .A2(new_n760), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n259), .B1(new_n766), .B2(new_n215), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n754), .A2(new_n763), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n764), .A2(new_n747), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n768), .B1(new_n566), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n764), .A2(new_n758), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n749), .B(new_n770), .C1(G58), .C2(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(KEYINPUT94), .B(G326), .ZN(new_n774));
  XNOR2_X1  g0574(.A(KEYINPUT33), .B(G317), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n765), .A2(new_n774), .B1(new_n761), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n756), .A2(G294), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n752), .A2(G329), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n776), .A2(new_n324), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G311), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n759), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G283), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n748), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G303), .ZN(new_n784));
  INV_X1    g0584(.A(G322), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n784), .A2(new_n769), .B1(new_n771), .B2(new_n785), .ZN(new_n786));
  NOR4_X1   g0586(.A1(new_n779), .A2(new_n781), .A3(new_n783), .A4(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n745), .B1(new_n773), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n693), .A2(new_n259), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(new_n579), .B2(new_n232), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(new_n250), .B2(new_n579), .ZN(new_n792));
  NAND3_X1  g0592(.A1(G355), .A2(new_n205), .A3(new_n259), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n792), .B(new_n793), .C1(G116), .C2(new_n205), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n745), .A2(new_n739), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(G13), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(G20), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n252), .B1(new_n798), .B2(G45), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n696), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n741), .A2(new_n788), .A3(new_n796), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n689), .A2(new_n800), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n688), .A2(G330), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(G396));
  NOR2_X1   g0605(.A1(new_n396), .A2(new_n678), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n393), .A2(new_n678), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n807), .A2(KEYINPUT97), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(KEYINPUT97), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n808), .B(new_n809), .C1(new_n437), .C2(new_n439), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n806), .B1(new_n810), .B2(new_n396), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n660), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n812), .B1(new_n813), .B2(new_n678), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n682), .B(new_n811), .C1(new_n650), .C2(new_n659), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n800), .B1(new_n816), .B2(new_n733), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(KEYINPUT98), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT98), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n819), .B(new_n800), .C1(new_n816), .C2(new_n733), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n816), .A2(new_n733), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n818), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT99), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n757), .B1(new_n211), .B2(new_n769), .C1(new_n780), .C2(new_n751), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n324), .B1(new_n771), .B2(new_n494), .ZN(new_n825));
  INV_X1    g0625(.A(G87), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n826), .A2(new_n748), .B1(new_n759), .B2(new_n605), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n824), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n828), .B1(new_n782), .B2(new_n762), .C1(new_n784), .C2(new_n766), .ZN(new_n829));
  INV_X1    g0629(.A(new_n759), .ZN(new_n830));
  AOI22_X1  g0630(.A1(G143), .A2(new_n772), .B1(new_n830), .B2(G159), .ZN(new_n831));
  INV_X1    g0631(.A(G137), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n831), .B1(new_n832), .B2(new_n766), .C1(new_n413), .C2(new_n762), .ZN(new_n833));
  XOR2_X1   g0633(.A(KEYINPUT96), .B(KEYINPUT34), .Z(new_n834));
  NOR2_X1   g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n769), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n835), .B1(G50), .B2(new_n836), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n837), .B1(new_n220), .B2(new_n755), .C1(new_n209), .C2(new_n748), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n833), .A2(new_n834), .B1(G132), .B2(new_n752), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n259), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n829), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n745), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n745), .A2(new_n737), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n800), .B1(new_n843), .B2(new_n217), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n842), .B(new_n844), .C1(new_n811), .C2(new_n738), .ZN(new_n845));
  AND3_X1   g0645(.A1(new_n822), .A2(new_n823), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n823), .B1(new_n822), .B2(new_n845), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(G384));
  NAND2_X1  g0649(.A1(new_n730), .A2(new_n731), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n452), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n851), .B(KEYINPUT100), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n342), .A2(new_n294), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n355), .ZN(new_n854));
  INV_X1    g0654(.A(new_n676), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n444), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n372), .A2(new_n373), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n373), .A2(new_n855), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT37), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n859), .A2(new_n860), .A3(new_n861), .A4(new_n363), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n854), .A2(new_n368), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n363), .A2(new_n856), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n862), .B1(new_n864), .B2(new_n861), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT38), .B1(new_n858), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n858), .A2(KEYINPUT38), .A3(new_n865), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n311), .A2(new_n678), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n445), .A2(new_n446), .A3(new_n870), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n311), .B(new_n678), .C1(new_n310), .C2(new_n317), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n850), .A2(new_n811), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT40), .B1(new_n869), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT38), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n860), .B1(new_n365), .B2(new_n664), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n860), .A2(new_n363), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT37), .B1(new_n878), .B2(new_n663), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n879), .A2(new_n862), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n876), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n868), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n882), .A2(KEYINPUT40), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n875), .B1(new_n874), .B2(new_n883), .ZN(new_n884));
  XOR2_X1   g0684(.A(new_n852), .B(new_n884), .Z(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(G330), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT39), .B1(new_n881), .B2(new_n868), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n445), .A2(new_n678), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n867), .A2(KEYINPUT39), .A3(new_n868), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n873), .ZN(new_n892));
  INV_X1    g0692(.A(new_n806), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n892), .B1(new_n815), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n869), .ZN(new_n895));
  OR2_X1    g0695(.A1(new_n664), .A2(new_n855), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n891), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n452), .B1(new_n710), .B2(new_n712), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n670), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n897), .B(new_n899), .Z(new_n900));
  XNOR2_X1  g0700(.A(new_n886), .B(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n252), .B2(new_n798), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n531), .A2(new_n533), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n605), .B1(new_n903), .B2(KEYINPUT35), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n904), .B(new_n230), .C1(KEYINPUT35), .C2(new_n903), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT36), .ZN(new_n906));
  OAI21_X1  g0706(.A(G77), .B1(new_n220), .B2(new_n209), .ZN(new_n907));
  OAI22_X1  g0707(.A1(new_n907), .A2(new_n231), .B1(G50), .B2(new_n209), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(G1), .A3(new_n797), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n902), .A2(new_n906), .A3(new_n909), .ZN(G367));
  OR2_X1    g0710(.A1(new_n597), .A2(new_n682), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n647), .B2(new_n648), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n911), .A2(new_n638), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n914), .A2(KEYINPUT43), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n915), .B(KEYINPUT101), .Z(new_n916));
  NOR2_X1   g0716(.A1(new_n916), .A2(KEYINPUT102), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n685), .A2(new_n678), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n679), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n640), .B1(new_n591), .B2(new_n682), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT42), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n657), .A2(new_n678), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n681), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n561), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n682), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n914), .A2(KEYINPUT43), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n916), .A2(KEYINPUT102), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n917), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AOI211_X1 g0731(.A(KEYINPUT102), .B(new_n916), .C1(new_n927), .C2(new_n928), .ZN(new_n932));
  INV_X1    g0732(.A(new_n690), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n920), .A2(new_n923), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OR3_X1    g0735(.A1(new_n931), .A2(new_n932), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n935), .B1(new_n931), .B2(new_n932), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n696), .B(KEYINPUT41), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n934), .A2(KEYINPUT45), .A3(new_n691), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT45), .B1(new_n934), .B2(new_n691), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n691), .A2(new_n640), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT44), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n943), .B(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT103), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n690), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n946), .A2(KEYINPUT103), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(KEYINPUT104), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n684), .B(new_n689), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(new_n918), .Z(new_n954));
  NOR2_X1   g0754(.A1(new_n954), .A2(new_n734), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT104), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n949), .A2(new_n956), .A3(new_n950), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n946), .A2(new_n690), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n952), .A2(new_n955), .A3(new_n957), .A4(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n938), .B1(new_n959), .B2(new_n735), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n799), .B(KEYINPUT105), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n936), .B(new_n937), .C1(new_n960), .C2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n914), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n800), .B1(new_n963), .B2(new_n740), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n795), .B1(new_n205), .B2(new_n389), .C1(new_n240), .C2(new_n790), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT46), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n769), .B2(new_n605), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n967), .A2(KEYINPUT106), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n836), .A2(KEYINPUT46), .A3(G116), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n761), .A2(G294), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n967), .A2(KEYINPUT106), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n968), .A2(new_n969), .A3(new_n970), .A4(new_n971), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n972), .A2(KEYINPUT107), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(KEYINPUT107), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n771), .A2(new_n784), .B1(new_n759), .B2(new_n782), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n259), .B(new_n975), .C1(G311), .C2(new_n765), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n973), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(G317), .B2(new_n752), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n978), .B1(new_n243), .B2(new_n748), .C1(new_n211), .C2(new_n755), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT108), .ZN(new_n980));
  XNOR2_X1  g0780(.A(KEYINPUT109), .B(G137), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n259), .B1(new_n982), .B2(new_n751), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n772), .A2(G150), .B1(new_n765), .B2(G143), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n984), .B1(new_n215), .B2(new_n759), .C1(new_n209), .C2(new_n755), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(G58), .B2(new_n836), .ZN(new_n986));
  INV_X1    g0786(.A(new_n748), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(G77), .ZN(new_n988));
  INV_X1    g0788(.A(G159), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n986), .B(new_n988), .C1(new_n989), .C2(new_n762), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n980), .B1(new_n983), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT47), .Z(new_n992));
  INV_X1    g0792(.A(new_n745), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n964), .B(new_n965), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n962), .A2(new_n994), .ZN(G387));
  INV_X1    g0795(.A(new_n353), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n215), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT50), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n209), .A2(new_n217), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n567), .A2(new_n605), .ZN(new_n1000));
  NOR4_X1   g0800(.A1(new_n998), .A2(G45), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n789), .B1(new_n237), .B2(new_n579), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1000), .A2(new_n205), .A3(new_n259), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1001), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n205), .A2(G107), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n795), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n800), .B1(new_n684), .B2(new_n740), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n766), .A2(new_n989), .B1(new_n755), .B2(new_n389), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n324), .B1(new_n752), .B2(G150), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n217), .B2(new_n769), .C1(new_n243), .C2(new_n748), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT110), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n1008), .B(new_n1011), .C1(G50), .C2(new_n772), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1012), .B1(new_n209), .B2(new_n759), .C1(new_n353), .C2(new_n762), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(G322), .A2(new_n765), .B1(new_n761), .B2(G311), .ZN(new_n1014));
  INV_X1    g0814(.A(G317), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1014), .B1(new_n784), .B2(new_n759), .C1(new_n1015), .C2(new_n771), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT48), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1017), .B1(new_n782), .B2(new_n755), .C1(new_n494), .C2(new_n769), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT49), .Z(new_n1019));
  AOI21_X1  g0819(.A(new_n259), .B1(new_n987), .B2(G116), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n752), .A2(new_n774), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1013), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT111), .Z(new_n1024));
  OAI211_X1 g0824(.A(new_n1006), .B(new_n1007), .C1(new_n1024), .C2(new_n993), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT112), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n961), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n696), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n954), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1028), .B1(new_n1029), .B2(new_n735), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1026), .B1(new_n954), .B2(new_n1027), .C1(new_n1030), .C2(new_n955), .ZN(G393));
  INV_X1    g0831(.A(new_n958), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n946), .A2(new_n690), .ZN(new_n1033));
  NOR3_X1   g0833(.A1(new_n1032), .A2(new_n1027), .A3(new_n1033), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n954), .A2(new_n734), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n959), .A2(new_n1028), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT114), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n959), .A2(KEYINPUT114), .A3(new_n1028), .A4(new_n1035), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1034), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n748), .A2(new_n211), .B1(new_n751), .B2(new_n785), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n324), .B1(new_n782), .B2(new_n769), .C1(new_n762), .C2(new_n784), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1041), .B(new_n1042), .C1(G294), .C2(new_n830), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n605), .B2(new_n755), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n772), .A2(G311), .B1(new_n765), .B2(G317), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT52), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n755), .A2(new_n217), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n766), .A2(new_n413), .B1(new_n771), .B2(new_n989), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT51), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n752), .A2(G143), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n324), .B1(new_n987), .B2(G87), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n769), .A2(new_n209), .B1(new_n759), .B2(new_n353), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(G50), .B2(new_n761), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .A4(new_n1053), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n1044), .A2(new_n1046), .B1(new_n1047), .B2(new_n1054), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT113), .Z(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n745), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n920), .A2(new_n739), .A3(new_n923), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n795), .B1(new_n243), .B2(new_n205), .C1(new_n247), .C2(new_n790), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1057), .A2(new_n801), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1040), .A2(new_n1060), .ZN(G390));
  INV_X1    g0861(.A(KEYINPUT119), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n815), .A2(new_n893), .ZN(new_n1063));
  AND4_X1   g0863(.A1(G330), .A2(new_n850), .A3(new_n811), .A4(new_n873), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n873), .B1(new_n732), .B2(new_n811), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1063), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(KEYINPUT117), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1064), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n810), .A2(new_n396), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n806), .B1(new_n708), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1065), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1068), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT117), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1063), .B(new_n1073), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1067), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n452), .A2(G330), .A3(new_n850), .ZN(new_n1076));
  AND3_X1   g0876(.A1(new_n898), .A2(new_n1076), .A3(new_n670), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(KEYINPUT118), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT118), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1075), .A2(new_n1077), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n868), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT39), .ZN(new_n1083));
  NOR3_X1   g0883(.A1(new_n1082), .A2(new_n866), .A3(new_n1083), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n1084), .A2(new_n887), .B1(new_n894), .B2(new_n889), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1064), .A2(KEYINPUT116), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n889), .B1(new_n881), .B2(new_n868), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n1070), .B2(new_n892), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1085), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(KEYINPUT116), .B1(new_n1064), .B2(KEYINPUT115), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1090), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1085), .A2(new_n1092), .A3(new_n1088), .A4(new_n1086), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1079), .A2(new_n1081), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1062), .B1(new_n1094), .B2(new_n696), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1097));
  OR2_X1    g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n1075), .A2(new_n1080), .A3(new_n1077), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1080), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1097), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1101), .A2(KEYINPUT119), .A3(new_n1028), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1095), .A2(new_n1098), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1097), .A2(new_n961), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n737), .B1(new_n1084), .B2(new_n887), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n494), .A2(new_n751), .B1(new_n755), .B2(new_n217), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n766), .A2(new_n782), .B1(new_n748), .B2(new_n209), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1106), .B(new_n1107), .C1(G97), .C2(new_n830), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n259), .B1(new_n772), .B2(G116), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n1110), .B1(new_n826), .B2(new_n769), .C1(new_n211), .C2(new_n762), .ZN(new_n1111));
  INV_X1    g0911(.A(G125), .ZN(new_n1112));
  INV_X1    g0912(.A(G132), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n259), .B1(new_n751), .B2(new_n1112), .C1(new_n1113), .C2(new_n771), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n836), .A2(G150), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT53), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n1114), .B(new_n1116), .C1(G159), .C2(new_n756), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(G50), .A2(new_n987), .B1(new_n765), .B2(G128), .ZN(new_n1118));
  XOR2_X1   g0918(.A(KEYINPUT54), .B(G143), .Z(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1117), .B(new_n1118), .C1(new_n759), .C2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n762), .A2(new_n982), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1111), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n800), .B1(new_n1123), .B2(new_n745), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n843), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1124), .B1(new_n996), .B2(new_n1125), .ZN(new_n1126));
  XOR2_X1   g0926(.A(new_n1126), .B(KEYINPUT120), .Z(new_n1127));
  NAND2_X1  g0927(.A1(new_n1105), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1104), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1103), .A2(new_n1130), .ZN(G378));
  INV_X1    g0931(.A(KEYINPUT57), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n898), .A2(new_n1076), .A3(new_n670), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1094), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n875), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n882), .A2(KEYINPUT40), .A3(new_n874), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1135), .A2(G330), .A3(new_n1136), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1137), .A2(new_n895), .A3(new_n896), .A4(new_n891), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n897), .A2(new_n884), .A3(G330), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n435), .ZN(new_n1141));
  OR2_X1    g0941(.A1(new_n1141), .A2(KEYINPUT122), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(KEYINPUT122), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n416), .A2(new_n676), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n1142), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1145), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1140), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1138), .A2(new_n1152), .A3(new_n1139), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1132), .B1(new_n1134), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1101), .A2(new_n1077), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1158), .A2(KEYINPUT57), .A3(new_n1155), .A4(new_n1154), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1157), .A2(new_n1159), .A3(new_n1028), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1152), .A2(new_n738), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n215), .B1(new_n322), .B2(G41), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n759), .A2(new_n832), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n766), .A2(new_n1112), .B1(new_n755), .B2(new_n413), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT121), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1163), .B(new_n1165), .C1(new_n836), .C2(new_n1119), .ZN(new_n1166));
  INV_X1    g0966(.A(G128), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n1166), .B1(new_n1167), .B2(new_n771), .C1(new_n1113), .C2(new_n762), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n987), .A2(G159), .ZN(new_n1170));
  AOI21_X1  g0970(.A(G41), .B1(new_n752), .B2(G124), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1169), .A2(new_n263), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1162), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n217), .A2(new_n769), .B1(new_n771), .B2(new_n211), .ZN(new_n1175));
  AOI211_X1 g0975(.A(G41), .B(new_n1175), .C1(G68), .C2(new_n756), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n259), .B1(new_n987), .B2(G58), .ZN(new_n1177));
  OR2_X1    g0977(.A1(new_n759), .A2(new_n389), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(G97), .A2(new_n761), .B1(new_n752), .B2(G283), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(G116), .B2(new_n765), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT58), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n745), .B1(new_n1174), .B2(new_n1182), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1183), .B(new_n801), .C1(G50), .C2(new_n1125), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n1156), .A2(new_n1027), .B1(new_n1161), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1160), .A2(new_n1186), .ZN(G375));
  NAND2_X1  g0987(.A1(new_n892), .A2(new_n737), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n748), .A2(new_n220), .B1(new_n751), .B2(new_n1167), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n324), .B(new_n1189), .C1(G50), .C2(new_n756), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1190), .B1(new_n413), .B2(new_n759), .C1(new_n989), .C2(new_n769), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT123), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n772), .A2(new_n981), .B1(new_n765), .B2(G132), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1192), .B(new_n1193), .C1(new_n762), .C2(new_n1120), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n988), .B1(new_n766), .B2(new_n494), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n324), .B1(new_n759), .B2(new_n211), .C1(new_n243), .C2(new_n769), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n755), .A2(new_n389), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n751), .A2(new_n784), .ZN(new_n1198));
  NOR4_X1   g0998(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1199), .B1(new_n605), .B2(new_n762), .C1(new_n782), .C2(new_n771), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n993), .B1(new_n1194), .B2(new_n1200), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n800), .B(new_n1201), .C1(new_n209), .C2(new_n843), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1075), .A2(new_n961), .B1(new_n1188), .B2(new_n1202), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1133), .A2(new_n1072), .A3(new_n1067), .A4(new_n1074), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n938), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1203), .B1(new_n1096), .B2(new_n1206), .ZN(new_n1207));
  XOR2_X1   g1007(.A(new_n1207), .B(KEYINPUT124), .Z(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(G381));
  NOR4_X1   g1009(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n1101), .A2(KEYINPUT119), .A3(new_n1028), .ZN(new_n1211));
  AOI21_X1  g1011(.A(KEYINPUT119), .B1(new_n1101), .B2(new_n1028), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(KEYINPUT125), .B1(new_n1214), .B2(new_n1129), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT125), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1103), .A2(new_n1216), .A3(new_n1130), .ZN(new_n1217));
  AOI21_X1  g1017(.A(G375), .B1(new_n1215), .B2(new_n1217), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1040), .A2(new_n962), .A3(new_n994), .A4(new_n1060), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1210), .A2(new_n1218), .A3(new_n1220), .ZN(G407));
  INV_X1    g1021(.A(G213), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n1218), .B2(new_n677), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(G407), .ZN(G409));
  NOR2_X1   g1024(.A1(new_n1222), .A2(G343), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1096), .A2(new_n1204), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1204), .A2(KEYINPUT126), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(KEYINPUT60), .ZN(new_n1229));
  OR2_X1    g1029(.A1(new_n1228), .A2(KEYINPUT60), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1227), .A2(new_n1028), .A3(new_n1229), .A4(new_n1230), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1231), .A2(new_n848), .A3(new_n1203), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n848), .B1(new_n1231), .B2(new_n1203), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1134), .A2(new_n1156), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1185), .B1(new_n1205), .B2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n1215), .B2(new_n1217), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1160), .A2(G378), .A3(new_n1186), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1226), .B(new_n1235), .C1(new_n1238), .C2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(KEYINPUT62), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1226), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1225), .A2(G2897), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1231), .A2(new_n1203), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(G384), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1231), .A2(new_n848), .A3(new_n1203), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1247), .A2(new_n1248), .A3(new_n1243), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1245), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1242), .A2(new_n1251), .ZN(new_n1252));
  XOR2_X1   g1052(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1253));
  NAND2_X1  g1053(.A1(new_n1236), .A2(new_n1205), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n1186), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1103), .A2(new_n1216), .A3(new_n1130), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1216), .B1(new_n1103), .B2(new_n1130), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1255), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1160), .A2(G378), .A3(new_n1186), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT62), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1260), .A2(new_n1261), .A3(new_n1226), .A4(new_n1235), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1241), .A2(new_n1252), .A3(new_n1253), .A4(new_n1262), .ZN(new_n1263));
  XOR2_X1   g1063(.A(G393), .B(G396), .Z(new_n1264));
  AOI22_X1  g1064(.A1(new_n1040), .A2(new_n1060), .B1(new_n962), .B2(new_n994), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1264), .B1(new_n1220), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(G390), .A2(G387), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1264), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1267), .A2(new_n1268), .A3(new_n1219), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1266), .A2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1263), .A2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1250), .B1(new_n1260), .B2(new_n1226), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT63), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1240), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  AOI211_X1 g1074(.A(new_n1225), .B(new_n1234), .C1(new_n1258), .C2(new_n1259), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1270), .B1(new_n1275), .B2(KEYINPUT63), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT61), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1274), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1271), .A2(new_n1278), .ZN(G405));
  INV_X1    g1079(.A(new_n1269), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1268), .B1(new_n1267), .B2(new_n1219), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1234), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1266), .A2(new_n1269), .A3(new_n1235), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1239), .B1(G375), .B2(new_n1285), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(new_n1284), .B(new_n1286), .ZN(G402));
endmodule


