//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 0 0 1 1 1 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 1 1 1 1 0 1 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063;
  XNOR2_X1  g000(.A(KEYINPUT2), .B(G113), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G116), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  AND2_X1   g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n188), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n190), .A2(new_n192), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(new_n187), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n199), .A2(new_n201), .A3(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n198), .B1(new_n201), .B2(KEYINPUT1), .ZN(new_n205));
  XNOR2_X1  g019(.A(G143), .B(G146), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT11), .ZN(new_n208));
  INV_X1    g022(.A(G134), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n208), .B1(new_n209), .B2(G137), .ZN(new_n210));
  INV_X1    g024(.A(G137), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(KEYINPUT11), .A3(G134), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n209), .A2(G137), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n210), .A2(new_n212), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n209), .A2(G137), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n211), .A2(G134), .ZN(new_n217));
  OAI21_X1  g031(.A(G131), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n197), .B1(new_n207), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n210), .A2(new_n212), .A3(new_n214), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G131), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n215), .ZN(new_n224));
  AND2_X1   g038(.A1(KEYINPUT0), .A2(G128), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n201), .A2(new_n203), .A3(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT0), .B(G128), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n226), .B1(new_n206), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n224), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(KEYINPUT28), .B1(new_n221), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT1), .B1(new_n202), .B2(G146), .ZN(new_n233));
  AOI22_X1  g047(.A1(new_n233), .A2(G128), .B1(new_n201), .B2(new_n203), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n199), .A2(new_n201), .A3(new_n203), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT64), .B1(new_n236), .B2(new_n219), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT64), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n207), .A2(new_n238), .A3(new_n215), .A4(new_n218), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n237), .A2(new_n230), .A3(new_n239), .ZN(new_n240));
  AND2_X1   g054(.A1(new_n240), .A2(new_n197), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n230), .A2(KEYINPUT65), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT65), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n224), .A2(new_n243), .A3(new_n229), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n242), .A2(new_n221), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT66), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n242), .A2(new_n221), .A3(KEYINPUT66), .A4(new_n244), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n241), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT28), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n232), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G237), .ZN(new_n252));
  INV_X1    g066(.A(G953), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n253), .A3(G210), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n254), .B(KEYINPUT27), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT26), .B(G101), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XOR2_X1   g071(.A(new_n257), .B(KEYINPUT68), .Z(new_n258));
  NAND2_X1  g072(.A1(new_n251), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n247), .A2(new_n248), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n220), .A2(new_n207), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n242), .A2(KEYINPUT30), .A3(new_n261), .A4(new_n244), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT30), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n240), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n262), .A2(new_n264), .A3(new_n197), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n260), .A2(new_n257), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT31), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n266), .A2(KEYINPUT67), .A3(KEYINPUT31), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT67), .B1(new_n266), .B2(KEYINPUT31), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n259), .B(new_n269), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(G472), .A2(G902), .ZN(new_n273));
  XOR2_X1   g087(.A(new_n273), .B(KEYINPUT69), .Z(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT32), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n274), .A2(new_n277), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n272), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT71), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n260), .A2(new_n265), .ZN(new_n282));
  INV_X1    g096(.A(new_n257), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT29), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n258), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n232), .B(new_n285), .C1(new_n249), .C2(new_n250), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT70), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n284), .A2(new_n286), .A3(new_n289), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n257), .A2(KEYINPUT29), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n242), .A2(new_n261), .A3(new_n244), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n247), .A2(new_n248), .B1(new_n197), .B2(new_n292), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n232), .B(new_n291), .C1(new_n293), .C2(new_n250), .ZN(new_n294));
  INV_X1    g108(.A(G902), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n288), .A2(new_n290), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G472), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT71), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n272), .A2(new_n300), .A3(new_n279), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n278), .A2(new_n281), .A3(new_n299), .A4(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT9), .B(G234), .ZN(new_n303));
  OAI21_X1  g117(.A(G221), .B1(new_n303), .B2(G902), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G469), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n306), .A2(new_n295), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n207), .A2(KEYINPUT10), .ZN(new_n308));
  INV_X1    g122(.A(G107), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G104), .ZN(new_n310));
  INV_X1    g124(.A(G104), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G107), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G101), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT3), .B1(new_n311), .B2(G107), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT3), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(new_n309), .A3(G104), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n315), .A2(new_n317), .A3(new_n312), .ZN(new_n318));
  XOR2_X1   g132(.A(KEYINPUT80), .B(G101), .Z(new_n319));
  OAI21_X1  g133(.A(new_n314), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n308), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n206), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT83), .ZN(new_n323));
  OAI21_X1  g137(.A(G128), .B1(new_n233), .B2(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(KEYINPUT83), .B1(new_n201), .B2(KEYINPUT1), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n322), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n204), .ZN(new_n327));
  INV_X1    g141(.A(new_n320), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT10), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n321), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT4), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n315), .A2(new_n317), .A3(new_n312), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT80), .B(G101), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n318), .A2(G101), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n228), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT82), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n318), .A2(new_n332), .A3(G101), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT81), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n318), .A2(KEYINPUT81), .A3(new_n332), .A4(G101), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n337), .A2(new_n338), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n338), .B1(new_n337), .B2(new_n343), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n331), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n224), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n253), .A2(G227), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n348), .B(KEYINPUT79), .ZN(new_n349));
  XNOR2_X1  g163(.A(G110), .B(G140), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n349), .B(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n320), .B1(new_n326), .B2(new_n204), .ZN(new_n352));
  OAI22_X1  g166(.A1(new_n352), .A2(KEYINPUT10), .B1(new_n320), .B2(new_n308), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n341), .A2(new_n342), .ZN(new_n354));
  INV_X1    g168(.A(new_n336), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT4), .B1(new_n318), .B2(new_n319), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n229), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT82), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n337), .A2(new_n338), .A3(new_n343), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n353), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  XOR2_X1   g174(.A(new_n224), .B(KEYINPUT84), .Z(new_n361));
  AOI21_X1  g175(.A(new_n351), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n331), .B(new_n361), .C1(new_n344), .C2(new_n345), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n333), .A2(new_n334), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n207), .B1(new_n364), .B2(new_n314), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n224), .B1(new_n352), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT12), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g182(.A(KEYINPUT12), .B(new_n224), .C1(new_n352), .C2(new_n365), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n363), .A2(new_n370), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n347), .A2(new_n362), .B1(new_n371), .B2(new_n351), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n307), .B1(new_n372), .B2(G469), .ZN(new_n373));
  INV_X1    g187(.A(new_n351), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n374), .B1(new_n347), .B2(new_n363), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n363), .A2(new_n370), .A3(new_n374), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n306), .B(new_n295), .C1(new_n375), .C2(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n305), .B1(new_n373), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n198), .A2(KEYINPUT23), .A3(G119), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n189), .A2(G128), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n189), .A2(G128), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n381), .B(new_n382), .C1(new_n383), .C2(KEYINPUT23), .ZN(new_n384));
  XNOR2_X1  g198(.A(G119), .B(G128), .ZN(new_n385));
  INV_X1    g199(.A(G110), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT24), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT24), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G110), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n384), .A2(G110), .B1(new_n385), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G140), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G125), .ZN(new_n393));
  INV_X1    g207(.A(G125), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G140), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(new_n395), .A3(KEYINPUT16), .ZN(new_n396));
  OR3_X1    g210(.A1(new_n394), .A2(KEYINPUT16), .A3(G140), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(G146), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(G146), .B1(new_n396), .B2(new_n397), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n391), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(KEYINPUT73), .B(G110), .ZN(new_n402));
  OAI22_X1  g216(.A1(new_n384), .A2(new_n402), .B1(new_n385), .B2(new_n390), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n393), .A2(new_n395), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT74), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT74), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n393), .A2(new_n395), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n405), .A2(new_n200), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n403), .A2(new_n408), .A3(new_n398), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT22), .B(G137), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n253), .A2(G221), .A3(G234), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n410), .B(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT75), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n410), .B(new_n411), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT75), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n401), .A2(new_n409), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n401), .A2(new_n409), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n418), .A2(KEYINPUT76), .B1(new_n420), .B2(new_n416), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n415), .A2(new_n417), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT76), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  XOR2_X1   g240(.A(KEYINPUT72), .B(G217), .Z(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G234), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n428), .B1(new_n429), .B2(G902), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n295), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(KEYINPUT77), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n426), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n433), .B(KEYINPUT78), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n420), .A2(new_n416), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n419), .A2(new_n422), .A3(KEYINPUT76), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n425), .A2(new_n435), .A3(new_n295), .A4(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT25), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n421), .A2(KEYINPUT25), .A3(new_n295), .A4(new_n425), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n430), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n434), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(G210), .B1(G237), .B2(G902), .ZN(new_n445));
  XOR2_X1   g259(.A(new_n445), .B(KEYINPUT89), .Z(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n190), .A2(new_n192), .A3(KEYINPUT5), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT5), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(new_n189), .A3(G116), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT85), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n449), .A2(new_n189), .A3(KEYINPUT85), .A4(G116), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n448), .A2(new_n452), .A3(G113), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n194), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n455), .A2(new_n320), .ZN(new_n456));
  AOI22_X1  g270(.A1(new_n335), .A2(new_n336), .B1(new_n194), .B2(new_n196), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n456), .B1(new_n457), .B2(new_n343), .ZN(new_n458));
  XNOR2_X1  g272(.A(G110), .B(G122), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n458), .A2(KEYINPUT6), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n207), .A2(new_n394), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n226), .B(G125), .C1(new_n206), .C2(new_n227), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(G224), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(G953), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n463), .B(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n328), .A2(new_n194), .A3(new_n454), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n197), .B1(new_n355), .B2(new_n356), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n467), .B(new_n459), .C1(new_n354), .C2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT86), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n458), .A2(KEYINPUT86), .A3(new_n459), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT6), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n467), .B1(new_n354), .B2(new_n468), .ZN(new_n475));
  INV_X1    g289(.A(new_n459), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI211_X1 g291(.A(new_n460), .B(new_n466), .C1(new_n473), .C2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT7), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n461), .B(new_n462), .C1(new_n479), .C2(new_n465), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT87), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n461), .A2(new_n462), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT87), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n482), .B(new_n483), .C1(new_n479), .C2(new_n465), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT88), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n479), .B1(new_n465), .B2(new_n485), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n463), .B(new_n486), .C1(new_n485), .C2(new_n465), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n459), .B(KEYINPUT8), .ZN(new_n488));
  AOI22_X1  g302(.A1(new_n364), .A2(new_n314), .B1(new_n454), .B2(new_n194), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n488), .B1(new_n456), .B2(new_n489), .ZN(new_n490));
  AND4_X1   g304(.A1(new_n481), .A2(new_n484), .A3(new_n487), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n473), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n295), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n447), .B1(new_n478), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n460), .B1(new_n473), .B2(new_n477), .ZN(new_n495));
  INV_X1    g309(.A(new_n466), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(G902), .B1(new_n473), .B2(new_n491), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(new_n446), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(G214), .B1(G237), .B2(G902), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n494), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NOR3_X1   g315(.A1(new_n380), .A2(new_n444), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT93), .ZN(new_n503));
  XNOR2_X1  g317(.A(G113), .B(G122), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(new_n311), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT19), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n405), .A2(new_n506), .A3(new_n407), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n404), .A2(KEYINPUT19), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(new_n200), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n398), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT91), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n252), .A2(new_n253), .A3(G214), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n202), .A2(KEYINPUT90), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT90), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n514), .A2(G143), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n512), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g330(.A1(G237), .A2(G953), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n517), .B(G214), .C1(new_n514), .C2(G143), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n213), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n516), .A2(new_n213), .A3(new_n518), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT91), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n509), .A2(new_n523), .A3(new_n398), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n511), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n404), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n408), .B1(new_n200), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n519), .A2(KEYINPUT18), .ZN(new_n528));
  NAND2_X1  g342(.A1(KEYINPUT18), .A2(G131), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n516), .A2(new_n518), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n505), .B1(new_n525), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT17), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n520), .A2(new_n533), .A3(new_n521), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n399), .A2(new_n400), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT92), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n519), .A2(new_n536), .A3(KEYINPUT17), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n536), .B1(new_n519), .B2(KEYINPUT17), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n534), .B(new_n535), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(new_n505), .A3(new_n531), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n503), .B1(new_n532), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(G475), .A2(G902), .ZN(new_n543));
  INV_X1    g357(.A(new_n531), .ZN(new_n544));
  AOI22_X1  g358(.A1(new_n510), .A2(KEYINPUT91), .B1(new_n520), .B2(new_n521), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n544), .B1(new_n545), .B2(new_n524), .ZN(new_n546));
  OAI211_X1 g360(.A(KEYINPUT93), .B(new_n540), .C1(new_n546), .C2(new_n505), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n542), .A2(new_n543), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n540), .B1(new_n546), .B2(new_n505), .ZN(new_n549));
  NOR3_X1   g363(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n548), .A2(KEYINPUT20), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(G475), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n505), .B1(new_n539), .B2(new_n531), .ZN(new_n553));
  OR2_X1    g367(.A1(new_n541), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n552), .B1(new_n554), .B2(new_n295), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(G122), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(G116), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n309), .B1(new_n558), .B2(KEYINPUT14), .ZN(new_n559));
  XNOR2_X1  g373(.A(G116), .B(G122), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n202), .A2(G128), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n198), .A2(G143), .ZN(new_n563));
  AOI21_X1  g377(.A(KEYINPUT95), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n562), .A2(new_n563), .A3(KEYINPUT95), .ZN(new_n566));
  AOI21_X1  g380(.A(G134), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n566), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n568), .A2(new_n209), .A3(new_n564), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n561), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n209), .B1(new_n568), .B2(new_n564), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n560), .B(new_n309), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT13), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n573), .B1(new_n198), .B2(G143), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n202), .A2(KEYINPUT13), .A3(G128), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(new_n575), .A3(new_n563), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n576), .A2(KEYINPUT94), .A3(G134), .ZN(new_n577));
  AOI21_X1  g391(.A(KEYINPUT94), .B1(new_n576), .B2(G134), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n571), .B(new_n572), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  NOR3_X1   g393(.A1(new_n427), .A2(G953), .A3(new_n303), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n570), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n580), .B1(new_n570), .B2(new_n579), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n295), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(KEYINPUT96), .ZN(new_n584));
  INV_X1    g398(.A(G478), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n585), .A2(KEYINPUT15), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n583), .A2(KEYINPUT96), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n588), .B1(KEYINPUT15), .B2(new_n585), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n253), .A2(G952), .ZN(new_n592));
  NAND2_X1  g406(.A1(G234), .A2(G237), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT21), .B(G898), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n593), .A2(G902), .A3(G953), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n594), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(KEYINPUT97), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n556), .A2(new_n591), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n302), .A2(new_n502), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(new_n319), .ZN(G3));
  NAND2_X1  g417(.A1(new_n266), .A2(KEYINPUT31), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT67), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n266), .A2(KEYINPUT67), .A3(KEYINPUT31), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI22_X1  g422(.A1(new_n251), .A2(new_n258), .B1(new_n267), .B2(new_n268), .ZN(new_n609));
  AOI21_X1  g423(.A(G902), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(G472), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n276), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n612), .A2(new_n444), .A3(new_n380), .ZN(new_n613));
  OR2_X1    g427(.A1(new_n583), .A2(G478), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n585), .A2(new_n295), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  OR3_X1    g431(.A1(new_n581), .A2(new_n582), .A3(KEYINPUT33), .ZN(new_n618));
  OAI21_X1  g432(.A(KEYINPUT33), .B1(new_n581), .B2(new_n582), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n617), .B1(G478), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n621), .B1(new_n551), .B2(new_n555), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n494), .A2(new_n499), .A3(new_n599), .A4(new_n500), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n613), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT34), .B(G104), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G6));
  NAND2_X1  g441(.A1(new_n548), .A2(KEYINPUT20), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT20), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n542), .A2(new_n547), .A3(new_n629), .A4(new_n543), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n555), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n632), .A2(new_n591), .A3(new_n623), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n613), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT35), .B(G107), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G9));
  NOR2_X1   g450(.A1(new_n600), .A2(new_n612), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n494), .A2(new_n499), .A3(new_n500), .ZN(new_n638));
  INV_X1    g452(.A(new_n432), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT98), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n419), .B(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n422), .A2(KEYINPUT36), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n419), .B(KEYINPUT98), .ZN(new_n644));
  INV_X1    g458(.A(new_n642), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n639), .B1(new_n643), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n647), .B1(new_n441), .B2(new_n442), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT99), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n430), .B1(new_n439), .B2(new_n440), .ZN(new_n651));
  OAI21_X1  g465(.A(KEYINPUT99), .B1(new_n651), .B2(new_n647), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n638), .A2(new_n379), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n637), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT37), .B(G110), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT100), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n655), .B(new_n657), .ZN(G12));
  XNOR2_X1  g472(.A(new_n594), .B(KEYINPUT102), .ZN(new_n659));
  NOR2_X1   g473(.A1(KEYINPUT101), .A2(G900), .ZN(new_n660));
  AND2_X1   g474(.A1(KEYINPUT101), .A2(G900), .ZN(new_n661));
  OR3_X1    g475(.A1(new_n597), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n631), .A2(new_n590), .A3(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n302), .A2(new_n654), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G128), .ZN(G30));
  INV_X1    g481(.A(new_n500), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n668), .B1(new_n587), .B2(new_n589), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n669), .B1(new_n551), .B2(new_n555), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n653), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n671), .B(KEYINPUT103), .Z(new_n672));
  OAI21_X1  g486(.A(new_n266), .B1(new_n285), .B2(new_n293), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n295), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(G472), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n278), .A2(new_n281), .A3(new_n301), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n663), .B(KEYINPUT39), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n379), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(KEYINPUT40), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n678), .A2(KEYINPUT40), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n494), .A2(new_n499), .A3(KEYINPUT38), .ZN(new_n681));
  AOI21_X1  g495(.A(KEYINPUT38), .B1(new_n494), .B2(new_n499), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n672), .A2(new_n676), .A3(new_n679), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G143), .ZN(G45));
  OAI211_X1 g500(.A(new_n621), .B(new_n663), .C1(new_n551), .C2(new_n555), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n281), .A2(new_n301), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n284), .A2(new_n289), .A3(new_n286), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n289), .B1(new_n284), .B2(new_n286), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n690), .A2(new_n691), .A3(new_n296), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n274), .B1(new_n608), .B2(new_n609), .ZN(new_n693));
  OAI22_X1  g507(.A1(new_n692), .A2(new_n611), .B1(new_n693), .B2(KEYINPUT32), .ZN(new_n694));
  OAI211_X1 g508(.A(new_n654), .B(new_n688), .C1(new_n689), .C2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G146), .ZN(G48));
  INV_X1    g510(.A(new_n444), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n295), .B1(new_n375), .B2(new_n377), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(G469), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n699), .A2(new_n304), .A3(new_n378), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n302), .A2(new_n624), .A3(new_n697), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT41), .B(G113), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G15));
  NAND4_X1  g518(.A1(new_n302), .A2(new_n697), .A3(new_n633), .A4(new_n701), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G116), .ZN(G18));
  INV_X1    g520(.A(new_n647), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n649), .B1(new_n443), .B2(new_n707), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n651), .A2(KEYINPUT99), .A3(new_n647), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n710), .A2(new_n700), .A3(new_n501), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n302), .A2(new_n601), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G119), .ZN(G21));
  NAND2_X1  g527(.A1(new_n292), .A2(new_n197), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n260), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n231), .B1(new_n715), .B2(KEYINPUT28), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT104), .ZN(new_n717));
  OR2_X1    g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n716), .A2(new_n717), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(new_n258), .A3(new_n719), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n269), .A2(new_n604), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n274), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT105), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n723), .B1(new_n610), .B2(new_n611), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n272), .A2(new_n295), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(KEYINPUT105), .A3(G472), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n722), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n599), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n494), .A2(new_n499), .ZN(new_n729));
  NOR4_X1   g543(.A1(new_n670), .A2(new_n700), .A3(new_n728), .A4(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n727), .A2(new_n730), .A3(new_n697), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  NAND2_X1  g546(.A1(new_n724), .A2(new_n726), .ZN(new_n733));
  INV_X1    g547(.A(new_n722), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n733), .A2(new_n688), .A3(new_n711), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT106), .B(G125), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G27));
  AOI22_X1  g551(.A1(new_n277), .A2(new_n276), .B1(new_n298), .B2(G472), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n444), .B1(new_n738), .B2(new_n280), .ZN(new_n739));
  INV_X1    g553(.A(new_n378), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n347), .A2(new_n363), .A3(new_n374), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n371), .A2(new_n351), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(new_n742), .A3(G469), .ZN(new_n743));
  INV_X1    g557(.A(new_n307), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g559(.A(KEYINPUT107), .B1(new_n740), .B2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT107), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n373), .A2(new_n747), .A3(new_n378), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n668), .B1(new_n494), .B2(new_n499), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n304), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n749), .A2(new_n751), .A3(new_n687), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n739), .A2(new_n752), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n272), .A2(new_n300), .A3(new_n279), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n300), .B1(new_n272), .B2(new_n279), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n444), .B1(new_n756), .B2(new_n738), .ZN(new_n757));
  NOR4_X1   g571(.A1(new_n749), .A2(new_n751), .A3(new_n687), .A4(KEYINPUT42), .ZN(new_n758));
  AOI22_X1  g572(.A1(new_n753), .A2(KEYINPUT42), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G131), .ZN(G33));
  NOR3_X1   g574(.A1(new_n749), .A2(new_n664), .A3(new_n751), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n757), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G134), .ZN(G36));
  NAND2_X1  g577(.A1(new_n741), .A2(new_n742), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n306), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n741), .A2(new_n742), .A3(KEYINPUT45), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n307), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n378), .B1(new_n768), .B2(KEYINPUT46), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n363), .A2(new_n374), .ZN(new_n770));
  INV_X1    g584(.A(new_n224), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n360), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n374), .B1(new_n363), .B2(new_n370), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n765), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(G469), .A3(new_n767), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n744), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT46), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n304), .B(new_n677), .C1(new_n769), .C2(new_n779), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n780), .A2(KEYINPUT108), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(KEYINPUT108), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n549), .A2(new_n550), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n628), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n555), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(new_n621), .A3(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(KEYINPUT43), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT43), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n789), .B1(new_n556), .B2(new_n621), .ZN(new_n790));
  OAI21_X1  g604(.A(KEYINPUT109), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n787), .A2(KEYINPUT43), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n556), .A2(new_n789), .A3(new_n621), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT109), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n693), .B1(G472), .B2(new_n725), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(new_n710), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n791), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(KEYINPUT44), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n729), .A2(new_n500), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n791), .A2(new_n795), .A3(new_n797), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT44), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n783), .A2(new_n799), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G137), .ZN(G39));
  OAI21_X1  g619(.A(new_n304), .B1(new_n769), .B2(new_n779), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT47), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI211_X1 g622(.A(KEYINPUT47), .B(new_n304), .C1(new_n769), .C2(new_n779), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n302), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n697), .A2(new_n687), .A3(new_n800), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G140), .ZN(G42));
  NAND2_X1  g628(.A1(new_n699), .A2(new_n378), .ZN(new_n815));
  AOI211_X1 g629(.A(new_n305), .B(new_n668), .C1(new_n815), .C2(KEYINPUT49), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n816), .B1(KEYINPUT49), .B2(new_n815), .ZN(new_n817));
  NOR4_X1   g631(.A1(new_n817), .A2(new_n681), .A3(new_n682), .A4(new_n787), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n676), .A2(new_n444), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT114), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT110), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n822), .B1(new_n648), .B2(new_n663), .ZN(new_n823));
  INV_X1    g637(.A(new_n663), .ZN(new_n824));
  NOR4_X1   g638(.A1(new_n651), .A2(new_n647), .A3(KEYINPUT110), .A4(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n304), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n749), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n785), .A2(new_n786), .ZN(new_n828));
  INV_X1    g642(.A(new_n729), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(new_n829), .A3(new_n669), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n676), .A2(new_n827), .A3(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n666), .A2(new_n832), .A3(new_n735), .A4(new_n695), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(KEYINPUT52), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n556), .A2(new_n590), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n623), .B1(new_n835), .B2(new_n622), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n613), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n602), .A3(new_n655), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n587), .A2(new_n589), .A3(new_n663), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n839), .B1(new_n650), .B2(new_n652), .ZN(new_n840));
  AND4_X1   g654(.A1(new_n379), .A2(new_n840), .A3(new_n631), .A4(new_n750), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n302), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n302), .A2(new_n697), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n749), .A2(new_n751), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n665), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n842), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n838), .A2(new_n846), .ZN(new_n847));
  AND4_X1   g661(.A1(new_n702), .A2(new_n705), .A3(new_n731), .A4(new_n712), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n752), .A2(new_n727), .A3(new_n653), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n847), .A2(new_n848), .A3(new_n759), .A4(new_n849), .ZN(new_n850));
  XNOR2_X1  g664(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n834), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n757), .A2(new_n761), .B1(new_n302), .B2(new_n841), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n613), .A2(new_n836), .B1(new_n637), .B2(new_n654), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n853), .A2(new_n602), .A3(new_n854), .A4(new_n849), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n753), .A2(KEYINPUT42), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n758), .A2(new_n757), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n702), .A2(new_n705), .A3(new_n731), .A4(new_n712), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n855), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n832), .A2(new_n695), .A3(KEYINPUT52), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n666), .A2(new_n735), .ZN(new_n862));
  OAI21_X1  g676(.A(KEYINPUT111), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n638), .A2(new_n653), .A3(new_n379), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n864), .B1(new_n756), .B2(new_n738), .ZN(new_n865));
  NOR4_X1   g679(.A1(new_n687), .A2(new_n710), .A3(new_n700), .A4(new_n501), .ZN(new_n866));
  AOI22_X1  g680(.A1(new_n865), .A2(new_n665), .B1(new_n866), .B2(new_n727), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT111), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT52), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n830), .A2(new_n749), .A3(new_n826), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n869), .B1(new_n870), .B2(new_n676), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n867), .A2(new_n868), .A3(new_n695), .A4(new_n871), .ZN(new_n872));
  XOR2_X1   g686(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n873));
  NAND2_X1  g687(.A1(new_n833), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n863), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT53), .B1(new_n860), .B2(new_n875), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n821), .B(KEYINPUT54), .C1(new_n852), .C2(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n851), .B1(new_n834), .B2(new_n850), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n860), .A2(KEYINPUT53), .A3(new_n875), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT54), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n863), .A2(new_n872), .A3(new_n874), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n883), .B1(new_n884), .B2(new_n850), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n833), .B(new_n869), .ZN(new_n886));
  INV_X1    g700(.A(new_n851), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n860), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n821), .B1(new_n889), .B2(KEYINPUT54), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT51), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n733), .A2(new_n697), .A3(new_n734), .ZN(new_n892));
  INV_X1    g706(.A(new_n659), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n792), .A2(new_n793), .A3(new_n893), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n892), .A2(new_n800), .A3(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n808), .A2(KEYINPUT115), .A3(new_n809), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n815), .A2(new_n304), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT115), .B1(new_n808), .B2(new_n809), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n896), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n892), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n792), .A2(new_n793), .A3(new_n893), .ZN(new_n905));
  NOR4_X1   g719(.A1(new_n681), .A2(new_n700), .A3(new_n682), .A4(new_n500), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n904), .A2(KEYINPUT50), .A3(new_n905), .A4(new_n906), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n905), .A2(new_n697), .A3(new_n727), .A4(new_n906), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT50), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT116), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n701), .A2(new_n912), .A3(new_n750), .ZN(new_n913));
  OAI21_X1  g727(.A(KEYINPUT116), .B1(new_n800), .B2(new_n700), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n594), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n828), .A2(new_n621), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n819), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n913), .A2(new_n914), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n905), .A2(new_n918), .A3(new_n653), .A4(new_n727), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n911), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n891), .B1(new_n903), .B2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT118), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n808), .A2(new_n809), .A3(new_n899), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n891), .B1(new_n925), .B2(new_n895), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n926), .A2(new_n911), .A3(new_n921), .ZN(new_n927));
  INV_X1    g741(.A(new_n622), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n819), .A2(new_n928), .A3(new_n915), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n700), .A2(new_n501), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n905), .A2(new_n697), .A3(new_n930), .A4(new_n727), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n929), .A2(new_n592), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(KEYINPUT117), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT117), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n929), .A2(new_n931), .A3(new_n934), .A4(new_n592), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n739), .A2(new_n905), .A3(new_n918), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(KEYINPUT48), .ZN(new_n937));
  OR2_X1    g751(.A1(new_n936), .A2(KEYINPUT48), .ZN(new_n938));
  AOI22_X1  g752(.A1(new_n933), .A2(new_n935), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n923), .A2(new_n924), .A3(new_n927), .A4(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n933), .A2(new_n935), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n938), .A2(new_n937), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n941), .A2(new_n927), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n897), .A2(new_n899), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n895), .B1(new_n944), .B2(new_n901), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n920), .B1(new_n910), .B2(new_n907), .ZN(new_n946));
  AOI21_X1  g760(.A(KEYINPUT51), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(KEYINPUT118), .B1(new_n943), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n940), .A2(new_n948), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n882), .A2(new_n890), .A3(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(G952), .A2(G953), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n820), .B1(new_n950), .B2(new_n951), .ZN(G75));
  NAND2_X1  g766(.A1(new_n878), .A2(new_n879), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n953), .A2(G902), .A3(new_n446), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT56), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n495), .A2(new_n496), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n956), .A2(new_n478), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT55), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n954), .A2(new_n955), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n958), .B1(new_n954), .B2(new_n955), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n253), .A2(G952), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(G51));
  XNOR2_X1  g776(.A(new_n307), .B(KEYINPUT57), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n878), .A2(new_n880), .A3(new_n879), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n880), .B1(new_n878), .B2(new_n879), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n966), .B1(new_n375), .B2(new_n377), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n953), .A2(G902), .ZN(new_n968));
  OR2_X1    g782(.A1(new_n968), .A2(new_n776), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n961), .B1(new_n967), .B2(new_n969), .ZN(G54));
  NAND2_X1  g784(.A1(new_n542), .A2(new_n547), .ZN(new_n971));
  NAND2_X1  g785(.A1(KEYINPUT58), .A2(G475), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n971), .B1(new_n968), .B2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n961), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n968), .A2(new_n971), .A3(new_n972), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n975), .A2(new_n976), .ZN(G60));
  XNOR2_X1  g791(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n616), .B(new_n978), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n620), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n964), .B2(new_n965), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n974), .ZN(new_n982));
  INV_X1    g796(.A(new_n979), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n983), .B1(new_n882), .B2(new_n890), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n982), .B1(new_n984), .B2(new_n620), .ZN(G63));
  NAND2_X1  g799(.A1(G217), .A2(G902), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT60), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n953), .A2(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(new_n426), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n961), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n987), .B1(new_n878), .B2(new_n879), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n643), .A2(new_n646), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(KEYINPUT120), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT121), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n991), .B(new_n995), .C1(new_n996), .C2(KEYINPUT61), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT61), .ZN(new_n998));
  OAI211_X1 g812(.A(new_n996), .B(new_n974), .C1(new_n992), .C2(new_n426), .ZN(new_n999));
  INV_X1    g813(.A(new_n995), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n974), .B1(new_n992), .B2(new_n426), .ZN(new_n1001));
  OAI211_X1 g815(.A(new_n998), .B(new_n999), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n997), .A2(new_n1002), .ZN(G66));
  OAI21_X1  g817(.A(G953), .B1(new_n595), .B2(new_n464), .ZN(new_n1004));
  OR2_X1    g818(.A1(new_n859), .A2(new_n838), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1004), .B1(new_n1006), .B2(G953), .ZN(new_n1007));
  INV_X1    g821(.A(G898), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n495), .B1(new_n1008), .B2(G953), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT122), .Z(new_n1010));
  XNOR2_X1  g824(.A(new_n1007), .B(new_n1010), .ZN(G69));
  INV_X1    g825(.A(KEYINPUT124), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n856), .A2(new_n857), .A3(new_n762), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT123), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n759), .A2(KEYINPUT123), .A3(new_n762), .ZN(new_n1016));
  AND2_X1   g830(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n783), .A2(new_n831), .A3(new_n739), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n862), .B1(new_n865), .B2(new_n688), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n804), .A2(new_n1018), .A3(new_n813), .A4(new_n1019), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1012), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1021));
  AND2_X1   g835(.A1(new_n804), .A2(new_n813), .ZN(new_n1022));
  AND2_X1   g836(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1024));
  NAND4_X1  g838(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .A4(KEYINPUT124), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n1021), .A2(new_n1025), .A3(new_n253), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n262), .A2(new_n264), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n507), .A2(new_n508), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1027), .B(new_n1028), .ZN(new_n1029));
  INV_X1    g843(.A(new_n1029), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n1030), .B1(G900), .B2(G953), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1026), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1019), .A2(new_n685), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1033), .A2(KEYINPUT62), .ZN(new_n1034));
  INV_X1    g848(.A(KEYINPUT62), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n1019), .A2(new_n1035), .A3(new_n685), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n835), .A2(new_n622), .ZN(new_n1037));
  NOR2_X1   g851(.A1(new_n678), .A2(new_n800), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n757), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n1034), .A2(new_n1036), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g854(.A(new_n1022), .ZN(new_n1041));
  OAI21_X1  g855(.A(new_n253), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1042), .A2(new_n1030), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1032), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g858(.A1(G227), .A2(G900), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1045), .A2(G953), .ZN(new_n1046));
  AOI21_X1  g860(.A(new_n1046), .B1(new_n1029), .B2(KEYINPUT125), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n1044), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g862(.A(new_n1047), .ZN(new_n1049));
  NAND3_X1  g863(.A1(new_n1032), .A2(new_n1043), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1048), .A2(new_n1050), .ZN(G72));
  NOR3_X1   g865(.A1(new_n1040), .A2(new_n1041), .A3(new_n1005), .ZN(new_n1052));
  NAND2_X1  g866(.A1(G472), .A2(G902), .ZN(new_n1053));
  XNOR2_X1  g867(.A(new_n1053), .B(KEYINPUT63), .ZN(new_n1054));
  XNOR2_X1  g868(.A(new_n1054), .B(KEYINPUT126), .ZN(new_n1055));
  OAI211_X1 g869(.A(new_n257), .B(new_n282), .C1(new_n1052), .C2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g870(.A1(new_n282), .A2(new_n283), .ZN(new_n1057));
  AOI21_X1  g871(.A(new_n1054), .B1(new_n1057), .B2(new_n266), .ZN(new_n1058));
  AOI21_X1  g872(.A(new_n961), .B1(new_n889), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g873(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g874(.A1(new_n1021), .A2(new_n1025), .A3(new_n1006), .ZN(new_n1061));
  INV_X1    g875(.A(new_n1055), .ZN(new_n1062));
  AOI211_X1 g876(.A(new_n257), .B(new_n282), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g877(.A1(new_n1060), .A2(new_n1063), .ZN(G57));
endmodule


