

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X1 U324 ( .A(n549), .B(KEYINPUT36), .ZN(n496) );
  XNOR2_X2 U325 ( .A(n357), .B(KEYINPUT82), .ZN(n388) );
  XNOR2_X2 U326 ( .A(G190GAT), .B(G218GAT), .ZN(n357) );
  XNOR2_X1 U327 ( .A(n400), .B(n399), .ZN(n443) );
  NOR2_X4 U328 ( .A1(n482), .A2(n292), .ZN(n566) );
  XOR2_X2 U329 ( .A(n443), .B(KEYINPUT83), .Z(n549) );
  XNOR2_X1 U330 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n444) );
  XNOR2_X1 U331 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U332 ( .A(n431), .B(n430), .ZN(n433) );
  XNOR2_X1 U333 ( .A(n398), .B(n293), .ZN(n399) );
  XOR2_X1 U334 ( .A(KEYINPUT55), .B(n457), .Z(n292) );
  XOR2_X1 U335 ( .A(n397), .B(n396), .Z(n293) );
  XOR2_X1 U336 ( .A(n425), .B(KEYINPUT33), .Z(n294) );
  INV_X1 U337 ( .A(KEYINPUT117), .ZN(n439) );
  XNOR2_X1 U338 ( .A(n440), .B(n439), .ZN(n441) );
  INV_X1 U339 ( .A(KEYINPUT32), .ZN(n428) );
  NOR2_X1 U340 ( .A1(n541), .A2(n441), .ZN(n442) );
  XNOR2_X1 U341 ( .A(n429), .B(n428), .ZN(n430) );
  INV_X1 U342 ( .A(KEYINPUT86), .ZN(n411) );
  XOR2_X1 U343 ( .A(G71GAT), .B(KEYINPUT13), .Z(n432) );
  XOR2_X1 U344 ( .A(G183GAT), .B(KEYINPUT84), .Z(n403) );
  XNOR2_X1 U345 ( .A(n414), .B(n413), .ZN(n422) );
  XNOR2_X1 U346 ( .A(n577), .B(n444), .ZN(n557) );
  XNOR2_X1 U347 ( .A(n458), .B(G190GAT), .ZN(n459) );
  XNOR2_X1 U348 ( .A(n460), .B(n459), .ZN(G1351GAT) );
  XOR2_X1 U349 ( .A(G176GAT), .B(G183GAT), .Z(n296) );
  XNOR2_X1 U350 ( .A(G169GAT), .B(G15GAT), .ZN(n295) );
  XNOR2_X1 U351 ( .A(n296), .B(n295), .ZN(n304) );
  NAND2_X1 U352 ( .A1(G227GAT), .A2(G233GAT), .ZN(n302) );
  XOR2_X1 U353 ( .A(KEYINPUT90), .B(G120GAT), .Z(n298) );
  XNOR2_X1 U354 ( .A(G134GAT), .B(G99GAT), .ZN(n297) );
  XNOR2_X1 U355 ( .A(n298), .B(n297), .ZN(n300) );
  XOR2_X1 U356 ( .A(G43GAT), .B(G190GAT), .Z(n299) );
  XNOR2_X1 U357 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U358 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U359 ( .A(n304), .B(n303), .ZN(n312) );
  XNOR2_X1 U360 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n305) );
  XNOR2_X1 U361 ( .A(n305), .B(G127GAT), .ZN(n325) );
  XOR2_X1 U362 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n307) );
  XNOR2_X1 U363 ( .A(KEYINPUT20), .B(G71GAT), .ZN(n306) );
  XNOR2_X1 U364 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U365 ( .A(n325), .B(n308), .ZN(n310) );
  XOR2_X1 U366 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n309) );
  XOR2_X1 U367 ( .A(KEYINPUT17), .B(n309), .Z(n350) );
  XOR2_X1 U368 ( .A(n310), .B(n350), .Z(n311) );
  XNOR2_X1 U369 ( .A(n312), .B(n311), .ZN(n482) );
  XOR2_X1 U370 ( .A(KEYINPUT6), .B(KEYINPUT97), .Z(n314) );
  XNOR2_X1 U371 ( .A(KEYINPUT1), .B(KEYINPUT98), .ZN(n313) );
  XNOR2_X1 U372 ( .A(n314), .B(n313), .ZN(n332) );
  XOR2_X1 U373 ( .A(G85GAT), .B(G162GAT), .Z(n316) );
  XNOR2_X1 U374 ( .A(G29GAT), .B(G148GAT), .ZN(n315) );
  XNOR2_X1 U375 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U376 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n318) );
  XNOR2_X1 U377 ( .A(G1GAT), .B(G141GAT), .ZN(n317) );
  XNOR2_X1 U378 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U379 ( .A(n320), .B(n319), .Z(n330) );
  XOR2_X1 U380 ( .A(G155GAT), .B(KEYINPUT2), .Z(n322) );
  XNOR2_X1 U381 ( .A(KEYINPUT3), .B(KEYINPUT94), .ZN(n321) );
  XNOR2_X1 U382 ( .A(n322), .B(n321), .ZN(n347) );
  XOR2_X1 U383 ( .A(n347), .B(KEYINPUT96), .Z(n324) );
  NAND2_X1 U384 ( .A1(G225GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U385 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U386 ( .A(G134GAT), .B(KEYINPUT81), .Z(n392) );
  XNOR2_X1 U387 ( .A(n325), .B(n392), .ZN(n326) );
  XOR2_X1 U388 ( .A(G120GAT), .B(G57GAT), .Z(n427) );
  XNOR2_X1 U389 ( .A(n326), .B(n427), .ZN(n327) );
  XNOR2_X1 U390 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U391 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U392 ( .A(n332), .B(n331), .ZN(n526) );
  INV_X1 U393 ( .A(n526), .ZN(n571) );
  XOR2_X1 U394 ( .A(KEYINPUT93), .B(KEYINPUT95), .Z(n334) );
  XNOR2_X1 U395 ( .A(G106GAT), .B(KEYINPUT24), .ZN(n333) );
  XNOR2_X1 U396 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U397 ( .A(KEYINPUT79), .B(G162GAT), .Z(n393) );
  XOR2_X1 U398 ( .A(G218GAT), .B(n393), .Z(n336) );
  XOR2_X1 U399 ( .A(G141GAT), .B(G22GAT), .Z(n380) );
  XNOR2_X1 U400 ( .A(G50GAT), .B(n380), .ZN(n335) );
  XNOR2_X1 U401 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U402 ( .A(n338), .B(n337), .Z(n340) );
  NAND2_X1 U403 ( .A1(G228GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U404 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U405 ( .A(n341), .B(KEYINPUT23), .Z(n344) );
  XNOR2_X1 U406 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n342) );
  XNOR2_X1 U407 ( .A(n342), .B(G211GAT), .ZN(n358) );
  XNOR2_X1 U408 ( .A(n358), .B(KEYINPUT22), .ZN(n343) );
  XNOR2_X1 U409 ( .A(n344), .B(n343), .ZN(n349) );
  XOR2_X1 U410 ( .A(G78GAT), .B(G148GAT), .Z(n346) );
  XNOR2_X1 U411 ( .A(KEYINPUT77), .B(G204GAT), .ZN(n345) );
  XNOR2_X1 U412 ( .A(n346), .B(n345), .ZN(n435) );
  XOR2_X1 U413 ( .A(n435), .B(n347), .Z(n348) );
  XNOR2_X1 U414 ( .A(n349), .B(n348), .ZN(n481) );
  AND2_X1 U415 ( .A1(n571), .A2(n481), .ZN(n454) );
  XOR2_X1 U416 ( .A(G176GAT), .B(G64GAT), .Z(n434) );
  XNOR2_X1 U417 ( .A(n434), .B(n403), .ZN(n362) );
  XOR2_X1 U418 ( .A(G169GAT), .B(G8GAT), .Z(n374) );
  XOR2_X1 U419 ( .A(n350), .B(n374), .Z(n352) );
  NAND2_X1 U420 ( .A1(G226GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U421 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U422 ( .A(KEYINPUT99), .B(G92GAT), .Z(n354) );
  XNOR2_X1 U423 ( .A(G36GAT), .B(G204GAT), .ZN(n353) );
  XNOR2_X1 U424 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U425 ( .A(n356), .B(n355), .Z(n360) );
  XNOR2_X1 U426 ( .A(n358), .B(n388), .ZN(n359) );
  XNOR2_X1 U427 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U428 ( .A(n362), .B(n361), .ZN(n472) );
  XOR2_X1 U429 ( .A(G29GAT), .B(G36GAT), .Z(n364) );
  XNOR2_X1 U430 ( .A(G50GAT), .B(G43GAT), .ZN(n363) );
  XNOR2_X1 U431 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U432 ( .A(KEYINPUT7), .B(KEYINPUT71), .Z(n366) );
  XNOR2_X1 U433 ( .A(KEYINPUT72), .B(KEYINPUT8), .ZN(n365) );
  XNOR2_X1 U434 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U435 ( .A(n368), .B(n367), .Z(n398) );
  XOR2_X1 U436 ( .A(KEYINPUT75), .B(KEYINPUT29), .Z(n370) );
  XNOR2_X1 U437 ( .A(KEYINPUT69), .B(KEYINPUT68), .ZN(n369) );
  XNOR2_X1 U438 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U439 ( .A(n398), .B(n371), .ZN(n385) );
  XOR2_X1 U440 ( .A(KEYINPUT70), .B(KEYINPUT67), .Z(n373) );
  XNOR2_X1 U441 ( .A(G197GAT), .B(G113GAT), .ZN(n372) );
  XNOR2_X1 U442 ( .A(n373), .B(n372), .ZN(n375) );
  XOR2_X1 U443 ( .A(n375), .B(n374), .Z(n383) );
  XOR2_X1 U444 ( .A(G1GAT), .B(KEYINPUT73), .Z(n377) );
  XNOR2_X1 U445 ( .A(G15GAT), .B(KEYINPUT74), .ZN(n376) );
  XNOR2_X1 U446 ( .A(n377), .B(n376), .ZN(n410) );
  XOR2_X1 U447 ( .A(n410), .B(KEYINPUT30), .Z(n379) );
  NAND2_X1 U448 ( .A1(G229GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U449 ( .A(n379), .B(n378), .ZN(n381) );
  XNOR2_X1 U450 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U451 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U452 ( .A(n385), .B(n384), .ZN(n574) );
  XNOR2_X1 U453 ( .A(n574), .B(KEYINPUT76), .ZN(n541) );
  XOR2_X1 U454 ( .A(G92GAT), .B(G85GAT), .Z(n387) );
  XNOR2_X1 U455 ( .A(G99GAT), .B(G106GAT), .ZN(n386) );
  XNOR2_X1 U456 ( .A(n387), .B(n386), .ZN(n425) );
  XNOR2_X1 U457 ( .A(n388), .B(KEYINPUT65), .ZN(n390) );
  AND2_X1 U458 ( .A1(G232GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U459 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U460 ( .A(n425), .B(n391), .ZN(n395) );
  XOR2_X1 U461 ( .A(n393), .B(n392), .Z(n394) );
  XNOR2_X1 U462 ( .A(n395), .B(n394), .ZN(n400) );
  XOR2_X1 U463 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n397) );
  XNOR2_X1 U464 ( .A(KEYINPUT11), .B(KEYINPUT80), .ZN(n396) );
  XOR2_X1 U465 ( .A(KEYINPUT88), .B(KEYINPUT14), .Z(n402) );
  XNOR2_X1 U466 ( .A(KEYINPUT89), .B(KEYINPUT12), .ZN(n401) );
  XNOR2_X1 U467 ( .A(n402), .B(n401), .ZN(n407) );
  XOR2_X1 U468 ( .A(n432), .B(n403), .Z(n405) );
  XNOR2_X1 U469 ( .A(G78GAT), .B(G211GAT), .ZN(n404) );
  XNOR2_X1 U470 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U471 ( .A(n407), .B(n406), .Z(n409) );
  NAND2_X1 U472 ( .A1(G231GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U473 ( .A(n409), .B(n408), .ZN(n414) );
  XNOR2_X1 U474 ( .A(n410), .B(KEYINPUT87), .ZN(n412) );
  XOR2_X1 U475 ( .A(KEYINPUT85), .B(KEYINPUT15), .Z(n416) );
  XNOR2_X1 U476 ( .A(G57GAT), .B(G64GAT), .ZN(n415) );
  XNOR2_X1 U477 ( .A(n416), .B(n415), .ZN(n420) );
  XOR2_X1 U478 ( .A(G155GAT), .B(G127GAT), .Z(n418) );
  XNOR2_X1 U479 ( .A(G22GAT), .B(G8GAT), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U481 ( .A(n420), .B(n419), .Z(n421) );
  XNOR2_X1 U482 ( .A(n422), .B(n421), .ZN(n467) );
  INV_X1 U483 ( .A(n467), .ZN(n581) );
  NAND2_X1 U484 ( .A1(n496), .A2(n581), .ZN(n424) );
  XOR2_X1 U485 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n423) );
  XNOR2_X1 U486 ( .A(n424), .B(n423), .ZN(n438) );
  NAND2_X1 U487 ( .A1(G230GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U488 ( .A(n294), .B(n426), .ZN(n431) );
  XNOR2_X1 U489 ( .A(n427), .B(KEYINPUT31), .ZN(n429) );
  XOR2_X1 U490 ( .A(n433), .B(n432), .Z(n437) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n577) );
  NAND2_X1 U493 ( .A1(n438), .A2(n577), .ZN(n440) );
  XNOR2_X1 U494 ( .A(n442), .B(KEYINPUT118), .ZN(n451) );
  NAND2_X1 U495 ( .A1(n557), .A2(n574), .ZN(n446) );
  XNOR2_X1 U496 ( .A(KEYINPUT116), .B(KEYINPUT46), .ZN(n445) );
  XNOR2_X1 U497 ( .A(n446), .B(n445), .ZN(n447) );
  NAND2_X1 U498 ( .A1(n447), .A2(n467), .ZN(n448) );
  NOR2_X1 U499 ( .A1(n443), .A2(n448), .ZN(n449) );
  XOR2_X1 U500 ( .A(KEYINPUT47), .B(n449), .Z(n450) );
  NOR2_X1 U501 ( .A1(n451), .A2(n450), .ZN(n452) );
  XNOR2_X1 U502 ( .A(KEYINPUT48), .B(n452), .ZN(n537) );
  NOR2_X1 U503 ( .A1(n472), .A2(n537), .ZN(n453) );
  XNOR2_X1 U504 ( .A(KEYINPUT54), .B(n453), .ZN(n570) );
  NAND2_X1 U505 ( .A1(n454), .A2(n570), .ZN(n456) );
  XOR2_X1 U506 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n455) );
  XNOR2_X1 U507 ( .A(n456), .B(n455), .ZN(n457) );
  NAND2_X1 U508 ( .A1(n566), .A2(n549), .ZN(n460) );
  XOR2_X1 U509 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n458) );
  NAND2_X1 U510 ( .A1(n541), .A2(n566), .ZN(n462) );
  XNOR2_X1 U511 ( .A(G169GAT), .B(KEYINPUT124), .ZN(n461) );
  XNOR2_X1 U512 ( .A(n462), .B(n461), .ZN(G1348GAT) );
  XNOR2_X1 U513 ( .A(n557), .B(KEYINPUT108), .ZN(n543) );
  NAND2_X1 U514 ( .A1(n566), .A2(n543), .ZN(n465) );
  XOR2_X1 U515 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n463) );
  XNOR2_X1 U516 ( .A(n463), .B(G176GAT), .ZN(n464) );
  XNOR2_X1 U517 ( .A(n465), .B(n464), .ZN(G1349GAT) );
  XOR2_X1 U518 ( .A(KEYINPUT34), .B(KEYINPUT105), .Z(n488) );
  NAND2_X1 U519 ( .A1(n541), .A2(n577), .ZN(n466) );
  XNOR2_X1 U520 ( .A(n466), .B(KEYINPUT78), .ZN(n501) );
  NOR2_X1 U521 ( .A1(n467), .A2(n549), .ZN(n468) );
  XNOR2_X1 U522 ( .A(KEYINPUT16), .B(n468), .ZN(n485) );
  INV_X1 U523 ( .A(n482), .ZN(n538) );
  INV_X1 U524 ( .A(n472), .ZN(n528) );
  NAND2_X1 U525 ( .A1(n538), .A2(n528), .ZN(n469) );
  NAND2_X1 U526 ( .A1(n469), .A2(n481), .ZN(n470) );
  XNOR2_X1 U527 ( .A(n470), .B(KEYINPUT102), .ZN(n471) );
  XOR2_X1 U528 ( .A(KEYINPUT25), .B(n471), .Z(n476) );
  XOR2_X1 U529 ( .A(n472), .B(KEYINPUT27), .Z(n479) );
  NOR2_X1 U530 ( .A1(n538), .A2(n481), .ZN(n474) );
  XNOR2_X1 U531 ( .A(KEYINPUT101), .B(KEYINPUT26), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n474), .B(n473), .ZN(n555) );
  INV_X1 U533 ( .A(n555), .ZN(n573) );
  NAND2_X1 U534 ( .A1(n479), .A2(n573), .ZN(n475) );
  NAND2_X1 U535 ( .A1(n476), .A2(n475), .ZN(n477) );
  NAND2_X1 U536 ( .A1(n571), .A2(n477), .ZN(n478) );
  XOR2_X1 U537 ( .A(KEYINPUT103), .B(n478), .Z(n484) );
  NAND2_X1 U538 ( .A1(n526), .A2(n479), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n480), .B(KEYINPUT100), .ZN(n553) );
  XOR2_X1 U540 ( .A(KEYINPUT28), .B(n481), .Z(n532) );
  NOR2_X1 U541 ( .A1(n553), .A2(n532), .ZN(n539) );
  NAND2_X1 U542 ( .A1(n482), .A2(n539), .ZN(n483) );
  NAND2_X1 U543 ( .A1(n484), .A2(n483), .ZN(n497) );
  NAND2_X1 U544 ( .A1(n485), .A2(n497), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n486), .B(KEYINPUT104), .ZN(n511) );
  NOR2_X1 U546 ( .A1(n501), .A2(n511), .ZN(n494) );
  NAND2_X1 U547 ( .A1(n494), .A2(n526), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U549 ( .A(G1GAT), .B(n489), .ZN(G1324GAT) );
  NAND2_X1 U550 ( .A1(n528), .A2(n494), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n490), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U552 ( .A(KEYINPUT35), .B(KEYINPUT106), .Z(n492) );
  NAND2_X1 U553 ( .A1(n494), .A2(n538), .ZN(n491) );
  XNOR2_X1 U554 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U555 ( .A(G15GAT), .B(n493), .ZN(G1326GAT) );
  NAND2_X1 U556 ( .A1(n532), .A2(n494), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n495), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U558 ( .A(G29GAT), .B(KEYINPUT39), .Z(n504) );
  NAND2_X1 U559 ( .A1(n496), .A2(n497), .ZN(n498) );
  NOR2_X1 U560 ( .A1(n581), .A2(n498), .ZN(n500) );
  XOR2_X1 U561 ( .A(KEYINPUT107), .B(KEYINPUT37), .Z(n499) );
  XNOR2_X1 U562 ( .A(n500), .B(n499), .ZN(n525) );
  NOR2_X1 U563 ( .A1(n525), .A2(n501), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n502), .B(KEYINPUT38), .ZN(n508) );
  NAND2_X1 U565 ( .A1(n508), .A2(n526), .ZN(n503) );
  XNOR2_X1 U566 ( .A(n504), .B(n503), .ZN(G1328GAT) );
  NAND2_X1 U567 ( .A1(n508), .A2(n528), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n505), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U569 ( .A1(n508), .A2(n538), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n506), .B(KEYINPUT40), .ZN(n507) );
  XNOR2_X1 U571 ( .A(G43GAT), .B(n507), .ZN(G1330GAT) );
  NAND2_X1 U572 ( .A1(n508), .A2(n532), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n509), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n513) );
  INV_X1 U575 ( .A(n574), .ZN(n510) );
  NAND2_X1 U576 ( .A1(n510), .A2(n543), .ZN(n524) );
  NOR2_X1 U577 ( .A1(n511), .A2(n524), .ZN(n519) );
  NAND2_X1 U578 ( .A1(n519), .A2(n526), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U580 ( .A(G57GAT), .B(n514), .ZN(G1332GAT) );
  NAND2_X1 U581 ( .A1(n528), .A2(n519), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n515), .B(KEYINPUT110), .ZN(n516) );
  XNOR2_X1 U583 ( .A(G64GAT), .B(n516), .ZN(G1333GAT) );
  XOR2_X1 U584 ( .A(G71GAT), .B(KEYINPUT111), .Z(n518) );
  NAND2_X1 U585 ( .A1(n519), .A2(n538), .ZN(n517) );
  XNOR2_X1 U586 ( .A(n518), .B(n517), .ZN(G1334GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT113), .B(KEYINPUT43), .Z(n521) );
  NAND2_X1 U588 ( .A1(n519), .A2(n532), .ZN(n520) );
  XNOR2_X1 U589 ( .A(n521), .B(n520), .ZN(n523) );
  XOR2_X1 U590 ( .A(G78GAT), .B(KEYINPUT112), .Z(n522) );
  XNOR2_X1 U591 ( .A(n523), .B(n522), .ZN(G1335GAT) );
  NOR2_X1 U592 ( .A1(n525), .A2(n524), .ZN(n533) );
  NAND2_X1 U593 ( .A1(n533), .A2(n526), .ZN(n527) );
  XNOR2_X1 U594 ( .A(G85GAT), .B(n527), .ZN(G1336GAT) );
  NAND2_X1 U595 ( .A1(n528), .A2(n533), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n529), .B(KEYINPUT114), .ZN(n530) );
  XNOR2_X1 U597 ( .A(G92GAT), .B(n530), .ZN(G1337GAT) );
  NAND2_X1 U598 ( .A1(n538), .A2(n533), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n531), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT44), .B(KEYINPUT115), .Z(n535) );
  NAND2_X1 U601 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U603 ( .A(G106GAT), .B(n536), .ZN(G1339GAT) );
  NAND2_X1 U604 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U605 ( .A1(n537), .A2(n540), .ZN(n550) );
  NAND2_X1 U606 ( .A1(n541), .A2(n550), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n542), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT119), .B(KEYINPUT49), .Z(n545) );
  NAND2_X1 U609 ( .A1(n550), .A2(n543), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U611 ( .A(G120GAT), .B(n546), .Z(G1341GAT) );
  NAND2_X1 U612 ( .A1(n550), .A2(n581), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n547), .B(KEYINPUT50), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G127GAT), .B(n548), .ZN(G1342GAT) );
  XOR2_X1 U615 ( .A(G134GAT), .B(KEYINPUT51), .Z(n552) );
  NAND2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(G1343GAT) );
  OR2_X1 U618 ( .A1(n537), .A2(n553), .ZN(n554) );
  NOR2_X1 U619 ( .A1(n555), .A2(n554), .ZN(n563) );
  NAND2_X1 U620 ( .A1(n574), .A2(n563), .ZN(n556) );
  XNOR2_X1 U621 ( .A(G141GAT), .B(n556), .ZN(G1344GAT) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n561) );
  XOR2_X1 U623 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n559) );
  NAND2_X1 U624 ( .A1(n563), .A2(n557), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(G1345GAT) );
  NAND2_X1 U627 ( .A1(n563), .A2(n581), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U629 ( .A(G162GAT), .B(KEYINPUT121), .Z(n565) );
  NAND2_X1 U630 ( .A1(n563), .A2(n443), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1347GAT) );
  NAND2_X1 U632 ( .A1(n566), .A2(n581), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n568), .B(KEYINPUT60), .ZN(n569) );
  XOR2_X1 U636 ( .A(KEYINPUT126), .B(n569), .Z(n576) );
  AND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  AND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n583) );
  NAND2_X1 U639 ( .A1(n583), .A2(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT61), .Z(n580) );
  INV_X1 U642 ( .A(n577), .ZN(n578) );
  NAND2_X1 U643 ( .A1(n583), .A2(n578), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  NAND2_X1 U645 ( .A1(n583), .A2(n581), .ZN(n582) );
  XNOR2_X1 U646 ( .A(n582), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n585) );
  NAND2_X1 U648 ( .A1(n583), .A2(n496), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

