//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 1 0 0 0 1 1 1 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0 0 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1289, new_n1290, new_n1291,
    new_n1292, new_n1293, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1344, new_n1345, new_n1346;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n206), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  OR2_X1    g0019(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n220));
  NOR2_X1   g0020(.A1(G58), .A2(G68), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n221), .A2(KEYINPUT64), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(KEYINPUT64), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n222), .A2(G50), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G20), .ZN(new_n227));
  OR2_X1    g0027(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n209), .A2(new_n220), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n219), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G68), .Z(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  NAND3_X1  g0045(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(new_n225), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n213), .A2(KEYINPUT15), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT15), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G87), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n204), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT8), .B(G58), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n204), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G77), .ZN(new_n258));
  OAI22_X1  g0058(.A1(new_n255), .A2(new_n257), .B1(new_n204), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n247), .B1(new_n254), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n260), .B(KEYINPUT66), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n262));
  AND3_X1   g0062(.A1(new_n262), .A2(new_n225), .A3(new_n246), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n258), .B1(new_n203), .B2(G20), .ZN(new_n264));
  INV_X1    g0064(.A(new_n262), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n263), .A2(new_n264), .B1(new_n258), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n226), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G274), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n274), .B1(new_n226), .B2(new_n269), .ZN(new_n275));
  INV_X1    g0075(.A(new_n271), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n273), .A2(G244), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  OR2_X1    g0077(.A1(new_n277), .A2(KEYINPUT65), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n225), .B1(G33), .B2(G41), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT3), .B(G33), .ZN(new_n280));
  INV_X1    g0080(.A(G1698), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(G232), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G107), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n282), .B1(new_n283), .B2(new_n280), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT3), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NOR3_X1   g0088(.A1(new_n288), .A2(new_n212), .A3(new_n281), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n279), .B1(new_n284), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n277), .A2(KEYINPUT65), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n278), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT67), .B(G200), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G190), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n268), .B(new_n294), .C1(new_n295), .C2(new_n292), .ZN(new_n296));
  INV_X1    g0096(.A(G169), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n298), .B(new_n267), .C1(G179), .C2(new_n292), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G150), .ZN(new_n301));
  OAI22_X1  g0101(.A1(new_n255), .A2(new_n253), .B1(new_n301), .B2(new_n257), .ZN(new_n302));
  INV_X1    g0102(.A(G50), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n204), .B1(new_n221), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n247), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n303), .B1(new_n203), .B2(G20), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n263), .A2(new_n306), .B1(new_n303), .B2(new_n265), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(G222), .A2(G1698), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n281), .A2(G223), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n280), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n311), .B(new_n279), .C1(G77), .C2(new_n280), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n275), .A2(new_n276), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n273), .A2(G226), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n308), .B1(new_n297), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n316), .B1(G179), .B2(new_n315), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n308), .A2(KEYINPUT9), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n318), .B(KEYINPUT68), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n308), .A2(KEYINPUT9), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n315), .A2(new_n293), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n315), .A2(new_n295), .ZN(new_n322));
  NOR3_X1   g0122(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT10), .ZN(new_n324));
  AND3_X1   g0124(.A1(new_n319), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n324), .B1(new_n319), .B2(new_n323), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n300), .B(new_n317), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n255), .B1(new_n203), .B2(G20), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n328), .A2(new_n263), .B1(new_n265), .B2(new_n255), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n247), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT74), .ZN(new_n332));
  INV_X1    g0132(.A(G159), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n332), .B1(new_n257), .B2(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(G20), .A2(G33), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n335), .A2(KEYINPUT74), .A3(G159), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g0137(.A(G58), .B(G68), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(G20), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT73), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n288), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n280), .A2(KEYINPUT73), .ZN(new_n343));
  NOR2_X1   g0143(.A1(KEYINPUT7), .A2(G20), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n288), .A2(new_n204), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n211), .B1(new_n346), .B2(KEYINPUT7), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n340), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n331), .B1(new_n348), .B2(KEYINPUT16), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT16), .ZN(new_n350));
  OAI21_X1  g0150(.A(KEYINPUT75), .B1(new_n256), .B2(KEYINPUT3), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT75), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n352), .A2(new_n285), .A3(G33), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n351), .A2(new_n353), .A3(new_n287), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT7), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n355), .A2(G20), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n355), .B1(new_n280), .B2(G20), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n211), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n350), .B1(new_n359), .B2(new_n340), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n330), .B1(new_n349), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G232), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n313), .B1(new_n362), .B2(new_n272), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  OR2_X1    g0164(.A1(G223), .A2(G1698), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n281), .A2(G226), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n280), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(G33), .A2(G87), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n270), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n297), .B1(new_n364), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G179), .ZN(new_n372));
  NOR3_X1   g0172(.A1(new_n363), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(KEYINPUT18), .B1(new_n361), .B2(new_n374), .ZN(new_n375));
  XOR2_X1   g0175(.A(KEYINPUT76), .B(G190), .Z(new_n376));
  NAND3_X1  g0176(.A1(new_n364), .A2(new_n370), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G200), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(new_n363), .B2(new_n369), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n361), .A2(KEYINPUT17), .A3(new_n380), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n337), .A2(new_n339), .ZN(new_n382));
  INV_X1    g0182(.A(new_n345), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n280), .A2(G20), .ZN(new_n384));
  OAI21_X1  g0184(.A(G68), .B1(new_n384), .B2(new_n355), .ZN(new_n385));
  OAI211_X1 g0185(.A(KEYINPUT16), .B(new_n382), .C1(new_n383), .C2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n386), .A2(new_n360), .A3(new_n247), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n329), .ZN(new_n388));
  INV_X1    g0188(.A(new_n374), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT18), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n387), .A2(new_n329), .A3(new_n380), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT17), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n375), .A2(new_n381), .A3(new_n391), .A4(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n327), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n263), .B(G68), .C1(G1), .C2(new_n204), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT12), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n398), .B1(new_n265), .B2(new_n211), .ZN(new_n399));
  NOR3_X1   g0199(.A1(new_n262), .A2(KEYINPUT12), .A3(G68), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n397), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI22_X1  g0201(.A1(new_n253), .A2(new_n258), .B1(new_n204), .B2(G68), .ZN(new_n402));
  OAI22_X1  g0202(.A1(new_n402), .A2(KEYINPUT70), .B1(new_n303), .B2(new_n257), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n402), .A2(KEYINPUT70), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n247), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT71), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT71), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n407), .B(new_n247), .C1(new_n403), .C2(new_n404), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n401), .B1(new_n409), .B2(KEYINPUT11), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(KEYINPUT11), .B2(new_n409), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n286), .A2(new_n287), .A3(G232), .A4(G1698), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT69), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT69), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n280), .A2(new_n414), .A3(G232), .A4(G1698), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n286), .A2(new_n287), .A3(G226), .A4(new_n281), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G33), .A2(G97), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n270), .B1(new_n416), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n313), .B1(new_n272), .B2(new_n212), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT13), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n422), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT13), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n419), .B1(new_n415), .B2(new_n413), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n424), .B(new_n425), .C1(new_n426), .C2(new_n270), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n423), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(new_n295), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n378), .B1(new_n423), .B2(new_n427), .ZN(new_n430));
  NOR3_X1   g0230(.A1(new_n411), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT72), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n428), .A2(G169), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n432), .B1(new_n433), .B2(KEYINPUT14), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(KEYINPUT14), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT14), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n428), .A2(KEYINPUT72), .A3(new_n436), .A4(G169), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n423), .A2(new_n427), .A3(G179), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n434), .A2(new_n435), .A3(new_n437), .A4(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n431), .B1(new_n439), .B2(new_n411), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n396), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n212), .A2(new_n281), .ZN(new_n443));
  INV_X1    g0243(.A(G244), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(G1698), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n286), .A2(new_n443), .A3(new_n287), .A4(new_n445), .ZN(new_n446));
  AND2_X1   g0246(.A1(G33), .A2(G116), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n446), .A2(KEYINPUT79), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT79), .B1(new_n446), .B2(new_n448), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n279), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(G45), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(G1), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n275), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n203), .A2(G45), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n270), .A2(G250), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  AND3_X1   g0258(.A1(new_n451), .A2(new_n372), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(G169), .B1(new_n451), .B2(new_n458), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT80), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT19), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n204), .B1(new_n418), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G97), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n213), .A2(new_n465), .A3(new_n283), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n286), .A2(new_n287), .A3(new_n204), .A4(G68), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n463), .B1(new_n253), .B2(new_n465), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n247), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n251), .A2(new_n262), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n462), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  AOI211_X1 g0274(.A(KEYINPUT80), .B(new_n472), .C1(new_n470), .C2(new_n247), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n203), .A2(G33), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n262), .A2(new_n476), .A3(new_n225), .A4(new_n246), .ZN(new_n477));
  OAI22_X1  g0277(.A1(new_n474), .A2(new_n475), .B1(new_n477), .B2(new_n252), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n451), .A2(new_n295), .A3(new_n458), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n446), .A2(new_n448), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT79), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n446), .A2(KEYINPUT79), .A3(new_n448), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n457), .B1(new_n484), .B2(new_n279), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n479), .B1(new_n485), .B2(new_n293), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n477), .A2(new_n213), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n471), .A2(new_n473), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT80), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n471), .A2(new_n462), .A3(new_n473), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n487), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n461), .A2(new_n478), .B1(new_n486), .B2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n286), .A2(new_n287), .A3(G244), .A4(new_n281), .ZN(new_n493));
  XOR2_X1   g0293(.A(KEYINPUT77), .B(KEYINPUT4), .Z(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G250), .A2(G1698), .ZN(new_n496));
  NAND2_X1  g0296(.A1(KEYINPUT4), .A2(G244), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n496), .B1(new_n497), .B2(G1698), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n280), .A2(new_n498), .B1(G33), .B2(G283), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n279), .ZN(new_n501));
  NAND2_X1  g0301(.A1(KEYINPUT5), .A2(G41), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(KEYINPUT5), .A2(G41), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n453), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(G257), .A3(new_n270), .ZN(new_n506));
  OR2_X1    g0306(.A1(KEYINPUT5), .A2(G41), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n455), .B1(new_n507), .B2(new_n502), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n275), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n501), .A2(G179), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n270), .B1(new_n495), .B2(new_n499), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n506), .A2(new_n509), .ZN(new_n513));
  OAI21_X1  g0313(.A(G169), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n283), .B1(new_n357), .B2(new_n358), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n335), .A2(G77), .ZN(new_n517));
  AND3_X1   g0317(.A1(new_n283), .A2(KEYINPUT6), .A3(G97), .ZN(new_n518));
  XNOR2_X1  g0318(.A(G97), .B(G107), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT6), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n517), .B1(new_n521), .B2(new_n204), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n247), .B1(new_n516), .B2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT78), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n265), .A2(new_n465), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n477), .B2(new_n465), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  AND3_X1   g0327(.A1(new_n523), .A2(new_n524), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n524), .B1(new_n523), .B2(new_n527), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n515), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n519), .A2(new_n520), .ZN(new_n531));
  INV_X1    g0331(.A(new_n518), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(G20), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n346), .A2(new_n355), .B1(new_n354), .B2(new_n356), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n534), .B(new_n517), .C1(new_n535), .C2(new_n283), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n526), .B1(new_n536), .B2(new_n247), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n501), .A2(new_n510), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G200), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n537), .B(new_n539), .C1(new_n295), .C2(new_n538), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT25), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n262), .B2(G107), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n262), .A2(new_n541), .A3(G107), .ZN(new_n544));
  OAI22_X1  g0344(.A1(new_n543), .A2(new_n544), .B1(new_n283), .B2(new_n477), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT23), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n204), .B2(G107), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n283), .A2(KEYINPUT23), .A3(G20), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n547), .A2(new_n548), .B1(new_n204), .B2(new_n447), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT22), .ZN(new_n550));
  OAI21_X1  g0350(.A(KEYINPUT86), .B1(new_n550), .B2(KEYINPUT85), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(KEYINPUT86), .B2(new_n550), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n286), .A2(new_n287), .A3(new_n204), .A4(G87), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n549), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT86), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT85), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n555), .B1(new_n556), .B2(KEYINPUT22), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(KEYINPUT24), .B1(new_n554), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n550), .A2(KEYINPUT86), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n561), .A2(new_n204), .A3(G87), .A4(new_n280), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT24), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n553), .A2(new_n557), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .A4(new_n549), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n559), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n545), .B1(new_n566), .B2(new_n247), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n286), .A2(new_n287), .A3(G257), .A4(G1698), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n286), .A2(new_n287), .A3(G250), .A4(new_n281), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G33), .A2(G294), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n279), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n505), .A2(G264), .A3(new_n270), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n572), .A2(new_n509), .A3(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n574), .A2(G190), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT87), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n505), .A2(KEYINPUT87), .A3(G264), .A4(new_n270), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n577), .A2(new_n578), .B1(new_n279), .B2(new_n571), .ZN(new_n579));
  AOI21_X1  g0379(.A(G200), .B1(new_n579), .B2(new_n509), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n567), .B1(new_n575), .B2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n492), .A2(new_n530), .A3(new_n540), .A4(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT88), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n577), .A2(new_n578), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n584), .A2(G179), .A3(new_n509), .A4(new_n572), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n574), .A2(G169), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n583), .B1(new_n587), .B2(new_n567), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n566), .A2(new_n247), .ZN(new_n589));
  INV_X1    g0389(.A(new_n545), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n585), .A2(new_n586), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(KEYINPUT88), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n507), .A2(new_n502), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n279), .B1(new_n453), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n596), .A2(G270), .B1(new_n275), .B2(new_n508), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n286), .A2(new_n287), .A3(G264), .A4(G1698), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n286), .A2(new_n287), .A3(G257), .A4(new_n281), .ZN(new_n599));
  INV_X1    g0399(.A(G303), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n598), .B(new_n599), .C1(new_n600), .C2(new_n280), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n279), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n297), .B1(new_n597), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT81), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n263), .A2(new_n604), .A3(G116), .A4(new_n476), .ZN(new_n605));
  INV_X1    g0405(.A(G116), .ZN(new_n606));
  OAI21_X1  g0406(.A(KEYINPUT81), .B1(new_n477), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n246), .A2(new_n225), .B1(G20), .B2(new_n606), .ZN(new_n609));
  NAND2_X1  g0409(.A1(G33), .A2(G283), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n610), .B(new_n204), .C1(G33), .C2(new_n465), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT20), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n609), .A2(KEYINPUT20), .A3(new_n611), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n203), .A2(new_n606), .A3(G13), .A4(G20), .ZN(new_n617));
  XNOR2_X1  g0417(.A(new_n617), .B(KEYINPUT82), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n608), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(KEYINPUT21), .B1(new_n603), .B2(new_n619), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n608), .A2(new_n616), .A3(new_n618), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n597), .A2(new_n602), .A3(G179), .ZN(new_n622));
  OAI21_X1  g0422(.A(KEYINPUT84), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n597), .A2(new_n602), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT84), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n625), .A2(new_n619), .A3(new_n626), .A4(G179), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n620), .B1(new_n623), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n603), .A2(new_n619), .A3(KEYINPUT21), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT83), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n603), .A2(new_n619), .A3(KEYINPUT83), .A4(KEYINPUT21), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n619), .B1(G200), .B2(new_n624), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n624), .B2(new_n376), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n628), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  NOR3_X1   g0436(.A1(new_n582), .A2(new_n594), .A3(new_n636), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n442), .A2(new_n637), .ZN(G372));
  AND2_X1   g0438(.A1(new_n375), .A2(new_n391), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n439), .A2(new_n411), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n640), .A2(new_n299), .ZN(new_n641));
  INV_X1    g0441(.A(new_n431), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n642), .A2(new_n394), .A3(new_n381), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n639), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n325), .A2(new_n326), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n317), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n451), .A2(new_n458), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n297), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n451), .A2(new_n372), .A3(new_n458), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n478), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n297), .B1(new_n501), .B2(new_n510), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n512), .A2(new_n513), .A3(new_n372), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(KEYINPUT90), .B1(new_n655), .B2(new_n537), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n486), .A2(new_n491), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT90), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n523), .A2(new_n527), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n515), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n656), .A2(new_n657), .A3(new_n652), .A4(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n652), .B1(new_n661), .B2(KEYINPUT26), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT26), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n659), .A2(KEYINPUT78), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n523), .A2(new_n524), .A3(new_n527), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n655), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n663), .B1(new_n492), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(KEYINPUT91), .B1(new_n662), .B2(new_n667), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n515), .A2(new_n658), .A3(new_n659), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n658), .B1(new_n515), .B2(new_n659), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n671), .A2(new_n663), .A3(new_n492), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n657), .A2(new_n652), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT26), .B1(new_n673), .B2(new_n530), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT91), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n672), .A2(new_n674), .A3(new_n675), .A4(new_n652), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n581), .A2(new_n657), .A3(new_n652), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n530), .A2(new_n540), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n591), .A2(new_n592), .ZN(new_n680));
  AND3_X1   g0480(.A1(new_n628), .A2(new_n633), .A3(KEYINPUT89), .ZN(new_n681));
  AOI21_X1  g0481(.A(KEYINPUT89), .B1(new_n628), .B2(new_n633), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n680), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AOI22_X1  g0483(.A1(new_n668), .A2(new_n676), .B1(new_n679), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n648), .B1(new_n441), .B2(new_n684), .ZN(G369));
  NOR2_X1   g0485(.A1(new_n681), .A2(new_n682), .ZN(new_n686));
  INV_X1    g0486(.A(G13), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n687), .A2(G1), .A3(G20), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(G213), .B1(new_n689), .B2(KEYINPUT27), .ZN(new_n690));
  AOI21_X1  g0490(.A(KEYINPUT92), .B1(new_n689), .B2(KEYINPUT27), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n689), .A2(KEYINPUT92), .A3(KEYINPUT27), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n690), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(G343), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(new_n621), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n686), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n636), .B2(new_n699), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(G330), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n594), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n704), .A2(new_n581), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n567), .B2(new_n698), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n680), .B2(new_n698), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n680), .A2(new_n697), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n697), .B1(new_n628), .B2(new_n633), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n709), .B1(new_n705), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n708), .A2(new_n711), .ZN(G399));
  INV_X1    g0512(.A(new_n207), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G41), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n466), .A2(G116), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n715), .A2(G1), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(new_n224), .B2(new_n715), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT28), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n668), .A2(new_n676), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n683), .A2(new_n679), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT29), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n722), .A2(new_n723), .A3(new_n698), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT96), .ZN(new_n725));
  AND4_X1   g0525(.A1(new_n588), .A2(new_n628), .A3(new_n593), .A4(new_n633), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n725), .B1(new_n726), .B2(new_n582), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n666), .A2(new_n663), .A3(new_n652), .A4(new_n657), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(new_n652), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n663), .B1(new_n671), .B2(new_n492), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n588), .A2(new_n628), .A3(new_n593), .A4(new_n633), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n679), .A2(KEYINPUT96), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n727), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n698), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(KEYINPUT29), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n724), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT30), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT93), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n622), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n512), .A2(new_n513), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n740), .A2(new_n741), .A3(new_n579), .A4(new_n485), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n622), .A2(new_n739), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n738), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  AND3_X1   g0544(.A1(new_n485), .A2(new_n741), .A3(new_n579), .ZN(new_n745));
  INV_X1    g0545(.A(new_n743), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n745), .A2(KEYINPUT30), .A3(new_n746), .A4(new_n740), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n579), .A2(new_n509), .ZN(new_n748));
  AOI21_X1  g0548(.A(G179), .B1(new_n597), .B2(new_n602), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n748), .A2(new_n538), .A3(new_n649), .A4(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT94), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n485), .A2(new_n741), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n753), .A2(KEYINPUT94), .A3(new_n748), .A4(new_n749), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n744), .A2(new_n747), .A3(new_n752), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(new_n697), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT31), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n744), .A2(new_n747), .A3(new_n750), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n698), .A2(new_n757), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n636), .A2(new_n594), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT95), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n763), .A2(new_n764), .A3(new_n679), .A4(new_n698), .ZN(new_n765));
  AND3_X1   g0565(.A1(new_n628), .A2(new_n633), .A3(new_n635), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n679), .A2(new_n704), .A3(new_n766), .A4(new_n698), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(KEYINPUT95), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n762), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G330), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n737), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT97), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n719), .B1(new_n773), .B2(G1), .ZN(G364));
  AOI21_X1  g0574(.A(new_n225), .B1(G20), .B2(new_n297), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n204), .A2(new_n372), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT99), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n777), .A2(G190), .A3(G200), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G311), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n204), .A2(G179), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n293), .A2(new_n295), .A3(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G283), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n779), .A2(new_n780), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n293), .A2(G190), .A3(new_n781), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n784), .B1(G303), .B2(new_n786), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n295), .A2(G179), .A3(G200), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n204), .ZN(new_n789));
  INV_X1    g0589(.A(G294), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G190), .A2(G200), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n781), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n280), .B1(new_n794), .B2(G329), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n776), .A2(G200), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(G190), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  XOR2_X1   g0598(.A(KEYINPUT33), .B(G317), .Z(new_n799));
  OAI21_X1  g0599(.A(new_n795), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n376), .A2(new_n796), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n791), .B(new_n800), .C1(G326), .C2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G322), .ZN(new_n803));
  NOR3_X1   g0603(.A1(new_n777), .A2(G200), .A3(new_n376), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT100), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n787), .B(new_n802), .C1(new_n803), .C2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT102), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n808), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G58), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n798), .A2(new_n211), .B1(new_n789), .B2(new_n465), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n814), .A2(KEYINPUT101), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n794), .A2(G159), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n816), .A2(KEYINPUT32), .B1(new_n801), .B2(G50), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n817), .B(new_n280), .C1(KEYINPUT32), .C2(new_n816), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(KEYINPUT101), .B2(new_n814), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n782), .A2(new_n283), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n785), .A2(new_n213), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n820), .B(new_n821), .C1(new_n778), .C2(G77), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n813), .A2(new_n815), .A3(new_n819), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n811), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n809), .A2(new_n810), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n775), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n687), .A2(G20), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n203), .B1(new_n827), .B2(G45), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n714), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n713), .A2(new_n288), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n832), .A2(G355), .B1(new_n606), .B2(new_n713), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n342), .A2(new_n343), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n713), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(G45), .B2(new_n224), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n244), .A2(new_n452), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n833), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(G13), .A2(G33), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(G20), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n841), .A2(new_n775), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n831), .B1(new_n838), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n841), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n826), .B(new_n843), .C1(new_n701), .C2(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n701), .A2(G330), .ZN(new_n846));
  XOR2_X1   g0646(.A(new_n846), .B(KEYINPUT98), .Z(new_n847));
  NAND2_X1  g0647(.A1(new_n702), .A2(new_n831), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n845), .B1(new_n847), .B2(new_n848), .ZN(G396));
  AOI21_X1  g0649(.A(new_n697), .B1(new_n720), .B2(new_n721), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n296), .B1(new_n268), .B2(new_n698), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n299), .ZN(new_n852));
  OR2_X1    g0652(.A1(new_n299), .A2(new_n697), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n850), .B(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n771), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n830), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n857), .B2(new_n856), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n288), .B1(new_n793), .B2(new_n780), .ZN(new_n860));
  INV_X1    g0660(.A(new_n801), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n861), .A2(new_n600), .B1(new_n798), .B2(new_n783), .ZN(new_n862));
  INV_X1    g0662(.A(new_n789), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n860), .B(new_n862), .C1(G97), .C2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n785), .A2(new_n283), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n782), .A2(new_n213), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n865), .B(new_n866), .C1(new_n778), .C2(G116), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n864), .B(new_n867), .C1(new_n790), .C2(new_n808), .ZN(new_n868));
  INV_X1    g0668(.A(new_n834), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(G132), .B2(new_n794), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n782), .A2(new_n211), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(G50), .B2(new_n786), .ZN(new_n872));
  INV_X1    g0672(.A(G58), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n870), .B(new_n872), .C1(new_n873), .C2(new_n789), .ZN(new_n874));
  XOR2_X1   g0674(.A(new_n874), .B(KEYINPUT103), .Z(new_n875));
  AOI22_X1  g0675(.A1(G137), .A2(new_n801), .B1(new_n797), .B2(G150), .ZN(new_n876));
  INV_X1    g0676(.A(G143), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n876), .B1(new_n333), .B2(new_n779), .C1(new_n808), .C2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n875), .B1(new_n879), .B2(KEYINPUT34), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT34), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n868), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n775), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n775), .A2(new_n839), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n831), .B1(new_n258), .B2(new_n885), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n884), .B(new_n886), .C1(new_n855), .C2(new_n840), .ZN(new_n887));
  AND2_X1   g0687(.A1(new_n859), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(G384));
  INV_X1    g0689(.A(KEYINPUT105), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n361), .B2(new_n374), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT37), .B1(new_n361), .B2(new_n380), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n388), .A2(new_n694), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n388), .A2(new_n389), .A3(KEYINPUT105), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n891), .A2(new_n892), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n382), .B1(new_n383), .B2(new_n385), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n350), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n330), .B1(new_n349), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n392), .B1(new_n898), .B2(new_n695), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n898), .A2(new_n374), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT37), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n895), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n898), .A2(new_n695), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n395), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n902), .A2(new_n904), .A3(KEYINPUT38), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT38), .B1(new_n902), .B2(new_n904), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT39), .ZN(new_n908));
  NOR3_X1   g0708(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n893), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n395), .A2(KEYINPUT106), .A3(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n891), .A2(new_n894), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT37), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n893), .A2(new_n914), .A3(new_n392), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n893), .B(new_n392), .C1(new_n361), .C2(new_n374), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n913), .A2(new_n915), .B1(new_n916), .B2(KEYINPUT37), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT106), .B1(new_n395), .B2(new_n910), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n912), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n905), .B1(new_n919), .B2(KEYINPUT38), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n909), .B1(new_n920), .B2(new_n908), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n439), .A2(new_n411), .A3(new_n698), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n639), .A2(new_n694), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n411), .A2(new_n697), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n640), .A2(new_n927), .A3(new_n642), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n411), .B(new_n697), .C1(new_n439), .C2(new_n431), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n722), .A2(new_n698), .A3(new_n855), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n930), .B1(new_n931), .B2(new_n853), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n906), .A2(new_n907), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n926), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT108), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT107), .B1(new_n737), .B2(new_n442), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT107), .ZN(new_n938));
  AOI211_X1 g0738(.A(new_n938), .B(new_n441), .C1(new_n724), .C2(new_n736), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n648), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n936), .B(new_n940), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n920), .A2(KEYINPUT40), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n768), .A2(new_n765), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n756), .A2(new_n757), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT31), .B1(new_n755), .B2(new_n697), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n854), .B1(new_n928), .B2(new_n929), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n933), .A2(new_n947), .A3(new_n948), .ZN(new_n950));
  XOR2_X1   g0750(.A(KEYINPUT109), .B(KEYINPUT40), .Z(new_n951));
  AOI22_X1  g0751(.A1(new_n942), .A2(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n442), .A2(new_n947), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n952), .B1(new_n442), .B2(new_n947), .ZN(new_n956));
  NOR3_X1   g0756(.A1(new_n955), .A2(new_n956), .A3(new_n770), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n941), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n941), .A2(new_n957), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n958), .B(new_n959), .C1(new_n203), .C2(new_n827), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n606), .B(new_n227), .C1(new_n533), .C2(KEYINPUT35), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(KEYINPUT35), .B2(new_n533), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT36), .ZN(new_n963));
  OAI21_X1  g0763(.A(G77), .B1(new_n873), .B2(new_n211), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n224), .A2(new_n964), .B1(G50), .B2(new_n211), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n965), .A2(G1), .A3(new_n687), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT104), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n960), .A2(new_n968), .ZN(G367));
  INV_X1    g0769(.A(new_n773), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n530), .B(new_n540), .C1(new_n537), .C2(new_n698), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n697), .A2(new_n515), .A3(new_n659), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n711), .A2(new_n973), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT45), .Z(new_n975));
  NOR2_X1   g0775(.A1(new_n711), .A2(new_n973), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT44), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n975), .A2(new_n708), .A3(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT111), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n978), .A2(new_n979), .ZN(new_n981));
  INV_X1    g0781(.A(new_n708), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n975), .A2(new_n977), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n980), .A2(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n705), .A2(new_n710), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n707), .B2(new_n710), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(new_n703), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n970), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n714), .B(KEYINPUT41), .Z(new_n989));
  OAI21_X1  g0789(.A(new_n828), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n698), .A2(new_n491), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n991), .A2(new_n478), .A3(new_n461), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n673), .B2(new_n991), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n705), .A2(new_n710), .A3(new_n973), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT42), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n973), .A2(new_n594), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n697), .B1(new_n997), .B2(new_n530), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n994), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT110), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1000), .B(new_n1001), .Z(new_n1002));
  INV_X1    g0802(.A(new_n973), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n708), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n990), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n835), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n842), .B1(new_n207), .B2(new_n252), .C1(new_n1009), .C2(new_n237), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n1010), .A2(new_n830), .ZN(new_n1011));
  INV_X1    g0811(.A(G317), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n869), .B1(new_n1012), .B2(new_n793), .C1(new_n779), .C2(new_n783), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n782), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1013), .B1(G97), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n812), .A2(G303), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n861), .A2(new_n780), .B1(new_n283), .B2(new_n789), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(G294), .B2(new_n797), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n786), .A2(G116), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT46), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1015), .A2(new_n1016), .A3(new_n1018), .A4(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n782), .A2(new_n258), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n779), .B2(new_n303), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(G58), .B2(new_n786), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n861), .A2(new_n877), .B1(new_n798), .B2(new_n333), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n789), .A2(new_n211), .ZN(new_n1027));
  INV_X1    g0827(.A(G137), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n280), .B1(new_n793), .B2(new_n1028), .ZN(new_n1029));
  NOR3_X1   g0829(.A1(new_n1026), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1025), .B(new_n1030), .C1(new_n301), .C2(new_n808), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1021), .A2(new_n1031), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT47), .Z(new_n1033));
  INV_X1    g0833(.A(new_n775), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1011), .B1(new_n844), .B2(new_n993), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1008), .A2(new_n1035), .ZN(G387));
  AND2_X1   g0836(.A1(new_n773), .A2(new_n987), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1037), .A2(new_n715), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n773), .B2(new_n987), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n987), .A2(new_n829), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n808), .A2(new_n1012), .B1(new_n600), .B2(new_n779), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1041), .A2(KEYINPUT113), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(KEYINPUT113), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G322), .A2(new_n801), .B1(new_n797), .B2(G311), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT48), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n786), .A2(G294), .B1(new_n863), .B2(G283), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT49), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n782), .A2(new_n606), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n834), .B(new_n1054), .C1(G326), .C2(new_n794), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1052), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n863), .A2(new_n251), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n808), .B2(new_n303), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT112), .Z(new_n1059));
  OAI21_X1  g0859(.A(new_n834), .B1(new_n301), .B2(new_n793), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n861), .A2(new_n333), .B1(new_n798), .B2(new_n255), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n786), .A2(G77), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(new_n465), .B2(new_n782), .C1(new_n779), .C2(new_n211), .ZN(new_n1063));
  OR4_X1    g0863(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .A4(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1034), .B1(new_n1056), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n716), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n832), .A2(new_n1066), .B1(new_n283), .B2(new_n713), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n234), .A2(new_n452), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n255), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n303), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT50), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n716), .B(new_n452), .C1(new_n211), .C2(new_n258), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n835), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1067), .B1(new_n1068), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n831), .B1(new_n1074), .B2(new_n842), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n707), .B2(new_n844), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1039), .B(new_n1040), .C1(new_n1065), .C2(new_n1076), .ZN(G393));
  NAND2_X1  g0877(.A1(new_n983), .A2(new_n982), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT114), .Z(new_n1079));
  AND2_X1   g0879(.A1(new_n980), .A2(new_n981), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OR2_X1    g0881(.A1(new_n1081), .A2(new_n1037), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n715), .B1(new_n1037), .B2(new_n984), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1081), .A2(new_n829), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n835), .A2(new_n241), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n841), .B(new_n775), .C1(new_n713), .C2(G97), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n831), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n866), .B(new_n869), .C1(G143), .C2(new_n794), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n211), .B2(new_n785), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT115), .Z(new_n1091));
  NAND2_X1  g0891(.A1(new_n778), .A2(new_n1069), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n863), .A2(G77), .B1(new_n797), .B2(G50), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n808), .A2(new_n333), .B1(new_n301), .B2(new_n861), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT51), .Z(new_n1096));
  OAI22_X1  g0896(.A1(new_n808), .A2(new_n780), .B1(new_n1012), .B2(new_n861), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT52), .Z(new_n1098));
  AOI22_X1  g0898(.A1(new_n863), .A2(G116), .B1(new_n797), .B2(G303), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n779), .B2(new_n790), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT116), .Z(new_n1101));
  NAND2_X1  g0901(.A1(new_n786), .A2(G283), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n280), .B(new_n820), .C1(G322), .C2(new_n794), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n1094), .A2(new_n1096), .B1(new_n1098), .B2(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT117), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n1088), .B1(new_n844), .B2(new_n973), .C1(new_n1106), .C2(new_n1034), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1084), .A2(new_n1085), .A3(new_n1107), .ZN(G390));
  NOR4_X1   g0908(.A1(new_n769), .A2(new_n930), .A3(new_n770), .A4(new_n854), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n734), .A2(new_n698), .A3(new_n852), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n930), .B1(new_n1110), .B2(new_n853), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n395), .A2(new_n910), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT106), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n916), .A2(KEYINPUT37), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1112), .A2(new_n1113), .B1(new_n1114), .B2(new_n895), .ZN(new_n1115));
  AOI21_X1  g0915(.A(KEYINPUT38), .B1(new_n1115), .B2(new_n911), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n922), .B1(new_n1116), .B2(new_n906), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1111), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n853), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n850), .B2(new_n855), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n922), .B1(new_n1120), .B2(new_n930), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n909), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1116), .A2(new_n906), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1122), .B1(new_n1123), .B2(KEYINPUT39), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n1109), .B(new_n1118), .C1(new_n1121), .C2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT118), .ZN(new_n1126));
  AND4_X1   g0926(.A1(new_n1126), .A2(new_n947), .A3(G330), .A4(new_n948), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n770), .B1(new_n943), .B2(new_n946), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1126), .B1(new_n1128), .B2(new_n948), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1124), .B1(new_n932), .B2(new_n923), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1118), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1130), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1125), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n829), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n831), .B1(new_n255), .B2(new_n885), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n288), .B1(new_n793), .B2(new_n790), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n861), .A2(new_n783), .B1(new_n798), .B2(new_n283), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n1137), .B(new_n1138), .C1(G77), .C2(new_n863), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n821), .B(new_n871), .C1(new_n778), .C2(G97), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(G116), .B2(new_n812), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n812), .A2(G132), .B1(G128), .B2(new_n801), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT121), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(KEYINPUT54), .B(G143), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n779), .A2(new_n1145), .B1(new_n782), .B2(new_n303), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n786), .A2(G150), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT53), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n288), .B1(new_n794), .B2(G125), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n1149), .B1(new_n333), .B2(new_n789), .C1(new_n798), .C2(new_n1028), .ZN(new_n1150));
  NOR3_X1   g0950(.A1(new_n1146), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1142), .B1(new_n1144), .B2(new_n1151), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1136), .B1(new_n1152), .B2(new_n1034), .C1(new_n921), .C2(new_n840), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1135), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT119), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n947), .A2(G330), .A3(new_n948), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(KEYINPUT118), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n945), .B1(new_n759), .B2(new_n760), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n764), .B1(new_n637), .B2(new_n698), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n765), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1159), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1162), .A2(G330), .A3(new_n855), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n930), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1128), .A2(new_n1126), .A3(new_n948), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1158), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1120), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1110), .A2(new_n853), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n770), .B(new_n854), .C1(new_n943), .C2(new_n1159), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n930), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1169), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1128), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n930), .B1(new_n1173), .B2(new_n854), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1168), .A2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1173), .A2(new_n441), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n723), .B1(new_n734), .B2(new_n698), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n723), .B2(new_n850), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n938), .B1(new_n1179), .B2(new_n441), .ZN(new_n1180));
  NOR3_X1   g0980(.A1(new_n684), .A2(KEYINPUT29), .A3(new_n697), .ZN(new_n1181));
  OAI211_X1 g0981(.A(KEYINPUT107), .B(new_n442), .C1(new_n1181), .C2(new_n1178), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n647), .B(new_n1177), .C1(new_n1180), .C2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1176), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1158), .A2(new_n1165), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n684), .A2(new_n697), .A3(new_n854), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1171), .B1(new_n1186), .B2(new_n1119), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n921), .B1(new_n1187), .B2(new_n922), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1185), .B1(new_n1188), .B2(new_n1118), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1109), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1131), .A2(new_n1132), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1156), .B1(new_n1184), .B2(new_n1192), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1166), .A2(new_n1167), .B1(new_n1174), .B2(new_n1172), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1177), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n648), .B(new_n1195), .C1(new_n937), .C2(new_n939), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1134), .A2(new_n1197), .A3(KEYINPUT119), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1193), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT120), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n1134), .B2(new_n1197), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1184), .A2(KEYINPUT120), .A3(new_n1192), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1202), .A2(new_n714), .A3(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1155), .B1(new_n1200), .B2(new_n1204), .ZN(G378));
  AOI22_X1  g1005(.A1(new_n863), .A2(G150), .B1(new_n797), .B2(G132), .ZN(new_n1206));
  INV_X1    g1006(.A(G125), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1206), .B1(new_n1207), .B2(new_n861), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n779), .A2(new_n1028), .B1(new_n785), .B2(new_n1145), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1208), .B(new_n1209), .C1(new_n812), .C2(G128), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT59), .ZN(new_n1211));
  OR2_X1    g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1014), .A2(G159), .ZN(new_n1213));
  AOI211_X1 g1013(.A(G33), .B(G41), .C1(new_n794), .C2(G124), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(new_n1211), .B2(new_n1210), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n834), .A2(G41), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n303), .B1(G33), .B2(G41), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n782), .A2(new_n873), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1217), .A2(new_n1062), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1220), .B(new_n1221), .C1(new_n251), .C2(new_n778), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n861), .A2(new_n606), .B1(new_n798), .B2(new_n465), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n1027), .B(new_n1223), .C1(G283), .C2(new_n794), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1222), .B(new_n1224), .C1(new_n283), .C2(new_n808), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT58), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1219), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n1226), .B2(new_n1225), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n775), .B1(new_n1216), .B2(new_n1228), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1229), .B(KEYINPUT122), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n885), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n830), .B1(G50), .B2(new_n1231), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(KEYINPUT123), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1230), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n645), .A2(new_n317), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n695), .A2(new_n308), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1235), .B(new_n1236), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1237), .B(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(new_n839), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1234), .A2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n952), .A2(G330), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n924), .A2(new_n925), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n934), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1239), .A2(KEYINPUT124), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n952), .B(G330), .C1(new_n926), .C2(new_n934), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1246), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1241), .B1(new_n1250), .B2(new_n828), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NOR3_X1   g1052(.A1(new_n1184), .A2(new_n1192), .A3(new_n1156), .ZN(new_n1253));
  AOI21_X1  g1053(.A(KEYINPUT119), .B1(new_n1134), .B2(new_n1197), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1183), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  OR2_X1    g1055(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT57), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1196), .B1(new_n1193), .B2(new_n1198), .ZN(new_n1258));
  OAI21_X1  g1058(.A(KEYINPUT57), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n714), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1252), .B1(new_n1257), .B2(new_n1260), .ZN(G375));
  NAND2_X1  g1061(.A1(new_n930), .A2(new_n839), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n830), .B1(G68), .B2(new_n1231), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(G294), .A2(new_n801), .B1(new_n797), .B2(G116), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n779), .B2(new_n283), .ZN(new_n1265));
  XOR2_X1   g1065(.A(new_n1265), .B(KEYINPUT125), .Z(new_n1266));
  AOI21_X1  g1066(.A(new_n280), .B1(new_n794), .B2(G303), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1023), .A2(new_n1057), .A3(new_n1267), .ZN(new_n1268));
  OAI221_X1 g1068(.A(new_n1268), .B1(new_n465), .B2(new_n785), .C1(new_n808), .C2(new_n783), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n808), .A2(new_n1028), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n1220), .B(new_n869), .C1(G128), .C2(new_n794), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n798), .A2(new_n1145), .B1(new_n789), .B2(new_n303), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(G132), .B2(new_n801), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n778), .A2(G150), .B1(G159), .B2(new_n786), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1271), .A2(new_n1273), .A3(new_n1274), .ZN(new_n1275));
  OAI22_X1  g1075(.A1(new_n1266), .A2(new_n1269), .B1(new_n1270), .B2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1263), .B1(new_n1276), .B2(new_n775), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n1176), .A2(new_n829), .B1(new_n1262), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1197), .A2(new_n989), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1279), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(G381));
  NOR2_X1   g1083(.A1(G393), .A2(G396), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1085), .A2(new_n1107), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1285), .B1(new_n1083), .B2(new_n1082), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1284), .A2(new_n1286), .A3(new_n888), .A4(new_n1282), .ZN(new_n1287));
  OR4_X1    g1087(.A1(G387), .A2(new_n1287), .A3(G378), .A4(G375), .ZN(G407));
  AND3_X1   g1088(.A1(new_n1202), .A2(new_n714), .A3(new_n1203), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1154), .B1(new_n1289), .B2(new_n1199), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n696), .A2(G213), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1293));
  OAI211_X1 g1093(.A(G407), .B(G213), .C1(G375), .C2(new_n1293), .ZN(G409));
  AND2_X1   g1094(.A1(G393), .A2(G396), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1295), .A2(new_n1284), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(G390), .A2(new_n1008), .A3(new_n1035), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1286), .A2(G387), .ZN(new_n1298));
  AND3_X1   g1098(.A1(new_n1296), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1296), .B1(new_n1298), .B2(new_n1297), .ZN(new_n1300));
  NOR3_X1   g1100(.A1(new_n1299), .A2(new_n1300), .A3(KEYINPUT61), .ZN(new_n1301));
  OAI211_X1 g1101(.A(G378), .B(new_n1252), .C1(new_n1257), .C2(new_n1260), .ZN(new_n1302));
  NOR3_X1   g1102(.A1(new_n1258), .A2(new_n989), .A3(new_n1250), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1290), .B1(new_n1303), .B2(new_n1251), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1292), .B1(new_n1302), .B2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1194), .A2(new_n1196), .A3(KEYINPUT60), .ZN(new_n1306));
  AND2_X1   g1106(.A1(new_n1306), .A2(new_n714), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT60), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1281), .B1(new_n1197), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1307), .A2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1310), .A2(G384), .A3(new_n1278), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(G384), .B1(new_n1310), .B2(new_n1278), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1305), .A2(KEYINPUT63), .A3(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1302), .A2(new_n1304), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1291), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1292), .A2(G2897), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1314), .A2(new_n1318), .ZN(new_n1319));
  OAI211_X1 g1119(.A(G2897), .B(new_n1292), .C1(new_n1312), .C2(new_n1313), .ZN(new_n1320));
  AND2_X1   g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1317), .A2(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1316), .A2(new_n1291), .A3(new_n1314), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT63), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1301), .A2(new_n1315), .A3(new_n1322), .A4(new_n1325), .ZN(new_n1326));
  OR2_X1    g1126(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1329), .B1(new_n1305), .B2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT62), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1323), .A2(new_n1332), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1305), .A2(KEYINPUT62), .A3(new_n1314), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1331), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT127), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1327), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1328), .B1(new_n1317), .B2(new_n1321), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1334), .ZN(new_n1339));
  AOI21_X1  g1139(.A(KEYINPUT62), .B1(new_n1305), .B2(new_n1314), .ZN(new_n1340));
  OAI211_X1 g1140(.A(new_n1336), .B(new_n1338), .C1(new_n1339), .C2(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1341), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1326), .B1(new_n1337), .B2(new_n1342), .ZN(G405));
  NAND2_X1  g1143(.A1(G375), .A2(new_n1290), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1344), .A2(new_n1302), .ZN(new_n1345));
  XNOR2_X1  g1145(.A(new_n1345), .B(new_n1314), .ZN(new_n1346));
  XNOR2_X1  g1146(.A(new_n1327), .B(new_n1346), .ZN(G402));
endmodule


