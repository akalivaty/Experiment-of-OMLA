//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 0 0 0 0 0 0 0 1 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n562, new_n563, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n608, new_n609, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1201, new_n1202, new_n1203,
    new_n1204;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT66), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT68), .Z(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n451), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n452), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  OR2_X1    g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(G137), .A3(new_n465), .ZN(new_n466));
  AND3_X1   g041(.A1(new_n465), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(KEYINPUT69), .B1(new_n465), .B2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(G101), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(G125), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n465), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n470), .A2(new_n475), .ZN(G160));
  AOI21_X1  g051(.A(new_n465), .B1(new_n462), .B2(new_n463), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT70), .ZN(new_n479));
  AOI21_X1  g054(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n465), .A2(G112), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n479), .B(new_n481), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n487), .B1(new_n471), .B2(new_n472), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT72), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n487), .B(KEYINPUT72), .C1(new_n472), .C2(new_n471), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n490), .A2(KEYINPUT4), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n488), .A2(new_n489), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n477), .A2(G126), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT71), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n465), .A2(G114), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(G114), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n500), .A2(new_n502), .A3(KEYINPUT71), .A4(G2104), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n492), .A2(new_n494), .A3(new_n495), .A4(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT5), .B(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G62), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT73), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n509), .A2(new_n510), .B1(G75), .B2(G543), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n508), .A2(KEYINPUT73), .A3(G62), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n507), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  AND2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n508), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n514), .A2(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n513), .A2(new_n521), .ZN(G166));
  NOR2_X1   g097(.A1(new_n515), .A2(new_n516), .ZN(new_n523));
  INV_X1    g098(.A(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n525), .A2(G51), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  XOR2_X1   g105(.A(KEYINPUT5), .B(G543), .Z(new_n531));
  NAND2_X1  g106(.A1(new_n517), .A2(G89), .ZN(new_n532));
  NAND2_X1  g107(.A1(G63), .A2(G651), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n530), .A2(new_n534), .ZN(G168));
  NOR2_X1   g110(.A1(new_n531), .A2(new_n523), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G90), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n525), .A2(G52), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(KEYINPUT74), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT74), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n537), .A2(new_n541), .A3(new_n538), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(new_n507), .ZN(new_n545));
  AND3_X1   g120(.A1(new_n543), .A2(KEYINPUT75), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g121(.A(KEYINPUT75), .B1(new_n543), .B2(new_n545), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n546), .A2(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  INV_X1    g124(.A(G43), .ZN(new_n550));
  INV_X1    g125(.A(G81), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n550), .A2(new_n518), .B1(new_n519), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(new_n507), .ZN(new_n554));
  OR2_X1    g129(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(KEYINPUT76), .ZN(new_n556));
  OR3_X1    g131(.A1(new_n552), .A2(KEYINPUT76), .A3(new_n554), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  NAND2_X1  g139(.A1(new_n525), .A2(G53), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n531), .B2(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n569), .A2(G651), .B1(new_n536), .B2(G91), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(G299));
  INV_X1    g146(.A(G168), .ZN(G286));
  OR2_X1    g147(.A1(new_n513), .A2(new_n521), .ZN(G303));
  NAND2_X1  g148(.A1(new_n525), .A2(G49), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n575));
  AND2_X1   g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(G87), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n519), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n576), .A2(new_n579), .ZN(G288));
  NAND2_X1  g155(.A1(new_n508), .A2(G61), .ZN(new_n581));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n507), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT77), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n583), .B(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n536), .A2(G86), .B1(new_n525), .B2(G48), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(G305));
  INV_X1    g162(.A(G47), .ZN(new_n588));
  INV_X1    g163(.A(G85), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n588), .A2(new_n518), .B1(new_n519), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(new_n507), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(new_n536), .A2(G92), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G66), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n531), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n600), .A2(G651), .B1(new_n525), .B2(G54), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(G171), .B2(G868), .ZN(G321));
  XOR2_X1   g179(.A(G321), .B(KEYINPUT78), .Z(G284));
  MUX2_X1   g180(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g181(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g182(.A(new_n602), .ZN(new_n608));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G860), .ZN(G148));
  NAND2_X1  g185(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(new_n559), .B2(G868), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g189(.A1(new_n480), .A2(G135), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT79), .ZN(new_n616));
  OAI21_X1  g191(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n617));
  INV_X1    g192(.A(G111), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G2105), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n619), .B1(G123), .B2(new_n477), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(G2096), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n467), .A2(new_n468), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(new_n464), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT13), .Z(new_n627));
  OAI21_X1  g202(.A(new_n623), .B1(new_n627), .B2(G2100), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(G2100), .B2(new_n627), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT80), .ZN(G156));
  XNOR2_X1  g205(.A(G2427), .B(G2438), .ZN(new_n631));
  INV_X1    g206(.A(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n631), .B(G2430), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(new_n634), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n636), .A2(new_n638), .A3(KEYINPUT14), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(KEYINPUT82), .ZN(new_n640));
  INV_X1    g215(.A(G1341), .ZN(new_n641));
  INV_X1    g216(.A(KEYINPUT82), .ZN(new_n642));
  NAND4_X1  g217(.A1(new_n636), .A2(new_n638), .A3(new_n642), .A4(KEYINPUT14), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n641), .B1(new_n640), .B2(new_n643), .ZN(new_n646));
  OAI21_X1  g221(.A(G1348), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(new_n646), .ZN(new_n648));
  INV_X1    g223(.A(G1348), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(new_n649), .A3(new_n644), .ZN(new_n650));
  XOR2_X1   g225(.A(G2451), .B(G2454), .Z(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n653), .B(new_n654), .Z(new_n655));
  NAND3_X1  g230(.A1(new_n647), .A2(new_n650), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(G14), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n655), .B1(new_n647), .B2(new_n650), .ZN(new_n658));
  OAI21_X1  g233(.A(KEYINPUT83), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n647), .A2(new_n650), .ZN(new_n660));
  INV_X1    g235(.A(new_n655), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT83), .ZN(new_n663));
  NAND4_X1  g238(.A1(new_n662), .A2(new_n663), .A3(G14), .A4(new_n656), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n659), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT84), .Z(G401));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2072), .B(G2078), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n669), .A2(KEYINPUT85), .ZN(new_n670));
  XOR2_X1   g245(.A(G2067), .B(G2678), .Z(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(KEYINPUT85), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(new_n672), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT17), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n668), .B(new_n673), .C1(new_n676), .C2(new_n671), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n668), .A2(new_n671), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT18), .Z(new_n680));
  NAND3_X1  g255(.A1(new_n676), .A2(new_n671), .A3(new_n667), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n677), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(G2096), .ZN(new_n683));
  NAND4_X1  g258(.A1(new_n677), .A2(new_n680), .A3(new_n622), .A4(new_n681), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT86), .B(G2100), .ZN(new_n685));
  AND3_X1   g260(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n685), .B1(new_n683), .B2(new_n684), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(G227));
  XOR2_X1   g263(.A(G1971), .B(G1976), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT19), .ZN(new_n690));
  XOR2_X1   g265(.A(G1956), .B(G2474), .Z(new_n691));
  XOR2_X1   g266(.A(G1961), .B(G1966), .Z(new_n692));
  AND2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT20), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n691), .A2(new_n692), .ZN(new_n696));
  NOR3_X1   g271(.A1(new_n690), .A2(new_n693), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n690), .B2(new_n696), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(G1991), .B(G1996), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT87), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n701), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1981), .B(G1986), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(G229));
  NOR2_X1   g282(.A1(G4), .A2(G16), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT89), .Z(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n709), .B1(new_n602), .B2(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT91), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT90), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(new_n649), .ZN(new_n714));
  NOR2_X1   g289(.A1(G5), .A2(G16), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G171), .B2(G16), .ZN(new_n716));
  INV_X1    g291(.A(G1961), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n559), .A2(new_n710), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n710), .B2(G19), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT92), .B(G1341), .Z(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT25), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n725), .A2(new_n465), .ZN(new_n726));
  AOI211_X1 g301(.A(new_n724), .B(new_n726), .C1(G139), .C2(new_n480), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n728), .B2(G33), .ZN(new_n730));
  INV_X1    g305(.A(G2072), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT31), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n734), .A2(G11), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(G11), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT30), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n737), .A2(G28), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n728), .B1(new_n737), .B2(G28), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n735), .B(new_n736), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n621), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n740), .B1(new_n741), .B2(G29), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n722), .A2(new_n732), .A3(new_n733), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n728), .A2(G27), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G164), .B2(new_n728), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT96), .B(G2078), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(G286), .A2(new_n710), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT95), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(KEYINPUT95), .B1(G16), .B2(G21), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(new_n748), .B2(new_n751), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n752), .A2(G1966), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(G1966), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n480), .A2(G140), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n477), .A2(G128), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n465), .A2(G116), .ZN(new_n757));
  OAI21_X1  g332(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n755), .B(new_n756), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G29), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n728), .A2(G26), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT28), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(G2067), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  AND2_X1   g340(.A1(KEYINPUT24), .A2(G34), .ZN(new_n766));
  NOR2_X1   g341(.A1(KEYINPUT24), .A2(G34), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n728), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT93), .Z(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G160), .B2(G29), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(G2084), .Z(new_n771));
  NAND4_X1  g346(.A1(new_n753), .A2(new_n754), .A3(new_n765), .A4(new_n771), .ZN(new_n772));
  NOR3_X1   g347(.A1(new_n743), .A2(new_n747), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n728), .A2(G32), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n477), .A2(G129), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n480), .A2(G141), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G105), .B2(new_n624), .ZN(new_n778));
  NAND3_X1  g353(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT94), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT26), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n774), .B1(new_n783), .B2(new_n728), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT27), .ZN(new_n785));
  INV_X1    g360(.A(G1996), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n710), .A2(G20), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT97), .Z(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT23), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G299), .B2(G16), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G1956), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n720), .B2(new_n721), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n728), .A2(G35), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G162), .B2(new_n728), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT29), .B(G2090), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NOR3_X1   g372(.A1(new_n787), .A2(new_n793), .A3(new_n797), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n714), .A2(new_n718), .A3(new_n773), .A4(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT36), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n710), .A2(G24), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n593), .B2(new_n710), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1986), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n480), .A2(G131), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n477), .A2(G119), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n465), .A2(G107), .ZN(new_n806));
  OAI21_X1  g381(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n804), .B(new_n805), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  MUX2_X1   g383(.A(G25), .B(new_n808), .S(G29), .Z(new_n809));
  XOR2_X1   g384(.A(KEYINPUT35), .B(G1991), .Z(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n809), .B(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT88), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(new_n576), .B2(new_n579), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n815));
  NOR3_X1   g390(.A1(new_n815), .A2(new_n578), .A3(KEYINPUT88), .ZN(new_n816));
  OAI21_X1  g391(.A(G16), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(G23), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(G16), .B2(new_n818), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT33), .Z(new_n820));
  AND2_X1   g395(.A1(new_n820), .A2(G1976), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n820), .A2(G1976), .ZN(new_n822));
  MUX2_X1   g397(.A(G6), .B(G305), .S(G16), .Z(new_n823));
  XOR2_X1   g398(.A(KEYINPUT32), .B(G1981), .Z(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n710), .A2(G22), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G166), .B2(new_n710), .ZN(new_n827));
  INV_X1    g402(.A(G1971), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  NOR3_X1   g405(.A1(new_n821), .A2(new_n822), .A3(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT34), .ZN(new_n832));
  AOI211_X1 g407(.A(new_n803), .B(new_n812), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n800), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n833), .A2(new_n800), .A3(new_n834), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n799), .B1(new_n836), .B2(new_n837), .ZN(G311));
  INV_X1    g413(.A(new_n799), .ZN(new_n839));
  INV_X1    g414(.A(new_n837), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n840), .B2(new_n835), .ZN(G150));
  NOR2_X1   g416(.A1(new_n602), .A2(new_n609), .ZN(new_n842));
  XOR2_X1   g417(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(G93), .ZN(new_n845));
  XNOR2_X1  g420(.A(KEYINPUT99), .B(G55), .ZN(new_n846));
  OAI22_X1  g421(.A1(new_n845), .A2(new_n519), .B1(new_n518), .B2(new_n846), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n848), .A2(new_n507), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n851), .A2(new_n555), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n852), .B1(new_n558), .B2(new_n851), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n844), .B(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT39), .ZN(new_n855));
  AOI21_X1  g430(.A(G860), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(new_n855), .B2(new_n854), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n851), .A2(G860), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT100), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT37), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT101), .Z(G145));
  NOR2_X1   g437(.A1(new_n727), .A2(KEYINPUT103), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n782), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n759), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(G164), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n865), .A2(G164), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n480), .A2(G142), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n477), .A2(G130), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n465), .A2(G118), .ZN(new_n871));
  OAI21_X1  g446(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n869), .B(new_n870), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT104), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n626), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n808), .ZN(new_n876));
  OAI22_X1  g451(.A1(new_n867), .A2(new_n868), .B1(KEYINPUT105), .B2(new_n876), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n865), .A2(G164), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n876), .A2(KEYINPUT105), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(new_n866), .A3(new_n879), .ZN(new_n880));
  XOR2_X1   g455(.A(G160), .B(KEYINPUT102), .Z(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(G162), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n621), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n877), .A2(new_n880), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n876), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n886), .B1(new_n867), .B2(new_n868), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n878), .A2(new_n866), .A3(new_n876), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n887), .A2(new_n888), .A3(new_n883), .ZN(new_n889));
  INV_X1    g464(.A(G37), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n885), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g467(.A(KEYINPUT111), .B1(new_n850), .B2(G868), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n853), .A2(new_n611), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n850), .B1(new_n556), .B2(new_n557), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n602), .A2(G559), .ZN(new_n896));
  NOR3_X1   g471(.A1(new_n895), .A2(new_n896), .A3(new_n852), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n602), .A2(G299), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n597), .A2(new_n566), .A3(new_n570), .A4(new_n601), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n898), .A2(KEYINPUT41), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(KEYINPUT41), .B1(new_n898), .B2(new_n899), .ZN(new_n901));
  OAI22_X1  g476(.A1(new_n894), .A2(new_n897), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n853), .A2(new_n611), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n896), .B1(new_n895), .B2(new_n852), .ZN(new_n904));
  AOI21_X1  g479(.A(KEYINPUT106), .B1(new_n898), .B2(new_n899), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n898), .A2(KEYINPUT106), .A3(new_n899), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n903), .B(new_n904), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  AND2_X1   g482(.A1(new_n902), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(G305), .A2(G303), .ZN(new_n909));
  NAND3_X1  g484(.A1(G166), .A2(new_n586), .A3(new_n585), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(G290), .B1(new_n814), .B2(new_n816), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n576), .A2(new_n813), .A3(new_n579), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT88), .B1(new_n815), .B2(new_n578), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n913), .A2(new_n593), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n911), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n917), .A2(KEYINPUT107), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT107), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n919), .B1(new_n911), .B2(new_n916), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n909), .A2(new_n912), .A3(new_n915), .A4(new_n910), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n921), .A2(KEYINPUT108), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(KEYINPUT108), .ZN(new_n923));
  OAI22_X1  g498(.A1(new_n918), .A2(new_n920), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OR2_X1    g499(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n925));
  NAND2_X1  g500(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n917), .B(KEYINPUT107), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n921), .B(KEYINPUT108), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n928), .A2(new_n929), .A3(KEYINPUT109), .A4(KEYINPUT42), .ZN(new_n930));
  AOI211_X1 g505(.A(KEYINPUT110), .B(new_n908), .C1(new_n927), .C2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n908), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n927), .A2(new_n930), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT110), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI22_X1  g510(.A1(new_n931), .A2(new_n935), .B1(new_n934), .B2(new_n933), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n893), .B1(new_n936), .B2(G868), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT111), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n936), .A2(G868), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(G295));
  AOI21_X1  g515(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(G331));
  OAI21_X1  g516(.A(G168), .B1(new_n546), .B2(new_n547), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n543), .A2(new_n545), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT75), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n543), .A2(KEYINPUT75), .A3(new_n545), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n945), .A2(G286), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n942), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n853), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n942), .A2(new_n947), .A3(new_n853), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n950), .A2(new_n898), .A3(new_n899), .A4(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n900), .A2(new_n901), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n942), .A2(new_n947), .A3(new_n853), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n853), .B1(new_n942), .B2(new_n947), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n952), .A2(new_n956), .A3(new_n924), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n952), .A2(new_n956), .ZN(new_n959));
  INV_X1    g534(.A(new_n924), .ZN(new_n960));
  AOI21_X1  g535(.A(G37), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT112), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n958), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n924), .B1(new_n952), .B2(new_n956), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT112), .B1(new_n964), .B2(G37), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT43), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  NOR4_X1   g541(.A1(new_n954), .A2(new_n955), .A3(new_n905), .A4(new_n906), .ZN(new_n967));
  INV_X1    g542(.A(new_n956), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n960), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AND4_X1   g544(.A1(KEYINPUT43), .A2(new_n969), .A3(new_n890), .A4(new_n957), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT44), .B1(new_n966), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n972), .B1(new_n963), .B2(new_n965), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n969), .A2(new_n972), .A3(new_n890), .A4(new_n957), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n971), .B1(new_n976), .B2(KEYINPUT44), .ZN(G397));
  XNOR2_X1  g552(.A(KEYINPUT113), .B(G1384), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n505), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G40), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n470), .A2(new_n982), .A3(new_n475), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  OR3_X1    g561(.A1(new_n986), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT46), .B1(new_n986), .B2(G1996), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n759), .B(G2067), .ZN(new_n989));
  OR2_X1    g564(.A1(new_n989), .A2(new_n782), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n987), .A2(new_n988), .B1(new_n985), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g566(.A(new_n991), .B(KEYINPUT47), .Z(new_n992));
  NOR2_X1   g567(.A1(new_n759), .A2(G2067), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n985), .A2(new_n786), .A3(new_n783), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n994), .B(KEYINPUT114), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n783), .A2(new_n786), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n985), .B1(new_n996), .B2(new_n989), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n808), .A2(new_n811), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n993), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n992), .B1(new_n1000), .B2(new_n986), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n808), .A2(new_n811), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n985), .B1(new_n1002), .B2(new_n999), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n998), .A2(KEYINPUT125), .A3(new_n1003), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n986), .A2(G1986), .A3(G290), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n1005), .B(KEYINPUT48), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n998), .A2(new_n1003), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT125), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1001), .B1(new_n1004), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G1384), .ZN(new_n1011));
  AND3_X1   g586(.A1(new_n490), .A2(KEYINPUT4), .A3(new_n491), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n494), .A2(new_n504), .A3(new_n495), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1011), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT50), .ZN(new_n1015));
  INV_X1    g590(.A(G2090), .ZN(new_n1016));
  XOR2_X1   g591(.A(KEYINPUT116), .B(KEYINPUT50), .Z(new_n1017));
  NAND3_X1  g592(.A1(new_n505), .A2(new_n1011), .A3(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1015), .A2(new_n1016), .A3(new_n983), .A4(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT117), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n494), .A2(new_n504), .A3(new_n495), .ZN(new_n1021));
  AOI21_X1  g596(.A(G1384), .B1(new_n1021), .B2(new_n492), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n984), .B1(new_n1022), .B2(new_n1017), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT117), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1023), .A2(new_n1024), .A3(new_n1016), .A4(new_n1015), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n978), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(new_n983), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(new_n1022), .B2(KEYINPUT45), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1014), .A2(KEYINPUT115), .A3(new_n980), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1027), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1020), .B(new_n1025), .C1(new_n1031), .C2(G1971), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G8), .ZN(new_n1035));
  NOR2_X1   g610(.A1(G166), .A2(new_n1035), .ZN(new_n1036));
  XOR2_X1   g611(.A(new_n1036), .B(KEYINPUT55), .Z(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n980), .B1(new_n1021), .B2(new_n492), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n984), .B1(new_n1039), .B2(new_n978), .ZN(new_n1040));
  AOI211_X1 g615(.A(new_n1028), .B(KEYINPUT45), .C1(new_n505), .C2(new_n1011), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT115), .B1(new_n1014), .B2(new_n980), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1040), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(new_n828), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1044), .A2(KEYINPUT118), .A3(new_n1020), .A4(new_n1025), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1034), .A2(G8), .A3(new_n1038), .A4(new_n1045), .ZN(new_n1046));
  OAI211_X1 g621(.A(KEYINPUT45), .B(new_n1011), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n983), .B(new_n1047), .C1(new_n1022), .C2(KEYINPUT45), .ZN(new_n1048));
  INV_X1    g623(.A(G1966), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  XOR2_X1   g625(.A(KEYINPUT119), .B(G2084), .Z(new_n1051));
  NAND4_X1  g626(.A1(new_n1015), .A2(new_n983), .A3(new_n1018), .A4(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1050), .A2(G168), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(G8), .ZN(new_n1054));
  AOI21_X1  g629(.A(G168), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT51), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1053), .A2(new_n1057), .A3(G8), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G1981), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n583), .A2(new_n584), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n583), .A2(new_n584), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n586), .B(new_n1060), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n586), .ZN(new_n1064));
  OAI21_X1  g639(.A(G1981), .B1(new_n1064), .B2(new_n583), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT49), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1063), .A2(new_n1065), .A3(KEYINPUT49), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1035), .B1(new_n1022), .B2(new_n983), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n913), .A2(new_n914), .A3(G1976), .ZN(new_n1072));
  INV_X1    g647(.A(G1976), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT52), .B1(G288), .B2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1070), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT52), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1071), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT50), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n505), .A2(new_n1079), .A3(new_n1011), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1080), .B(new_n983), .C1(new_n1022), .C2(new_n1017), .ZN(new_n1081));
  OAI22_X1  g656(.A1(new_n1031), .A2(G1971), .B1(G2090), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(G8), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1078), .B1(new_n1083), .B2(new_n1037), .ZN(new_n1084));
  INV_X1    g659(.A(G2078), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1085), .B(new_n1040), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT53), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1048), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1087), .A2(G2078), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1015), .A2(new_n983), .A3(new_n1018), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1089), .A2(new_n1090), .B1(new_n1091), .B2(new_n717), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1088), .A2(new_n1092), .A3(G301), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1017), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n983), .B1(new_n1014), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1079), .B1(new_n505), .B2(new_n1011), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n717), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n981), .A2(new_n983), .A3(new_n1026), .A4(new_n1090), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1099), .B1(new_n1087), .B2(new_n1086), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1093), .B(KEYINPUT54), .C1(new_n1100), .C2(G301), .ZN(new_n1101));
  AND4_X1   g676(.A1(new_n1046), .A2(new_n1059), .A3(new_n1084), .A4(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(G299), .B(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g680(.A(KEYINPUT56), .B(G2072), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1040), .B(new_n1106), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1107));
  INV_X1    g682(.A(G1956), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1081), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1105), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT121), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(new_n1014), .B2(new_n984), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1022), .A2(KEYINPUT121), .A3(new_n983), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1114), .A2(new_n764), .B1(new_n1091), .B2(new_n649), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1115), .A2(new_n602), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1105), .B1(new_n1109), .B2(new_n1107), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1110), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT121), .B1(new_n1022), .B2(new_n983), .ZN(new_n1119));
  AND4_X1   g694(.A1(KEYINPUT121), .A2(new_n505), .A3(new_n983), .A4(new_n1011), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n764), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n649), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT60), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n602), .B1(new_n1115), .B2(KEYINPUT60), .ZN(new_n1126));
  AND4_X1   g701(.A1(KEYINPUT60), .A2(new_n1121), .A3(new_n602), .A4(new_n1122), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1125), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT61), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1110), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1129), .B1(new_n1130), .B2(new_n1117), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1105), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1135), .A2(KEYINPUT61), .A3(new_n1110), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT59), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n786), .B(new_n1040), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1138));
  XOR2_X1   g713(.A(KEYINPUT58), .B(G1341), .Z(new_n1139));
  NAND3_X1  g714(.A1(new_n1112), .A2(new_n1113), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1137), .B1(new_n1141), .B2(new_n559), .ZN(new_n1142));
  AOI211_X1 g717(.A(KEYINPUT59), .B(new_n558), .C1(new_n1138), .C2(new_n1140), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1136), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1118), .B1(new_n1132), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT54), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT122), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1100), .A2(new_n1147), .A3(G301), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1088), .A2(new_n1092), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(G171), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1147), .B1(new_n1100), .B2(G301), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1146), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1102), .A2(new_n1145), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT123), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1053), .A2(new_n1057), .A3(G8), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(G286), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1158), .A2(G8), .A3(new_n1053), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1156), .B1(new_n1159), .B2(KEYINPUT51), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT62), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1155), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1150), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1163));
  AND2_X1   g738(.A1(new_n1046), .A2(new_n1084), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1059), .A2(KEYINPUT123), .A3(KEYINPUT62), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .A4(new_n1165), .ZN(new_n1166));
  AOI211_X1 g741(.A(new_n1035), .B(G286), .C1(new_n1050), .C2(new_n1052), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1046), .A2(new_n1084), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT63), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1034), .A2(G8), .A3(new_n1045), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(new_n1037), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1078), .ZN(new_n1173));
  AND3_X1   g748(.A1(new_n1173), .A2(KEYINPUT63), .A3(new_n1167), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1172), .A2(new_n1046), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1170), .A2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1046), .A2(new_n1078), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1071), .A2(new_n1073), .A3(new_n579), .A4(new_n576), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(new_n1063), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1177), .B1(new_n1070), .B2(new_n1179), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1154), .A2(new_n1166), .A3(new_n1176), .A4(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n593), .B(G1986), .Z(new_n1183));
  AOI21_X1  g758(.A(new_n1007), .B1(new_n985), .B2(new_n1183), .ZN(new_n1184));
  AND3_X1   g759(.A1(new_n1181), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1182), .B1(new_n1181), .B2(new_n1184), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1010), .B1(new_n1185), .B2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g762(.A(new_n891), .B1(new_n973), .B2(new_n975), .ZN(new_n1189));
  OAI21_X1  g763(.A(G319), .B1(new_n686), .B2(new_n687), .ZN(new_n1190));
  INV_X1    g764(.A(new_n1190), .ZN(new_n1191));
  AOI21_X1  g765(.A(KEYINPUT126), .B1(new_n665), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n1193));
  AOI211_X1 g767(.A(new_n1193), .B(new_n1190), .C1(new_n659), .C2(new_n664), .ZN(new_n1194));
  OAI21_X1  g768(.A(new_n706), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n1196));
  NAND2_X1  g770(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  OAI211_X1 g771(.A(new_n706), .B(KEYINPUT127), .C1(new_n1192), .C2(new_n1194), .ZN(new_n1198));
  NAND2_X1  g772(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g773(.A1(new_n1189), .A2(new_n1199), .ZN(G308));
  NAND2_X1  g774(.A1(new_n961), .A2(new_n962), .ZN(new_n1201));
  NAND3_X1  g775(.A1(new_n1201), .A2(new_n965), .A3(new_n957), .ZN(new_n1202));
  NAND2_X1  g776(.A1(new_n1202), .A2(KEYINPUT43), .ZN(new_n1203));
  NAND2_X1  g777(.A1(new_n1203), .A2(new_n974), .ZN(new_n1204));
  NAND4_X1  g778(.A1(new_n1204), .A2(new_n891), .A3(new_n1198), .A4(new_n1197), .ZN(G225));
endmodule


