//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n549, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n561,
    new_n562, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n601, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1168, new_n1169;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT66), .Z(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT67), .Z(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n462), .A2(KEYINPUT70), .A3(G137), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n468), .A2(G137), .A3(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT70), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n465), .A2(G2105), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n463), .A2(new_n472), .B1(G101), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g049(.A(KEYINPUT68), .B1(new_n459), .B2(new_n460), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n466), .A2(new_n476), .A3(new_n467), .ZN(new_n477));
  AND3_X1   g052(.A1(new_n475), .A2(new_n477), .A3(G125), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT69), .ZN(new_n480));
  OAI21_X1  g055(.A(G2105), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n474), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  NAND2_X1  g058(.A1(new_n462), .A2(G136), .ZN(new_n484));
  NOR2_X1   g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(new_n469), .B2(G112), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g062(.A(G2105), .B1(new_n459), .B2(new_n460), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(KEYINPUT71), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT71), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2105), .C1(new_n459), .C2(new_n460), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n487), .B1(G124), .B2(new_n492), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n493), .B(KEYINPUT72), .ZN(G162));
  OAI21_X1  g069(.A(G2104), .B1(new_n469), .B2(G114), .ZN(new_n495));
  INV_X1    g070(.A(G102), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n495), .B1(new_n496), .B2(new_n469), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT73), .ZN(new_n498));
  INV_X1    g073(.A(G126), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n498), .B1(new_n488), .B2(new_n499), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n468), .A2(KEYINPUT73), .A3(G126), .A4(G2105), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n497), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n469), .A2(KEYINPUT4), .A3(G138), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n461), .A2(new_n503), .ZN(new_n504));
  AND2_X1   g079(.A1(new_n469), .A2(G138), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n475), .A2(new_n477), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n504), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n502), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  OR2_X1    g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G50), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n516), .A2(new_n522), .ZN(G166));
  NAND3_X1  g098(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n524));
  INV_X1    g099(.A(G51), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n524), .B1(new_n520), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  INV_X1    g103(.A(G89), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n528), .B1(new_n518), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT74), .ZN(new_n531));
  OR3_X1    g106(.A1(new_n526), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n526), .B2(new_n530), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(G168));
  AOI22_X1  g109(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n515), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  INV_X1    g112(.A(G52), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n518), .A2(new_n537), .B1(new_n520), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(G171));
  AOI22_X1  g115(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n515), .ZN(new_n542));
  INV_X1    g117(.A(G81), .ZN(new_n543));
  INV_X1    g118(.A(G43), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n518), .A2(new_n543), .B1(new_n520), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT75), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  NAND3_X1  g127(.A1(new_n517), .A2(G53), .A3(G543), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT9), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n513), .A2(new_n517), .A3(G91), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n513), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n556), .A2(new_n515), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n554), .A2(new_n555), .A3(new_n557), .ZN(G299));
  INV_X1    g133(.A(G171), .ZN(G301));
  INV_X1    g134(.A(G168), .ZN(G286));
  OR2_X1    g135(.A1(G166), .A2(KEYINPUT76), .ZN(new_n561));
  NAND2_X1  g136(.A1(G166), .A2(KEYINPUT76), .ZN(new_n562));
  AND2_X1   g137(.A1(new_n561), .A2(new_n562), .ZN(G303));
  NAND3_X1  g138(.A1(new_n517), .A2(G49), .A3(G543), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT77), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n566));
  INV_X1    g141(.A(G87), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n518), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(G288));
  INV_X1    g145(.A(G61), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n571), .B1(new_n511), .B2(new_n512), .ZN(new_n572));
  AND2_X1   g147(.A1(G73), .A2(G543), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n513), .A2(new_n517), .A3(G86), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n517), .A2(G48), .A3(G543), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G305));
  AOI22_X1  g152(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n578), .A2(new_n515), .ZN(new_n579));
  INV_X1    g154(.A(G85), .ZN(new_n580));
  XOR2_X1   g155(.A(KEYINPUT78), .B(G47), .Z(new_n581));
  OAI22_X1  g156(.A1(new_n518), .A2(new_n580), .B1(new_n520), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n583), .B(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n513), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G54), .ZN(new_n588));
  OAI22_X1  g163(.A1(new_n587), .A2(new_n515), .B1(new_n520), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT80), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n589), .B(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n513), .A2(new_n517), .A3(G92), .ZN(new_n592));
  XOR2_X1   g167(.A(new_n592), .B(KEYINPUT10), .Z(new_n593));
  NAND2_X1  g168(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n586), .B1(new_n595), .B2(G868), .ZN(G284));
  OAI21_X1  g171(.A(new_n586), .B1(new_n595), .B2(G868), .ZN(G321));
  NOR2_X1   g172(.A1(G299), .A2(G868), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g174(.A(new_n598), .B1(G868), .B2(G168), .ZN(G280));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n595), .B1(new_n601), .B2(G860), .ZN(G148));
  NAND2_X1  g177(.A1(new_n595), .A2(new_n601), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G868), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g181(.A1(new_n462), .A2(G135), .ZN(new_n607));
  NOR2_X1   g182(.A1(G99), .A2(G2105), .ZN(new_n608));
  OAI21_X1  g183(.A(G2104), .B1(new_n469), .B2(G111), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(G123), .B2(new_n492), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(KEYINPUT82), .Z(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(G2096), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n475), .A2(new_n477), .A3(new_n473), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT12), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT13), .Z(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G2100), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT81), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n613), .B(new_n618), .C1(G2100), .C2(new_n616), .ZN(G156));
  XOR2_X1   g194(.A(G2451), .B(G2454), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT16), .ZN(new_n621));
  XNOR2_X1  g196(.A(G1341), .B(G1348), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(G2443), .B(G2446), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2427), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT15), .B(G2435), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n629), .A2(new_n630), .A3(KEYINPUT14), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n625), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n625), .A2(new_n632), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n633), .A2(new_n634), .A3(G14), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(G401));
  XNOR2_X1  g211(.A(G2072), .B(G2078), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT17), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2067), .B(G2678), .ZN(new_n639));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  NOR3_X1   g216(.A1(new_n638), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT83), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n638), .A2(new_n639), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n644), .B(new_n641), .C1(new_n637), .C2(new_n639), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n640), .A2(new_n637), .A3(new_n639), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT18), .Z(new_n647));
  NAND3_X1  g222(.A1(new_n643), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(G2096), .Z(new_n649));
  OR2_X1    g224(.A1(new_n649), .A2(G2100), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(G2100), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(G227));
  XOR2_X1   g227(.A(G1971), .B(G1976), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT84), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT19), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1956), .B(G2474), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1961), .B(G1966), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT20), .ZN(new_n660));
  AND2_X1   g235(.A1(new_n656), .A2(new_n657), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n655), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n662), .B1(new_n655), .B2(new_n661), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1991), .B(G1996), .ZN(new_n665));
  INV_X1    g240(.A(G1981), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n664), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(KEYINPUT85), .B(G1986), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G229));
  INV_X1    g247(.A(KEYINPUT87), .ZN(new_n673));
  INV_X1    g248(.A(G29), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(G25), .ZN(new_n675));
  OR2_X1    g250(.A1(G95), .A2(G2105), .ZN(new_n676));
  INV_X1    g251(.A(G107), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n465), .B1(new_n677), .B2(G2105), .ZN(new_n678));
  AOI22_X1  g253(.A1(new_n462), .A2(G131), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(G119), .B2(new_n492), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n675), .B1(new_n681), .B2(new_n674), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT35), .B(G1991), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT86), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n673), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  MUX2_X1   g260(.A(G24), .B(G290), .S(G16), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(G1986), .ZN(new_n687));
  AOI211_X1 g262(.A(new_n685), .B(new_n687), .C1(new_n684), .C2(new_n682), .ZN(new_n688));
  MUX2_X1   g263(.A(G6), .B(G305), .S(G16), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT32), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n690), .A2(G1981), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(G1981), .ZN(new_n692));
  INV_X1    g267(.A(G16), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G23), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(new_n569), .B2(new_n693), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT33), .B(G1976), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n693), .A2(G22), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G166), .B2(new_n693), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n700), .A2(G1971), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  AOI22_X1  g277(.A1(new_n695), .A2(new_n697), .B1(new_n700), .B2(G1971), .ZN(new_n703));
  NAND4_X1  g278(.A1(new_n691), .A2(new_n692), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n704), .A2(KEYINPUT34), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(KEYINPUT34), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n688), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT36), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT100), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n674), .A2(G35), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G162), .B2(new_n674), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT29), .B(G2090), .Z(new_n712));
  XOR2_X1   g287(.A(new_n711), .B(new_n712), .Z(new_n713));
  NOR2_X1   g288(.A1(G164), .A2(new_n674), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(G27), .B2(new_n674), .ZN(new_n715));
  INV_X1    g290(.A(G2078), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n693), .A2(G20), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT99), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT23), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G299), .B2(G16), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G1956), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n715), .A2(new_n716), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n674), .B1(KEYINPUT24), .B2(G34), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(KEYINPUT24), .B2(G34), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n482), .B2(G29), .ZN(new_n726));
  INV_X1    g301(.A(G2084), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g303(.A1(new_n717), .A2(new_n722), .A3(new_n723), .A4(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(G29), .A2(G33), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT89), .Z(new_n731));
  NAND3_X1  g306(.A1(new_n475), .A2(new_n477), .A3(G127), .ZN(new_n732));
  INV_X1    g307(.A(G115), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n733), .B2(new_n465), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G2105), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT25), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n736), .A2(new_n737), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n462), .A2(G139), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n735), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n731), .B1(new_n742), .B2(new_n674), .ZN(new_n743));
  INV_X1    g318(.A(G2072), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n693), .A2(G21), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G168), .B2(new_n693), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n743), .A2(new_n744), .B1(new_n746), .B2(G1966), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n674), .A2(G26), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT28), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n492), .A2(G128), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n462), .A2(G140), .ZN(new_n751));
  OR2_X1    g326(.A1(G104), .A2(G2105), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n752), .B(G2104), .C1(G116), .C2(new_n469), .ZN(new_n753));
  AND3_X1   g328(.A1(new_n750), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n749), .B1(new_n754), .B2(new_n674), .ZN(new_n755));
  INV_X1    g330(.A(G2067), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n693), .A2(G19), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n546), .B2(new_n693), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT88), .B(G1341), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n693), .A2(G5), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G171), .B2(new_n693), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(G1961), .Z(new_n764));
  NAND4_X1  g339(.A1(new_n747), .A2(new_n757), .A3(new_n761), .A4(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n726), .A2(new_n727), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT90), .Z(new_n767));
  NOR4_X1   g342(.A1(new_n713), .A2(new_n729), .A3(new_n765), .A4(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n746), .A2(G1966), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT98), .Z(new_n770));
  NAND2_X1  g345(.A1(new_n693), .A2(G4), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n595), .B2(new_n693), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G1348), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n743), .A2(new_n744), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT91), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT31), .B(G11), .Z(new_n777));
  INV_X1    g352(.A(KEYINPUT30), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n674), .B1(new_n778), .B2(G28), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT96), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI22_X1  g356(.A1(new_n779), .A2(new_n780), .B1(new_n778), .B2(G28), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n777), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(new_n612), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(new_n674), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT97), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n768), .A2(new_n774), .A3(new_n776), .A4(new_n786), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n468), .A2(G141), .A3(new_n469), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n473), .A2(G105), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g365(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n791), .A2(KEYINPUT93), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(KEYINPUT93), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n794), .A2(KEYINPUT26), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT26), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n792), .A2(new_n796), .A3(new_n793), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n790), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT92), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(new_n492), .B2(G129), .ZN(new_n800));
  INV_X1    g375(.A(G129), .ZN(new_n801));
  AOI211_X1 g376(.A(KEYINPUT92), .B(new_n801), .C1(new_n489), .C2(new_n491), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n798), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT94), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n805), .A2(new_n674), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n674), .B2(G32), .ZN(new_n807));
  INV_X1    g382(.A(G1996), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT95), .B(KEYINPUT27), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n807), .A2(new_n808), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n809), .A2(new_n811), .ZN(new_n813));
  INV_X1    g388(.A(new_n810), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n787), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  AND3_X1   g391(.A1(new_n708), .A2(new_n709), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n709), .B1(new_n708), .B2(new_n816), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n817), .A2(new_n818), .ZN(G311));
  NAND2_X1  g394(.A1(new_n708), .A2(new_n816), .ZN(G150));
  AOI22_X1  g395(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n821), .A2(new_n515), .ZN(new_n822));
  INV_X1    g397(.A(G93), .ZN(new_n823));
  INV_X1    g398(.A(G55), .ZN(new_n824));
  OAI22_X1  g399(.A1(new_n518), .A2(new_n823), .B1(new_n520), .B2(new_n824), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT101), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OR3_X1    g403(.A1(new_n822), .A2(new_n825), .A3(new_n827), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n828), .A2(new_n546), .A3(new_n829), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n826), .B(new_n827), .C1(new_n542), .C2(new_n545), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT38), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n595), .A2(G559), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT39), .ZN(new_n836));
  AOI21_X1  g411(.A(G860), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n836), .B2(new_n835), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT102), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n826), .A2(G860), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT37), .Z(new_n841));
  NAND2_X1  g416(.A1(new_n839), .A2(new_n841), .ZN(G145));
  XNOR2_X1  g417(.A(new_n612), .B(G160), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(G162), .Z(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n462), .A2(G142), .ZN(new_n846));
  NOR2_X1   g421(.A1(G106), .A2(G2105), .ZN(new_n847));
  OAI21_X1  g422(.A(G2104), .B1(new_n469), .B2(G118), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n849), .B1(G130), .B2(new_n492), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n803), .A2(new_n754), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n750), .A2(new_n751), .A3(new_n753), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n852), .B(new_n798), .C1(new_n800), .C2(new_n802), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT104), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT103), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n502), .B1(new_n508), .B2(new_n856), .ZN(new_n857));
  AOI211_X1 g432(.A(KEYINPUT103), .B(new_n504), .C1(new_n506), .C2(new_n507), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n855), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n506), .A2(new_n507), .ZN(new_n860));
  INV_X1    g435(.A(new_n504), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(KEYINPUT103), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n508), .A2(new_n856), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n863), .A2(KEYINPUT104), .A3(new_n502), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n859), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n854), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n851), .A2(new_n859), .A3(new_n853), .A4(new_n865), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n741), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  AND4_X1   g445(.A1(new_n859), .A2(new_n851), .A3(new_n865), .A4(new_n853), .ZN(new_n871));
  AOI22_X1  g446(.A1(new_n851), .A2(new_n853), .B1(new_n859), .B2(new_n865), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n804), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n867), .A2(KEYINPUT94), .A3(new_n868), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n742), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT105), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n870), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI211_X1 g452(.A(KEYINPUT105), .B(new_n742), .C1(new_n873), .C2(new_n874), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n850), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n681), .B(KEYINPUT106), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n880), .B(new_n615), .Z(new_n881));
  AND3_X1   g456(.A1(new_n867), .A2(KEYINPUT94), .A3(new_n868), .ZN(new_n882));
  AOI21_X1  g457(.A(KEYINPUT94), .B1(new_n867), .B2(new_n868), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n741), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(KEYINPUT105), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n875), .A2(new_n876), .ZN(new_n886));
  INV_X1    g461(.A(new_n850), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n885), .A2(new_n886), .A3(new_n887), .A4(new_n870), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n879), .A2(new_n881), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n881), .B1(new_n879), .B2(new_n888), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n845), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n881), .ZN(new_n892));
  NOR3_X1   g467(.A1(new_n877), .A2(new_n850), .A3(new_n878), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n869), .B1(new_n884), .B2(KEYINPUT105), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n887), .B1(new_n894), .B2(new_n886), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n892), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n879), .A2(new_n881), .A3(new_n888), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(new_n844), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(G37), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n891), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT40), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n891), .A2(new_n898), .A3(KEYINPUT40), .A4(new_n899), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(G395));
  INV_X1    g479(.A(G868), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n826), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n595), .A2(G299), .ZN(new_n907));
  INV_X1    g482(.A(G299), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n594), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT41), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n907), .A2(new_n909), .A3(KEYINPUT41), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n832), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(new_n603), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  XOR2_X1   g492(.A(new_n917), .B(KEYINPUT107), .Z(new_n918));
  INV_X1    g493(.A(new_n910), .ZN(new_n919));
  OR2_X1    g494(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  XOR2_X1   g495(.A(G290), .B(G166), .Z(new_n921));
  XNOR2_X1  g496(.A(new_n569), .B(G305), .ZN(new_n922));
  XOR2_X1   g497(.A(new_n921), .B(new_n922), .Z(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(KEYINPUT42), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n918), .B(new_n920), .C1(new_n924), .C2(KEYINPUT108), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n924), .A2(KEYINPUT108), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n925), .B(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n906), .B1(new_n927), .B2(new_n905), .ZN(G295));
  OAI21_X1  g503(.A(new_n906), .B1(new_n927), .B2(new_n905), .ZN(G331));
  NAND2_X1  g504(.A1(G286), .A2(KEYINPUT109), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT109), .ZN(new_n931));
  AOI21_X1  g506(.A(G301), .B1(G168), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(G286), .A2(KEYINPUT109), .A3(G301), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n933), .A2(new_n915), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n915), .B1(new_n933), .B2(new_n934), .ZN(new_n937));
  NOR3_X1   g512(.A1(new_n936), .A2(new_n937), .A3(new_n919), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n933), .A2(new_n934), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n832), .ZN(new_n940));
  AOI22_X1  g515(.A1(new_n940), .A2(new_n935), .B1(new_n912), .B2(new_n913), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n921), .B(new_n922), .ZN(new_n942));
  NOR3_X1   g517(.A1(new_n938), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n942), .B1(new_n941), .B2(new_n938), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n899), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT110), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n944), .A2(KEYINPUT110), .A3(new_n899), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT43), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n941), .ZN(new_n950));
  INV_X1    g525(.A(new_n938), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(new_n951), .A3(new_n923), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n899), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n912), .A2(KEYINPUT111), .A3(new_n913), .ZN(new_n954));
  OAI221_X1 g529(.A(new_n954), .B1(KEYINPUT111), .B2(new_n912), .C1(new_n936), .C2(new_n937), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n923), .B1(new_n955), .B2(new_n951), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n953), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT44), .B1(new_n949), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n957), .B1(new_n947), .B2(new_n948), .ZN(new_n960));
  NOR3_X1   g535(.A1(new_n953), .A2(new_n956), .A3(KEYINPUT43), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n959), .B1(new_n962), .B2(KEYINPUT44), .ZN(G397));
  XNOR2_X1  g538(.A(KEYINPUT123), .B(G1961), .ZN(new_n964));
  INV_X1    g539(.A(G1384), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n509), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n965), .B1(new_n857), .B2(new_n858), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n968), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n474), .A2(G40), .A3(new_n481), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n964), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT125), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT53), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n975), .A2(G1384), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n859), .A2(new_n865), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n971), .B1(new_n975), .B2(new_n966), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n974), .B1(new_n979), .B2(G2078), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n975), .B1(new_n866), .B2(G1384), .ZN(new_n981));
  XOR2_X1   g556(.A(new_n474), .B(KEYINPUT126), .Z(new_n982));
  NOR2_X1   g557(.A1(new_n974), .A2(G2078), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n481), .A2(G40), .A3(new_n983), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n981), .A2(new_n977), .A3(new_n982), .A4(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n971), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n863), .A2(new_n502), .A3(new_n864), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT50), .B1(new_n987), .B2(new_n965), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n986), .B1(new_n988), .B2(new_n968), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT125), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n989), .A2(new_n990), .A3(new_n964), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n973), .A2(new_n980), .A3(new_n985), .A4(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT127), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n992), .A2(new_n993), .A3(G171), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n993), .B1(new_n992), .B2(G171), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT54), .ZN(new_n997));
  INV_X1    g572(.A(new_n980), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT116), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n509), .A2(new_n999), .A3(new_n976), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n999), .B1(new_n509), .B2(new_n976), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n986), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT45), .B1(new_n987), .B2(new_n965), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n983), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n972), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT124), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT124), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(new_n972), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n998), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n997), .B1(new_n1010), .B2(G301), .ZN(new_n1011));
  INV_X1    g586(.A(G1348), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n989), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n986), .A2(new_n987), .A3(new_n965), .ZN(new_n1014));
  OR2_X1    g589(.A1(new_n1014), .A2(G2067), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1013), .A2(new_n594), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n594), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT60), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AND2_X1   g593(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT60), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1019), .A2(new_n1020), .A3(new_n595), .ZN(new_n1021));
  XOR2_X1   g596(.A(KEYINPUT58), .B(G1341), .Z(new_n1022));
  NAND2_X1  g597(.A1(new_n1014), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(new_n979), .B2(G1996), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n546), .ZN(new_n1025));
  AND2_X1   g600(.A1(new_n1025), .A2(KEYINPUT59), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1025), .A2(KEYINPUT59), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1018), .B(new_n1021), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  XOR2_X1   g603(.A(G299), .B(KEYINPUT57), .Z(new_n1029));
  XNOR2_X1  g604(.A(KEYINPUT56), .B(G2072), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n977), .A2(new_n978), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT120), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n1031), .B(new_n1032), .ZN(new_n1033));
  XOR2_X1   g608(.A(KEYINPUT118), .B(G1956), .Z(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n986), .B1(KEYINPUT50), .B2(new_n966), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n967), .B1(new_n987), .B2(new_n965), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1035), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT119), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT119), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1040), .B(new_n1035), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1029), .B1(new_n1033), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1033), .A2(new_n1042), .A3(new_n1029), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1043), .B1(new_n1044), .B2(new_n1017), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n996), .A2(new_n1011), .B1(new_n1028), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT51), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n727), .B(new_n986), .C1(new_n988), .C2(new_n968), .ZN(new_n1048));
  INV_X1    g623(.A(G1966), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1049), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1048), .A2(new_n1050), .A3(G168), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1047), .B1(new_n1051), .B2(G8), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(G168), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1054));
  OAI211_X1 g629(.A(G8), .B(new_n1051), .C1(new_n1054), .C2(new_n1047), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT122), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n561), .A2(G8), .A3(new_n562), .ZN(new_n1059));
  XOR2_X1   g634(.A(new_n1059), .B(KEYINPUT55), .Z(new_n1060));
  AOI21_X1  g635(.A(G1971), .B1(new_n977), .B2(new_n978), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(G2090), .B2(new_n989), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1065));
  OAI211_X1 g640(.A(G8), .B(new_n1060), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT61), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1033), .A2(new_n1042), .A3(new_n1067), .A4(new_n1029), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1060), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n1036), .A2(new_n1037), .A3(G2090), .ZN(new_n1070));
  OAI21_X1  g645(.A(G8), .B1(new_n1070), .B2(new_n1061), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT115), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1014), .A2(G8), .ZN(new_n1074));
  NAND2_X1  g649(.A1(G305), .A2(G1981), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n574), .A2(new_n575), .A3(new_n576), .A4(new_n666), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1075), .A2(KEYINPUT49), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT49), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1073), .B1(new_n1074), .B2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1014), .A2(new_n1079), .A3(KEYINPUT115), .A4(G8), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n569), .A2(G1976), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1014), .A2(G8), .A3(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n569), .A2(G1976), .ZN(new_n1086));
  OR3_X1    g661(.A1(new_n1085), .A2(KEYINPUT52), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1085), .A2(KEYINPUT52), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1083), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1066), .A2(new_n1068), .A3(new_n1072), .A4(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1056), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n1058), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n985), .A2(new_n980), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1093), .A2(G301), .A3(new_n973), .A4(new_n991), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1094), .B1(new_n1010), .B2(G301), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1067), .A2(KEYINPUT121), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n1019), .B2(new_n594), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1043), .B1(new_n1097), .B2(new_n1044), .ZN(new_n1098));
  OR2_X1    g673(.A1(new_n1044), .A2(KEYINPUT121), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1095), .A2(new_n997), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1046), .A2(new_n1092), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1102), .A2(G8), .A3(G168), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1066), .A2(KEYINPUT63), .A3(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(G8), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n1069), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT117), .B1(new_n1106), .B2(new_n1089), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT117), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1083), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1109));
  AOI211_X1 g684(.A(new_n1108), .B(new_n1109), .C1(new_n1105), .C2(new_n1069), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1104), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT63), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1066), .A2(new_n1072), .A3(new_n1089), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1103), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1112), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1111), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1117), .B1(new_n1058), .B2(new_n1091), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1091), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1119), .A2(KEYINPUT62), .A3(new_n1057), .ZN(new_n1120));
  NOR3_X1   g695(.A1(new_n1113), .A2(G301), .A3(new_n1010), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1118), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1066), .A2(new_n1109), .ZN(new_n1123));
  INV_X1    g698(.A(G1976), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1083), .A2(new_n1124), .A3(new_n569), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1074), .B1(new_n1125), .B2(new_n1076), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1101), .A2(new_n1116), .A3(new_n1122), .A4(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n981), .A2(new_n971), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n808), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1130), .B(KEYINPUT112), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n805), .ZN(new_n1132));
  INV_X1    g707(.A(new_n684), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n681), .B(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1129), .A2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n852), .B(new_n756), .ZN(new_n1136));
  INV_X1    g711(.A(new_n803), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1136), .B1(new_n1137), .B2(new_n808), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1129), .A2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(G290), .A2(G1986), .ZN(new_n1140));
  AND2_X1   g715(.A1(G290), .A2(G1986), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1129), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1132), .A2(new_n1135), .A3(new_n1139), .A4(new_n1142), .ZN(new_n1143));
  XOR2_X1   g718(.A(new_n1143), .B(KEYINPUT113), .Z(new_n1144));
  NAND2_X1  g719(.A1(new_n1128), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1129), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1146), .B1(new_n1137), .B2(new_n1136), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT46), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1131), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT112), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1130), .B(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(KEYINPUT46), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1147), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT47), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  AOI211_X1 g730(.A(KEYINPUT47), .B(new_n1147), .C1(new_n1149), .C2(new_n1152), .ZN(new_n1156));
  AND2_X1   g731(.A1(new_n1132), .A2(new_n1139), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(new_n1135), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1129), .A2(new_n1140), .ZN(new_n1159));
  XOR2_X1   g734(.A(new_n1159), .B(KEYINPUT48), .Z(new_n1160));
  OAI22_X1  g735(.A1(new_n1155), .A2(new_n1156), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1157), .A2(new_n1133), .A3(new_n681), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n754), .A2(new_n756), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1146), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1145), .A2(new_n1165), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g741(.A1(new_n635), .A2(G319), .ZN(new_n1168));
  NOR3_X1   g742(.A1(G229), .A2(G227), .A3(new_n1168), .ZN(new_n1169));
  OAI211_X1 g743(.A(new_n900), .B(new_n1169), .C1(new_n960), .C2(new_n961), .ZN(G225));
  INV_X1    g744(.A(G225), .ZN(G308));
endmodule


