

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U553 ( .A1(G2104), .A2(G2105), .ZN(n903) );
  NAND2_X1 U554 ( .A1(G8), .A2(n726), .ZN(n745) );
  NAND2_X2 U555 ( .A1(n781), .A2(n693), .ZN(n726) );
  NOR2_X2 U556 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  AND2_X1 U557 ( .A1(n729), .A2(n728), .ZN(n740) );
  XNOR2_X1 U558 ( .A(n587), .B(KEYINPUT15), .ZN(n994) );
  INV_X2 U559 ( .A(n726), .ZN(n700) );
  NOR2_X2 U560 ( .A1(n653), .A2(G651), .ZN(n522) );
  AND2_X2 U561 ( .A1(n529), .A2(G2104), .ZN(n907) );
  XNOR2_X1 U562 ( .A(n539), .B(G543), .ZN(n653) );
  NOR2_X2 U563 ( .A1(G2104), .A2(n529), .ZN(n556) );
  XNOR2_X1 U564 ( .A(n707), .B(n706), .ZN(n708) );
  NAND2_X1 U565 ( .A1(n738), .A2(n519), .ZN(n743) );
  NAND2_X1 U566 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U567 ( .A(KEYINPUT23), .B(KEYINPUT65), .ZN(n523) );
  NAND2_X1 U568 ( .A1(G171), .A2(n734), .ZN(n518) );
  XOR2_X1 U569 ( .A(n737), .B(KEYINPUT31), .Z(n519) );
  XOR2_X1 U570 ( .A(n720), .B(KEYINPUT29), .Z(n520) );
  NOR2_X1 U571 ( .A1(n765), .A2(n764), .ZN(n521) );
  NOR2_X2 U572 ( .A1(n563), .A2(n562), .ZN(G164) );
  INV_X1 U573 ( .A(KEYINPUT27), .ZN(n706) );
  INV_X1 U574 ( .A(KEYINPUT105), .ZN(n730) );
  XNOR2_X1 U575 ( .A(n740), .B(n730), .ZN(n731) );
  NAND2_X1 U576 ( .A1(n520), .A2(n518), .ZN(n738) );
  OR2_X1 U577 ( .A1(n761), .A2(KEYINPUT33), .ZN(n766) );
  INV_X1 U578 ( .A(KEYINPUT72), .ZN(n580) );
  NOR2_X1 U579 ( .A1(G164), .A2(G1384), .ZN(n781) );
  XNOR2_X1 U580 ( .A(n581), .B(n580), .ZN(n582) );
  INV_X1 U581 ( .A(KEYINPUT17), .ZN(n525) );
  INV_X1 U582 ( .A(KEYINPUT0), .ZN(n539) );
  XNOR2_X1 U583 ( .A(n526), .B(n525), .ZN(n552) );
  NOR2_X1 U584 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U585 ( .A1(n552), .A2(G138), .ZN(n553) );
  INV_X1 U586 ( .A(KEYINPUT87), .ZN(n560) );
  XNOR2_X1 U587 ( .A(n524), .B(n523), .ZN(n528) );
  INV_X1 U588 ( .A(G2105), .ZN(n529) );
  NAND2_X1 U589 ( .A1(G101), .A2(n907), .ZN(n524) );
  BUF_X2 U590 ( .A(n552), .Z(n908) );
  NAND2_X1 U591 ( .A1(G137), .A2(n908), .ZN(n527) );
  NAND2_X1 U592 ( .A1(n528), .A2(n527), .ZN(n533) );
  NAND2_X1 U593 ( .A1(G113), .A2(n903), .ZN(n531) );
  BUF_X1 U594 ( .A(n556), .Z(n904) );
  NAND2_X1 U595 ( .A1(G125), .A2(n904), .ZN(n530) );
  NAND2_X1 U596 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X2 U597 ( .A1(n533), .A2(n532), .ZN(G160) );
  INV_X1 U598 ( .A(G651), .ZN(n540) );
  NOR2_X1 U599 ( .A1(G543), .A2(n540), .ZN(n535) );
  XNOR2_X1 U600 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(n658) );
  NAND2_X1 U602 ( .A1(G65), .A2(n658), .ZN(n538) );
  NOR2_X1 U603 ( .A1(G651), .A2(G543), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n536), .B(KEYINPUT64), .ZN(n645) );
  NAND2_X1 U605 ( .A1(G91), .A2(n645), .ZN(n537) );
  NAND2_X1 U606 ( .A1(n538), .A2(n537), .ZN(n544) );
  NOR2_X1 U607 ( .A1(n653), .A2(n540), .ZN(n644) );
  NAND2_X1 U608 ( .A1(G78), .A2(n644), .ZN(n542) );
  NAND2_X1 U609 ( .A1(G53), .A2(n522), .ZN(n541) );
  NAND2_X1 U610 ( .A1(n542), .A2(n541), .ZN(n543) );
  OR2_X1 U611 ( .A1(n544), .A2(n543), .ZN(G299) );
  NAND2_X1 U612 ( .A1(G64), .A2(n658), .ZN(n546) );
  NAND2_X1 U613 ( .A1(G52), .A2(n522), .ZN(n545) );
  NAND2_X1 U614 ( .A1(n546), .A2(n545), .ZN(n551) );
  NAND2_X1 U615 ( .A1(G77), .A2(n644), .ZN(n548) );
  NAND2_X1 U616 ( .A1(G90), .A2(n645), .ZN(n547) );
  NAND2_X1 U617 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U618 ( .A(KEYINPUT9), .B(n549), .Z(n550) );
  NOR2_X1 U619 ( .A1(n551), .A2(n550), .ZN(G171) );
  INV_X1 U620 ( .A(G171), .ZN(G301) );
  AND2_X1 U621 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U622 ( .A(G57), .ZN(G237) );
  INV_X1 U623 ( .A(G108), .ZN(G238) );
  INV_X1 U624 ( .A(G132), .ZN(G219) );
  INV_X1 U625 ( .A(G82), .ZN(G220) );
  NAND2_X1 U626 ( .A1(G102), .A2(n907), .ZN(n554) );
  NAND2_X1 U627 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U628 ( .A(n555), .B(KEYINPUT88), .ZN(n563) );
  NAND2_X1 U629 ( .A1(n556), .A2(G126), .ZN(n557) );
  XNOR2_X1 U630 ( .A(n557), .B(KEYINPUT86), .ZN(n559) );
  NAND2_X1 U631 ( .A1(G114), .A2(n903), .ZN(n558) );
  NAND2_X1 U632 ( .A1(n559), .A2(n558), .ZN(n561) );
  XNOR2_X1 U633 ( .A(n561), .B(n560), .ZN(n562) );
  NAND2_X1 U634 ( .A1(G7), .A2(G661), .ZN(n564) );
  XNOR2_X1 U635 ( .A(n564), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U636 ( .A(G567), .ZN(n688) );
  NOR2_X1 U637 ( .A1(G223), .A2(n688), .ZN(n566) );
  XNOR2_X1 U638 ( .A(KEYINPUT68), .B(KEYINPUT11), .ZN(n565) );
  XNOR2_X1 U639 ( .A(n566), .B(n565), .ZN(G234) );
  NAND2_X1 U640 ( .A1(G56), .A2(n658), .ZN(n567) );
  XOR2_X1 U641 ( .A(KEYINPUT14), .B(n567), .Z(n573) );
  NAND2_X1 U642 ( .A1(G81), .A2(n645), .ZN(n568) );
  XNOR2_X1 U643 ( .A(n568), .B(KEYINPUT12), .ZN(n570) );
  NAND2_X1 U644 ( .A1(G68), .A2(n644), .ZN(n569) );
  NAND2_X1 U645 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U646 ( .A(KEYINPUT13), .B(n571), .Z(n572) );
  NOR2_X1 U647 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U648 ( .A1(n522), .A2(G43), .ZN(n574) );
  NAND2_X1 U649 ( .A1(n575), .A2(n574), .ZN(n979) );
  INV_X1 U650 ( .A(G860), .ZN(n602) );
  OR2_X1 U651 ( .A1(n979), .A2(n602), .ZN(G153) );
  NAND2_X1 U652 ( .A1(G868), .A2(G301), .ZN(n589) );
  NAND2_X1 U653 ( .A1(n645), .A2(G92), .ZN(n576) );
  XNOR2_X1 U654 ( .A(n576), .B(KEYINPUT70), .ZN(n583) );
  NAND2_X1 U655 ( .A1(n522), .A2(G54), .ZN(n577) );
  XOR2_X1 U656 ( .A(KEYINPUT71), .B(n577), .Z(n579) );
  NAND2_X1 U657 ( .A1(n644), .A2(G79), .ZN(n578) );
  NAND2_X1 U658 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U659 ( .A1(G66), .A2(n658), .ZN(n584) );
  XNOR2_X1 U660 ( .A(KEYINPUT69), .B(n584), .ZN(n585) );
  INV_X1 U661 ( .A(G868), .ZN(n671) );
  NAND2_X1 U662 ( .A1(n994), .A2(n671), .ZN(n588) );
  NAND2_X1 U663 ( .A1(n589), .A2(n588), .ZN(G284) );
  NAND2_X1 U664 ( .A1(G89), .A2(n645), .ZN(n590) );
  XNOR2_X1 U665 ( .A(n590), .B(KEYINPUT4), .ZN(n592) );
  NAND2_X1 U666 ( .A1(G76), .A2(n644), .ZN(n591) );
  NAND2_X1 U667 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U668 ( .A(n593), .B(KEYINPUT5), .ZN(n598) );
  NAND2_X1 U669 ( .A1(G63), .A2(n658), .ZN(n595) );
  NAND2_X1 U670 ( .A1(G51), .A2(n522), .ZN(n594) );
  NAND2_X1 U671 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U672 ( .A(KEYINPUT6), .B(n596), .Z(n597) );
  NAND2_X1 U673 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U674 ( .A(n599), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U675 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U676 ( .A1(G286), .A2(n671), .ZN(n601) );
  NOR2_X1 U677 ( .A1(G868), .A2(G299), .ZN(n600) );
  NOR2_X1 U678 ( .A1(n601), .A2(n600), .ZN(G297) );
  NAND2_X1 U679 ( .A1(n602), .A2(G559), .ZN(n603) );
  INV_X1 U680 ( .A(n994), .ZN(n618) );
  NAND2_X1 U681 ( .A1(n603), .A2(n618), .ZN(n604) );
  XNOR2_X1 U682 ( .A(n604), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U683 ( .A1(G868), .A2(n979), .ZN(n607) );
  NAND2_X1 U684 ( .A1(G868), .A2(n618), .ZN(n605) );
  NOR2_X1 U685 ( .A1(G559), .A2(n605), .ZN(n606) );
  NOR2_X1 U686 ( .A1(n607), .A2(n606), .ZN(G282) );
  NAND2_X1 U687 ( .A1(G123), .A2(n904), .ZN(n608) );
  XOR2_X1 U688 ( .A(KEYINPUT73), .B(n608), .Z(n609) );
  XNOR2_X1 U689 ( .A(n609), .B(KEYINPUT18), .ZN(n611) );
  NAND2_X1 U690 ( .A1(G111), .A2(n903), .ZN(n610) );
  NAND2_X1 U691 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U692 ( .A1(G99), .A2(n907), .ZN(n613) );
  NAND2_X1 U693 ( .A1(G135), .A2(n908), .ZN(n612) );
  NAND2_X1 U694 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U695 ( .A1(n615), .A2(n614), .ZN(n934) );
  XNOR2_X1 U696 ( .A(n934), .B(G2096), .ZN(n617) );
  INV_X1 U697 ( .A(G2100), .ZN(n616) );
  NAND2_X1 U698 ( .A1(n617), .A2(n616), .ZN(G156) );
  XNOR2_X1 U699 ( .A(KEYINPUT74), .B(n979), .ZN(n619) );
  NAND2_X1 U700 ( .A1(n618), .A2(G559), .ZN(n669) );
  XNOR2_X1 U701 ( .A(n619), .B(n669), .ZN(n620) );
  NOR2_X1 U702 ( .A1(G860), .A2(n620), .ZN(n629) );
  NAND2_X1 U703 ( .A1(G67), .A2(n658), .ZN(n621) );
  XNOR2_X1 U704 ( .A(n621), .B(KEYINPUT76), .ZN(n628) );
  NAND2_X1 U705 ( .A1(n522), .A2(G55), .ZN(n623) );
  NAND2_X1 U706 ( .A1(G93), .A2(n645), .ZN(n622) );
  NAND2_X1 U707 ( .A1(n623), .A2(n622), .ZN(n626) );
  NAND2_X1 U708 ( .A1(G80), .A2(n644), .ZN(n624) );
  XNOR2_X1 U709 ( .A(KEYINPUT75), .B(n624), .ZN(n625) );
  NOR2_X1 U710 ( .A1(n626), .A2(n625), .ZN(n627) );
  NAND2_X1 U711 ( .A1(n628), .A2(n627), .ZN(n672) );
  XOR2_X1 U712 ( .A(n629), .B(n672), .Z(G145) );
  NAND2_X1 U713 ( .A1(n522), .A2(G47), .ZN(n631) );
  NAND2_X1 U714 ( .A1(G85), .A2(n645), .ZN(n630) );
  NAND2_X1 U715 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U716 ( .A1(G72), .A2(n644), .ZN(n632) );
  XOR2_X1 U717 ( .A(KEYINPUT66), .B(n632), .Z(n633) );
  NOR2_X1 U718 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U719 ( .A1(n658), .A2(G60), .ZN(n635) );
  NAND2_X1 U720 ( .A1(n636), .A2(n635), .ZN(G290) );
  NAND2_X1 U721 ( .A1(G61), .A2(n658), .ZN(n638) );
  NAND2_X1 U722 ( .A1(G86), .A2(n645), .ZN(n637) );
  NAND2_X1 U723 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U724 ( .A1(n644), .A2(G73), .ZN(n639) );
  XOR2_X1 U725 ( .A(KEYINPUT2), .B(n639), .Z(n640) );
  NOR2_X1 U726 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U727 ( .A1(n522), .A2(G48), .ZN(n642) );
  NAND2_X1 U728 ( .A1(n643), .A2(n642), .ZN(G305) );
  NAND2_X1 U729 ( .A1(G75), .A2(n644), .ZN(n647) );
  NAND2_X1 U730 ( .A1(G88), .A2(n645), .ZN(n646) );
  NAND2_X1 U731 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U732 ( .A(KEYINPUT79), .B(n648), .ZN(n652) );
  NAND2_X1 U733 ( .A1(G62), .A2(n658), .ZN(n650) );
  NAND2_X1 U734 ( .A1(G50), .A2(n522), .ZN(n649) );
  AND2_X1 U735 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U736 ( .A1(n652), .A2(n651), .ZN(G303) );
  INV_X1 U737 ( .A(G303), .ZN(G166) );
  NAND2_X1 U738 ( .A1(n653), .A2(G87), .ZN(n654) );
  XNOR2_X1 U739 ( .A(KEYINPUT78), .B(n654), .ZN(n661) );
  NAND2_X1 U740 ( .A1(G49), .A2(n522), .ZN(n656) );
  NAND2_X1 U741 ( .A1(G74), .A2(G651), .ZN(n655) );
  NAND2_X1 U742 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U743 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U744 ( .A(KEYINPUT77), .B(n659), .Z(n660) );
  NAND2_X1 U745 ( .A1(n661), .A2(n660), .ZN(G288) );
  XNOR2_X1 U746 ( .A(G290), .B(G305), .ZN(n668) );
  XOR2_X1 U747 ( .A(KEYINPUT19), .B(KEYINPUT80), .Z(n662) );
  XNOR2_X1 U748 ( .A(G288), .B(n662), .ZN(n663) );
  XNOR2_X1 U749 ( .A(n663), .B(n979), .ZN(n664) );
  XNOR2_X1 U750 ( .A(n664), .B(G299), .ZN(n665) );
  XNOR2_X1 U751 ( .A(G166), .B(n665), .ZN(n666) );
  XNOR2_X1 U752 ( .A(n666), .B(n672), .ZN(n667) );
  XNOR2_X1 U753 ( .A(n668), .B(n667), .ZN(n854) );
  XOR2_X1 U754 ( .A(n854), .B(n669), .Z(n670) );
  NOR2_X1 U755 ( .A1(n671), .A2(n670), .ZN(n674) );
  NOR2_X1 U756 ( .A1(G868), .A2(n672), .ZN(n673) );
  NOR2_X1 U757 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U758 ( .A(KEYINPUT81), .B(n675), .Z(G295) );
  NAND2_X1 U759 ( .A1(G2078), .A2(G2084), .ZN(n676) );
  XOR2_X1 U760 ( .A(KEYINPUT20), .B(n676), .Z(n677) );
  NAND2_X1 U761 ( .A1(G2090), .A2(n677), .ZN(n678) );
  XNOR2_X1 U762 ( .A(KEYINPUT21), .B(n678), .ZN(n679) );
  NAND2_X1 U763 ( .A1(n679), .A2(G2072), .ZN(n680) );
  XNOR2_X1 U764 ( .A(KEYINPUT82), .B(n680), .ZN(G158) );
  XNOR2_X1 U765 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U766 ( .A1(G220), .A2(G219), .ZN(n681) );
  XOR2_X1 U767 ( .A(KEYINPUT22), .B(n681), .Z(n682) );
  NOR2_X1 U768 ( .A1(G218), .A2(n682), .ZN(n683) );
  NAND2_X1 U769 ( .A1(G96), .A2(n683), .ZN(n840) );
  NAND2_X1 U770 ( .A1(G2106), .A2(n840), .ZN(n684) );
  XNOR2_X1 U771 ( .A(n684), .B(KEYINPUT83), .ZN(n690) );
  NAND2_X1 U772 ( .A1(G120), .A2(G69), .ZN(n685) );
  NOR2_X1 U773 ( .A1(G237), .A2(n685), .ZN(n686) );
  XOR2_X1 U774 ( .A(KEYINPUT84), .B(n686), .Z(n687) );
  NOR2_X1 U775 ( .A1(G238), .A2(n687), .ZN(n842) );
  NOR2_X1 U776 ( .A1(n688), .A2(n842), .ZN(n689) );
  NOR2_X1 U777 ( .A1(n690), .A2(n689), .ZN(G319) );
  INV_X1 U778 ( .A(G319), .ZN(n919) );
  NAND2_X1 U779 ( .A1(G661), .A2(G483), .ZN(n691) );
  XOR2_X1 U780 ( .A(KEYINPUT85), .B(n691), .Z(n692) );
  NOR2_X1 U781 ( .A1(n919), .A2(n692), .ZN(n837) );
  NAND2_X1 U782 ( .A1(n837), .A2(G36), .ZN(G176) );
  NAND2_X1 U783 ( .A1(G160), .A2(G40), .ZN(n782) );
  INV_X1 U784 ( .A(n782), .ZN(n693) );
  XNOR2_X1 U785 ( .A(G1996), .B(KEYINPUT102), .ZN(n957) );
  NAND2_X1 U786 ( .A1(n700), .A2(n957), .ZN(n694) );
  XNOR2_X1 U787 ( .A(n694), .B(KEYINPUT26), .ZN(n696) );
  INV_X1 U788 ( .A(n700), .ZN(n746) );
  NAND2_X1 U789 ( .A1(G1341), .A2(n746), .ZN(n695) );
  NAND2_X1 U790 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U791 ( .A(KEYINPUT103), .B(n697), .ZN(n698) );
  INV_X1 U792 ( .A(n698), .ZN(n699) );
  NOR2_X1 U793 ( .A1(n979), .A2(n699), .ZN(n704) );
  NAND2_X1 U794 ( .A1(G1348), .A2(n746), .ZN(n702) );
  NAND2_X1 U795 ( .A1(G2067), .A2(n700), .ZN(n701) );
  NAND2_X1 U796 ( .A1(n702), .A2(n701), .ZN(n710) );
  NAND2_X1 U797 ( .A1(n710), .A2(n994), .ZN(n703) );
  NAND2_X1 U798 ( .A1(n704), .A2(n703), .ZN(n714) );
  NAND2_X1 U799 ( .A1(G1956), .A2(n746), .ZN(n705) );
  XOR2_X1 U800 ( .A(KEYINPUT101), .B(n705), .Z(n709) );
  NAND2_X1 U801 ( .A1(n700), .A2(G2072), .ZN(n707) );
  NAND2_X1 U802 ( .A1(n709), .A2(n708), .ZN(n716) );
  NOR2_X1 U803 ( .A1(G299), .A2(n716), .ZN(n712) );
  NOR2_X1 U804 ( .A1(n710), .A2(n994), .ZN(n711) );
  NOR2_X1 U805 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U806 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U807 ( .A(n715), .B(KEYINPUT104), .ZN(n719) );
  NAND2_X1 U808 ( .A1(G299), .A2(n716), .ZN(n717) );
  XNOR2_X1 U809 ( .A(KEYINPUT28), .B(n717), .ZN(n718) );
  NAND2_X1 U810 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U811 ( .A(G1961), .B(KEYINPUT98), .ZN(n1007) );
  NAND2_X1 U812 ( .A1(n746), .A2(n1007), .ZN(n723) );
  XNOR2_X1 U813 ( .A(G2078), .B(KEYINPUT25), .ZN(n721) );
  XNOR2_X1 U814 ( .A(n721), .B(KEYINPUT99), .ZN(n958) );
  NAND2_X1 U815 ( .A1(n700), .A2(n958), .ZN(n722) );
  NAND2_X1 U816 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U817 ( .A(n724), .B(KEYINPUT100), .Z(n734) );
  NOR2_X1 U818 ( .A1(G1966), .A2(n745), .ZN(n725) );
  XNOR2_X1 U819 ( .A(n725), .B(KEYINPUT97), .ZN(n729) );
  NOR2_X1 U820 ( .A1(G2084), .A2(n726), .ZN(n727) );
  XOR2_X1 U821 ( .A(KEYINPUT96), .B(n727), .Z(n728) );
  NAND2_X1 U822 ( .A1(n731), .A2(G8), .ZN(n732) );
  XNOR2_X1 U823 ( .A(KEYINPUT30), .B(n732), .ZN(n733) );
  NOR2_X1 U824 ( .A1(G168), .A2(n733), .ZN(n736) );
  NOR2_X1 U825 ( .A1(G171), .A2(n734), .ZN(n735) );
  NOR2_X1 U826 ( .A1(n736), .A2(n735), .ZN(n737) );
  INV_X1 U827 ( .A(n743), .ZN(n742) );
  NOR2_X1 U828 ( .A1(G8), .A2(KEYINPUT97), .ZN(n739) );
  NOR2_X1 U829 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U830 ( .A1(n742), .A2(n741), .ZN(n756) );
  INV_X1 U831 ( .A(KEYINPUT32), .ZN(n754) );
  NAND2_X1 U832 ( .A1(n743), .A2(G286), .ZN(n744) );
  XNOR2_X1 U833 ( .A(n744), .B(KEYINPUT106), .ZN(n751) );
  NOR2_X1 U834 ( .A1(G1971), .A2(n745), .ZN(n748) );
  NOR2_X1 U835 ( .A1(G2090), .A2(n746), .ZN(n747) );
  NOR2_X1 U836 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U837 ( .A1(n749), .A2(G303), .ZN(n750) );
  NAND2_X1 U838 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U839 ( .A1(n752), .A2(G8), .ZN(n753) );
  XNOR2_X1 U840 ( .A(n754), .B(n753), .ZN(n755) );
  NOR2_X1 U841 ( .A1(n756), .A2(n755), .ZN(n773) );
  NOR2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n762) );
  INV_X1 U843 ( .A(n762), .ZN(n758) );
  INV_X1 U844 ( .A(G1971), .ZN(n1001) );
  NAND2_X1 U845 ( .A1(G166), .A2(n1001), .ZN(n757) );
  NAND2_X1 U846 ( .A1(n758), .A2(n757), .ZN(n991) );
  NOR2_X1 U847 ( .A1(n773), .A2(n991), .ZN(n760) );
  NAND2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n992) );
  INV_X1 U849 ( .A(n745), .ZN(n775) );
  NAND2_X1 U850 ( .A1(n992), .A2(n775), .ZN(n759) );
  NOR2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U852 ( .A(G1981), .B(G305), .Z(n984) );
  INV_X1 U853 ( .A(n984), .ZN(n765) );
  NAND2_X1 U854 ( .A1(n762), .A2(KEYINPUT33), .ZN(n763) );
  NOR2_X1 U855 ( .A1(n745), .A2(n763), .ZN(n764) );
  NAND2_X1 U856 ( .A1(n766), .A2(n521), .ZN(n779) );
  NOR2_X1 U857 ( .A1(G1981), .A2(G305), .ZN(n767) );
  XOR2_X1 U858 ( .A(n767), .B(KEYINPUT24), .Z(n768) );
  NOR2_X1 U859 ( .A1(n745), .A2(n768), .ZN(n777) );
  INV_X1 U860 ( .A(G8), .ZN(n771) );
  NOR2_X1 U861 ( .A1(G2090), .A2(G303), .ZN(n769) );
  XNOR2_X1 U862 ( .A(n769), .B(KEYINPUT107), .ZN(n770) );
  NOR2_X1 U863 ( .A1(n771), .A2(n770), .ZN(n772) );
  NOR2_X1 U864 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X1 U865 ( .A1(n775), .A2(n774), .ZN(n776) );
  NOR2_X1 U866 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U868 ( .A(n780), .B(KEYINPUT108), .ZN(n817) );
  NOR2_X1 U869 ( .A1(n781), .A2(n782), .ZN(n830) );
  XNOR2_X1 U870 ( .A(G1986), .B(G290), .ZN(n990) );
  AND2_X1 U871 ( .A1(n830), .A2(n990), .ZN(n815) );
  NAND2_X1 U872 ( .A1(G104), .A2(n907), .ZN(n784) );
  NAND2_X1 U873 ( .A1(G140), .A2(n908), .ZN(n783) );
  NAND2_X1 U874 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U875 ( .A(KEYINPUT34), .B(n785), .ZN(n790) );
  NAND2_X1 U876 ( .A1(G116), .A2(n903), .ZN(n787) );
  NAND2_X1 U877 ( .A1(G128), .A2(n904), .ZN(n786) );
  NAND2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n788) );
  XOR2_X1 U879 ( .A(KEYINPUT35), .B(n788), .Z(n789) );
  NOR2_X1 U880 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U881 ( .A(KEYINPUT36), .B(n791), .ZN(n884) );
  XNOR2_X1 U882 ( .A(G2067), .B(KEYINPUT37), .ZN(n828) );
  NOR2_X1 U883 ( .A1(n884), .A2(n828), .ZN(n927) );
  NAND2_X1 U884 ( .A1(n927), .A2(n830), .ZN(n792) );
  XOR2_X1 U885 ( .A(KEYINPUT89), .B(n792), .Z(n827) );
  NAND2_X1 U886 ( .A1(G117), .A2(n903), .ZN(n794) );
  NAND2_X1 U887 ( .A1(G129), .A2(n904), .ZN(n793) );
  NAND2_X1 U888 ( .A1(n794), .A2(n793), .ZN(n797) );
  NAND2_X1 U889 ( .A1(n908), .A2(G141), .ZN(n795) );
  XOR2_X1 U890 ( .A(KEYINPUT94), .B(n795), .Z(n796) );
  NOR2_X1 U891 ( .A1(n797), .A2(n796), .ZN(n801) );
  XOR2_X1 U892 ( .A(KEYINPUT93), .B(KEYINPUT38), .Z(n799) );
  NAND2_X1 U893 ( .A1(G105), .A2(n907), .ZN(n798) );
  XNOR2_X1 U894 ( .A(n799), .B(n798), .ZN(n800) );
  NAND2_X1 U895 ( .A1(n801), .A2(n800), .ZN(n802) );
  XOR2_X1 U896 ( .A(KEYINPUT95), .B(n802), .Z(n895) );
  NAND2_X1 U897 ( .A1(G1996), .A2(n895), .ZN(n813) );
  NAND2_X1 U898 ( .A1(G95), .A2(n907), .ZN(n803) );
  XOR2_X1 U899 ( .A(KEYINPUT92), .B(n803), .Z(n809) );
  NAND2_X1 U900 ( .A1(n904), .A2(G119), .ZN(n804) );
  XNOR2_X1 U901 ( .A(n804), .B(KEYINPUT90), .ZN(n806) );
  NAND2_X1 U902 ( .A1(G107), .A2(n903), .ZN(n805) );
  NAND2_X1 U903 ( .A1(n806), .A2(n805), .ZN(n807) );
  XOR2_X1 U904 ( .A(KEYINPUT91), .B(n807), .Z(n808) );
  NOR2_X1 U905 ( .A1(n809), .A2(n808), .ZN(n811) );
  NAND2_X1 U906 ( .A1(n908), .A2(G131), .ZN(n810) );
  NAND2_X1 U907 ( .A1(n811), .A2(n810), .ZN(n885) );
  NAND2_X1 U908 ( .A1(G1991), .A2(n885), .ZN(n812) );
  NAND2_X1 U909 ( .A1(n813), .A2(n812), .ZN(n929) );
  NAND2_X1 U910 ( .A1(n830), .A2(n929), .ZN(n819) );
  NAND2_X1 U911 ( .A1(n827), .A2(n819), .ZN(n814) );
  NOR2_X1 U912 ( .A1(n815), .A2(n814), .ZN(n816) );
  AND2_X1 U913 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U914 ( .A(n818), .B(KEYINPUT109), .ZN(n833) );
  NOR2_X1 U915 ( .A1(G1996), .A2(n895), .ZN(n938) );
  INV_X1 U916 ( .A(n819), .ZN(n822) );
  NOR2_X1 U917 ( .A1(G1986), .A2(G290), .ZN(n820) );
  NOR2_X1 U918 ( .A1(G1991), .A2(n885), .ZN(n930) );
  NOR2_X1 U919 ( .A1(n820), .A2(n930), .ZN(n821) );
  NOR2_X1 U920 ( .A1(n822), .A2(n821), .ZN(n823) );
  NOR2_X1 U921 ( .A1(n938), .A2(n823), .ZN(n824) );
  XNOR2_X1 U922 ( .A(n824), .B(KEYINPUT39), .ZN(n825) );
  XNOR2_X1 U923 ( .A(n825), .B(KEYINPUT110), .ZN(n826) );
  NAND2_X1 U924 ( .A1(n827), .A2(n826), .ZN(n829) );
  NAND2_X1 U925 ( .A1(n884), .A2(n828), .ZN(n926) );
  NAND2_X1 U926 ( .A1(n829), .A2(n926), .ZN(n831) );
  NAND2_X1 U927 ( .A1(n831), .A2(n830), .ZN(n832) );
  NAND2_X1 U928 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U929 ( .A(n834), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U930 ( .A(G223), .ZN(n835) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n835), .ZN(G217) );
  AND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n836) );
  NAND2_X1 U933 ( .A1(G661), .A2(n836), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U935 ( .A1(n838), .A2(n837), .ZN(n839) );
  XOR2_X1 U936 ( .A(KEYINPUT113), .B(n839), .Z(G188) );
  XOR2_X1 U937 ( .A(G96), .B(KEYINPUT114), .Z(G221) );
  INV_X1 U939 ( .A(G120), .ZN(G236) );
  INV_X1 U940 ( .A(G69), .ZN(G235) );
  INV_X1 U941 ( .A(n840), .ZN(n841) );
  NAND2_X1 U942 ( .A1(n842), .A2(n841), .ZN(G261) );
  INV_X1 U943 ( .A(G261), .ZN(G325) );
  XOR2_X1 U944 ( .A(G2454), .B(G2435), .Z(n844) );
  XNOR2_X1 U945 ( .A(G2438), .B(G2427), .ZN(n843) );
  XNOR2_X1 U946 ( .A(n844), .B(n843), .ZN(n851) );
  XOR2_X1 U947 ( .A(KEYINPUT111), .B(G2446), .Z(n846) );
  XNOR2_X1 U948 ( .A(G2443), .B(G2430), .ZN(n845) );
  XNOR2_X1 U949 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U950 ( .A(n847), .B(G2451), .Z(n849) );
  XNOR2_X1 U951 ( .A(G1348), .B(G1341), .ZN(n848) );
  XNOR2_X1 U952 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(n852) );
  NAND2_X1 U954 ( .A1(n852), .A2(G14), .ZN(n853) );
  XOR2_X1 U955 ( .A(KEYINPUT112), .B(n853), .Z(G401) );
  XNOR2_X1 U956 ( .A(G286), .B(n994), .ZN(n855) );
  XNOR2_X1 U957 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n856), .B(G301), .ZN(n857) );
  NOR2_X1 U959 ( .A1(G37), .A2(n857), .ZN(G397) );
  XOR2_X1 U960 ( .A(KEYINPUT115), .B(G1956), .Z(n859) );
  XNOR2_X1 U961 ( .A(G1986), .B(G1961), .ZN(n858) );
  XNOR2_X1 U962 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U963 ( .A(n860), .B(KEYINPUT41), .Z(n862) );
  XNOR2_X1 U964 ( .A(G1996), .B(G1991), .ZN(n861) );
  XNOR2_X1 U965 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U966 ( .A(G1976), .B(G1981), .Z(n864) );
  XNOR2_X1 U967 ( .A(G1966), .B(G1971), .ZN(n863) );
  XNOR2_X1 U968 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U969 ( .A(n866), .B(n865), .Z(n868) );
  XNOR2_X1 U970 ( .A(G2474), .B(KEYINPUT116), .ZN(n867) );
  XNOR2_X1 U971 ( .A(n868), .B(n867), .ZN(G229) );
  XOR2_X1 U972 ( .A(G2100), .B(G2096), .Z(n870) );
  XNOR2_X1 U973 ( .A(KEYINPUT42), .B(G2678), .ZN(n869) );
  XNOR2_X1 U974 ( .A(n870), .B(n869), .ZN(n874) );
  XOR2_X1 U975 ( .A(KEYINPUT43), .B(G2090), .Z(n872) );
  XNOR2_X1 U976 ( .A(G2067), .B(G2072), .ZN(n871) );
  XNOR2_X1 U977 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U978 ( .A(n874), .B(n873), .Z(n876) );
  XNOR2_X1 U979 ( .A(G2078), .B(G2084), .ZN(n875) );
  XNOR2_X1 U980 ( .A(n876), .B(n875), .ZN(G227) );
  NAND2_X1 U981 ( .A1(G124), .A2(n904), .ZN(n877) );
  XNOR2_X1 U982 ( .A(n877), .B(KEYINPUT44), .ZN(n879) );
  NAND2_X1 U983 ( .A1(n903), .A2(G112), .ZN(n878) );
  NAND2_X1 U984 ( .A1(n879), .A2(n878), .ZN(n883) );
  NAND2_X1 U985 ( .A1(G100), .A2(n907), .ZN(n881) );
  NAND2_X1 U986 ( .A1(G136), .A2(n908), .ZN(n880) );
  NAND2_X1 U987 ( .A1(n881), .A2(n880), .ZN(n882) );
  NOR2_X1 U988 ( .A1(n883), .A2(n882), .ZN(G162) );
  XNOR2_X1 U989 ( .A(G164), .B(n884), .ZN(n886) );
  XNOR2_X1 U990 ( .A(n886), .B(n885), .ZN(n897) );
  NAND2_X1 U991 ( .A1(G103), .A2(n907), .ZN(n888) );
  NAND2_X1 U992 ( .A1(G139), .A2(n908), .ZN(n887) );
  NAND2_X1 U993 ( .A1(n888), .A2(n887), .ZN(n893) );
  NAND2_X1 U994 ( .A1(G115), .A2(n903), .ZN(n890) );
  NAND2_X1 U995 ( .A1(G127), .A2(n904), .ZN(n889) );
  NAND2_X1 U996 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U997 ( .A(KEYINPUT47), .B(n891), .Z(n892) );
  NOR2_X1 U998 ( .A1(n893), .A2(n892), .ZN(n941) );
  XOR2_X1 U999 ( .A(G162), .B(n941), .Z(n894) );
  XNOR2_X1 U1000 ( .A(n895), .B(n894), .ZN(n896) );
  XOR2_X1 U1001 ( .A(n897), .B(n896), .Z(n902) );
  XOR2_X1 U1002 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n899) );
  XNOR2_X1 U1003 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n898) );
  XNOR2_X1 U1004 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U1005 ( .A(KEYINPUT117), .B(n900), .ZN(n901) );
  XNOR2_X1 U1006 ( .A(n902), .B(n901), .ZN(n917) );
  NAND2_X1 U1007 ( .A1(G118), .A2(n903), .ZN(n906) );
  NAND2_X1 U1008 ( .A1(G130), .A2(n904), .ZN(n905) );
  NAND2_X1 U1009 ( .A1(n906), .A2(n905), .ZN(n913) );
  NAND2_X1 U1010 ( .A1(G106), .A2(n907), .ZN(n910) );
  NAND2_X1 U1011 ( .A1(G142), .A2(n908), .ZN(n909) );
  NAND2_X1 U1012 ( .A1(n910), .A2(n909), .ZN(n911) );
  XOR2_X1 U1013 ( .A(KEYINPUT45), .B(n911), .Z(n912) );
  NOR2_X1 U1014 ( .A1(n913), .A2(n912), .ZN(n915) );
  XOR2_X1 U1015 ( .A(G160), .B(n934), .Z(n914) );
  XNOR2_X1 U1016 ( .A(n915), .B(n914), .ZN(n916) );
  XNOR2_X1 U1017 ( .A(n917), .B(n916), .ZN(n918) );
  NOR2_X1 U1018 ( .A1(G37), .A2(n918), .ZN(G395) );
  NOR2_X1 U1019 ( .A1(n919), .A2(G401), .ZN(n923) );
  NOR2_X1 U1020 ( .A1(G229), .A2(G227), .ZN(n920) );
  XNOR2_X1 U1021 ( .A(KEYINPUT49), .B(n920), .ZN(n921) );
  NOR2_X1 U1022 ( .A1(G397), .A2(n921), .ZN(n922) );
  NAND2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1024 ( .A1(n924), .A2(G395), .ZN(n925) );
  XNOR2_X1 U1025 ( .A(n925), .B(KEYINPUT120), .ZN(G308) );
  INV_X1 U1026 ( .A(G308), .ZN(G225) );
  INV_X1 U1027 ( .A(n926), .ZN(n928) );
  NOR2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n936) );
  XNOR2_X1 U1029 ( .A(G160), .B(G2084), .ZN(n932) );
  NOR2_X1 U1030 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n948) );
  XOR2_X1 U1034 ( .A(G2090), .B(G162), .Z(n937) );
  NOR2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1036 ( .A(KEYINPUT51), .B(n939), .Z(n940) );
  XOR2_X1 U1037 ( .A(KEYINPUT121), .B(n940), .Z(n946) );
  XOR2_X1 U1038 ( .A(G2072), .B(n941), .Z(n943) );
  XOR2_X1 U1039 ( .A(G164), .B(G2078), .Z(n942) );
  NOR2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1041 ( .A(KEYINPUT50), .B(n944), .ZN(n945) );
  NAND2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1044 ( .A(KEYINPUT52), .B(n949), .ZN(n950) );
  XOR2_X1 U1045 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n973) );
  NAND2_X1 U1046 ( .A1(n950), .A2(n973), .ZN(n951) );
  NAND2_X1 U1047 ( .A1(n951), .A2(G29), .ZN(n1031) );
  XNOR2_X1 U1048 ( .A(KEYINPUT54), .B(G34), .ZN(n952) );
  XNOR2_X1 U1049 ( .A(n952), .B(KEYINPUT125), .ZN(n953) );
  XNOR2_X1 U1050 ( .A(G2084), .B(n953), .ZN(n971) );
  XOR2_X1 U1051 ( .A(KEYINPUT53), .B(KEYINPUT123), .Z(n954) );
  XNOR2_X1 U1052 ( .A(KEYINPUT124), .B(n954), .ZN(n967) );
  XNOR2_X1 U1053 ( .A(G1991), .B(G25), .ZN(n956) );
  XNOR2_X1 U1054 ( .A(G33), .B(G2072), .ZN(n955) );
  NOR2_X1 U1055 ( .A1(n956), .A2(n955), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(n957), .B(G32), .ZN(n960) );
  XNOR2_X1 U1057 ( .A(G27), .B(n958), .ZN(n959) );
  NOR2_X1 U1058 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1059 ( .A1(n962), .A2(n961), .ZN(n965) );
  XOR2_X1 U1060 ( .A(G2067), .B(G26), .Z(n963) );
  NAND2_X1 U1061 ( .A1(G28), .A2(n963), .ZN(n964) );
  NOR2_X1 U1062 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1063 ( .A(n967), .B(n966), .ZN(n969) );
  XNOR2_X1 U1064 ( .A(G35), .B(G2090), .ZN(n968) );
  NOR2_X1 U1065 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(n973), .B(n972), .ZN(n975) );
  INV_X1 U1068 ( .A(G29), .ZN(n974) );
  NAND2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1070 ( .A1(G11), .A2(n976), .ZN(n1029) );
  XNOR2_X1 U1071 ( .A(G16), .B(KEYINPUT56), .ZN(n1000) );
  XNOR2_X1 U1072 ( .A(G301), .B(G1961), .ZN(n978) );
  XNOR2_X1 U1073 ( .A(G299), .B(G1956), .ZN(n977) );
  NOR2_X1 U1074 ( .A1(n978), .A2(n977), .ZN(n983) );
  XNOR2_X1 U1075 ( .A(n979), .B(G1341), .ZN(n981) );
  NOR2_X1 U1076 ( .A1(n1001), .A2(G166), .ZN(n980) );
  NOR2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n989) );
  XNOR2_X1 U1079 ( .A(G168), .B(G1966), .ZN(n985) );
  NAND2_X1 U1080 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1081 ( .A(n986), .B(KEYINPUT57), .ZN(n987) );
  XOR2_X1 U1082 ( .A(KEYINPUT126), .B(n987), .Z(n988) );
  NOR2_X1 U1083 ( .A1(n989), .A2(n988), .ZN(n998) );
  NOR2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n993) );
  NAND2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(G1348), .B(n994), .ZN(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1027) );
  INV_X1 U1090 ( .A(G16), .ZN(n1025) );
  XOR2_X1 U1091 ( .A(G1986), .B(G24), .Z(n1003) );
  XNOR2_X1 U1092 ( .A(n1001), .B(G22), .ZN(n1002) );
  NAND2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(G23), .B(G1976), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1096 ( .A(KEYINPUT58), .B(n1006), .ZN(n1011) );
  XNOR2_X1 U1097 ( .A(n1007), .B(G5), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(G21), .B(G1966), .ZN(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1022) );
  XNOR2_X1 U1101 ( .A(KEYINPUT59), .B(G4), .ZN(n1012) );
  XNOR2_X1 U1102 ( .A(n1012), .B(KEYINPUT127), .ZN(n1013) );
  XNOR2_X1 U1103 ( .A(G1348), .B(n1013), .ZN(n1015) );
  XNOR2_X1 U1104 ( .A(G1956), .B(G20), .ZN(n1014) );
  NOR2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(G1341), .B(G19), .ZN(n1017) );
  XNOR2_X1 U1107 ( .A(G1981), .B(G6), .ZN(n1016) );
  NOR2_X1 U1108 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1109 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1110 ( .A(KEYINPUT60), .B(n1020), .ZN(n1021) );
  NOR2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1112 ( .A(KEYINPUT61), .B(n1023), .ZN(n1024) );
  NAND2_X1 U1113 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1114 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NOR2_X1 U1115 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1116 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XOR2_X1 U1117 ( .A(KEYINPUT62), .B(n1032), .Z(G311) );
  INV_X1 U1118 ( .A(G311), .ZN(G150) );
endmodule

