//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 1 1 0 0 0 0 1 1 1 1 1 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n993, new_n994;
  XOR2_X1   g000(.A(G134gat), .B(G162gat), .Z(new_n202));
  AOI21_X1  g001(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT101), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT89), .ZN(new_n206));
  INV_X1    g005(.A(G29gat), .ZN(new_n207));
  INV_X1    g006(.A(G36gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT89), .B1(G29gat), .B2(G36gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(KEYINPUT14), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT14), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n212), .B(KEYINPUT89), .C1(G29gat), .C2(G36gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(G29gat), .A2(G36gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n211), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT15), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G50gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(G43gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n216), .B1(new_n219), .B2(KEYINPUT90), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n211), .A2(new_n220), .A3(new_n213), .A4(new_n214), .ZN(new_n221));
  XNOR2_X1  g020(.A(G43gat), .B(G50gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n217), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n211), .A2(new_n214), .ZN(new_n224));
  INV_X1    g023(.A(new_n222), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n224), .A2(new_n220), .A3(new_n213), .A4(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT91), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT91), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n223), .A2(new_n229), .A3(new_n226), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT99), .ZN(new_n231));
  NAND2_X1  g030(.A1(G99gat), .A2(G106gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT98), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(KEYINPUT98), .A2(G99gat), .A3(G106gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(KEYINPUT8), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT97), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT7), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(KEYINPUT97), .A2(KEYINPUT7), .ZN(new_n240));
  AND2_X1   g039(.A1(G85gat), .A2(G92gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(G85gat), .ZN(new_n243));
  INV_X1    g042(.A(G92gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n237), .B(new_n238), .C1(new_n243), .C2(new_n244), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n236), .A2(new_n242), .A3(new_n245), .A4(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(G99gat), .B(G106gat), .Z(new_n248));
  AOI21_X1  g047(.A(new_n231), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  AND2_X1   g048(.A1(new_n242), .A2(new_n246), .ZN(new_n250));
  INV_X1    g049(.A(new_n248), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n250), .A2(new_n251), .A3(new_n245), .A4(new_n236), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  OR3_X1    g052(.A1(new_n247), .A2(KEYINPUT99), .A3(new_n248), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n228), .A2(new_n230), .A3(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT100), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n256), .A2(KEYINPUT100), .A3(new_n257), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT17), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n228), .A2(new_n263), .A3(new_n230), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT92), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n255), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n223), .A2(KEYINPUT17), .A3(new_n226), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n228), .A2(KEYINPUT92), .A3(new_n263), .A4(new_n230), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n266), .A2(new_n267), .A3(new_n268), .A4(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(G190gat), .B(G218gat), .Z(new_n271));
  NAND3_X1  g070(.A1(new_n262), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n271), .ZN(new_n273));
  INV_X1    g072(.A(new_n270), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n256), .A2(KEYINPUT100), .A3(new_n257), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT100), .B1(new_n256), .B2(new_n257), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n273), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n205), .B(new_n272), .C1(new_n278), .C2(new_n204), .ZN(new_n279));
  XOR2_X1   g078(.A(G57gat), .B(G64gat), .Z(new_n280));
  NAND2_X1  g079(.A1(G71gat), .A2(G78gat), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT9), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OR2_X1    g082(.A1(G71gat), .A2(G78gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(new_n281), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n280), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G57gat), .B(G64gat), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n281), .B(new_n284), .C1(new_n287), .C2(new_n282), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT95), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n286), .A2(new_n288), .A3(KEYINPUT95), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(KEYINPUT21), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(G183gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(G15gat), .B(G22gat), .ZN(new_n294));
  OR2_X1    g093(.A1(new_n294), .A2(G1gat), .ZN(new_n295));
  INV_X1    g094(.A(G8gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT16), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n294), .B1(new_n297), .B2(G1gat), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n295), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n296), .B1(new_n295), .B2(new_n298), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n292), .A2(new_n293), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n293), .B1(new_n292), .B2(new_n301), .ZN(new_n304));
  OAI21_X1  g103(.A(G127gat), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n286), .A2(new_n288), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  XOR2_X1   g106(.A(KEYINPUT96), .B(G211gat), .Z(new_n308));
  NOR3_X1   g107(.A1(new_n307), .A2(KEYINPUT21), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G231gat), .A2(G233gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n308), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT21), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n311), .B1(new_n306), .B2(new_n312), .ZN(new_n313));
  OR3_X1    g112(.A1(new_n309), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n310), .B1(new_n309), .B2(new_n313), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n301), .ZN(new_n317));
  AND3_X1   g116(.A1(new_n286), .A2(new_n288), .A3(KEYINPUT95), .ZN(new_n318));
  NOR3_X1   g117(.A1(new_n318), .A2(new_n289), .A3(new_n312), .ZN(new_n319));
  OAI21_X1  g118(.A(G183gat), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G127gat), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(new_n321), .A3(new_n302), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n316), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n316), .B1(new_n305), .B2(new_n322), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n326), .B(G155gat), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NOR3_X1   g127(.A1(new_n324), .A2(new_n325), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n305), .A2(new_n322), .ZN(new_n330));
  INV_X1    g129(.A(new_n316), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n327), .B1(new_n332), .B2(new_n323), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n205), .ZN(new_n335));
  AND3_X1   g134(.A1(new_n262), .A2(new_n270), .A3(new_n271), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n271), .B1(new_n262), .B2(new_n270), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AND3_X1   g137(.A1(new_n279), .A2(new_n334), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  AND2_X1   g139(.A1(G228gat), .A2(G233gat), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT79), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT2), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT2), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT79), .ZN(new_n345));
  NAND2_X1  g144(.A1(G155gat), .A2(G162gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n343), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(G141gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G148gat), .ZN(new_n349));
  INV_X1    g148(.A(G148gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(G141gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(G155gat), .ZN(new_n354));
  INV_X1    g153(.A(G162gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n346), .A2(KEYINPUT78), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT78), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n358), .A2(G155gat), .A3(G162gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n353), .A2(new_n356), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT80), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n347), .A2(new_n352), .B1(new_n357), .B2(new_n359), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n364), .A2(KEYINPUT80), .A3(new_n356), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n366), .A2(new_n348), .A3(G148gat), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT81), .B1(new_n350), .B2(G141gat), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n350), .A2(G141gat), .ZN(new_n369));
  OAI211_X1 g168(.A(KEYINPUT82), .B(new_n367), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n366), .B1(new_n348), .B2(G148gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(new_n349), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT82), .B1(new_n373), .B2(new_n367), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n346), .B1(new_n356), .B2(KEYINPUT2), .ZN(new_n376));
  AOI22_X1  g175(.A1(new_n363), .A2(new_n365), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G197gat), .B(G204gat), .ZN(new_n378));
  XOR2_X1   g177(.A(KEYINPUT73), .B(KEYINPUT22), .Z(new_n379));
  INV_X1    g178(.A(G211gat), .ZN(new_n380));
  INV_X1    g179(.A(G218gat), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n378), .B1(new_n379), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT74), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  XOR2_X1   g184(.A(G211gat), .B(G218gat), .Z(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n385), .B(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT29), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT3), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n377), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n373), .A2(new_n367), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT82), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n395), .A2(new_n376), .A3(new_n370), .ZN(new_n396));
  XOR2_X1   g195(.A(KEYINPUT83), .B(KEYINPUT3), .Z(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  AND4_X1   g197(.A1(KEYINPUT80), .A2(new_n353), .A3(new_n356), .A4(new_n360), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT80), .B1(new_n364), .B2(new_n356), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n396), .B(new_n398), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n388), .B1(new_n389), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n341), .B1(new_n392), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n383), .A2(KEYINPUT86), .A3(new_n387), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n387), .B(KEYINPUT86), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n389), .B(new_n404), .C1(new_n405), .C2(new_n383), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n377), .B1(new_n406), .B2(new_n398), .ZN(new_n407));
  OR2_X1    g206(.A1(new_n407), .A2(new_n341), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n403), .B1(new_n402), .B2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G78gat), .B(G106gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(G22gat), .ZN(new_n411));
  XOR2_X1   g210(.A(KEYINPUT31), .B(G50gat), .Z(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n409), .B(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n388), .ZN(new_n416));
  NAND2_X1  g215(.A1(G226gat), .A2(G233gat), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT66), .ZN(new_n419));
  NAND2_X1  g218(.A1(G183gat), .A2(G190gat), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n420), .A2(KEYINPUT24), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT24), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n422), .B1(G183gat), .B2(G190gat), .ZN(new_n423));
  NOR2_X1   g222(.A1(G183gat), .A2(G190gat), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n421), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(G169gat), .A2(G176gat), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT65), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n427), .B(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT25), .ZN(new_n430));
  INV_X1    g229(.A(G169gat), .ZN(new_n431));
  INV_X1    g230(.A(G176gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT23), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n430), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n426), .A2(new_n429), .A3(new_n435), .ZN(new_n436));
  NOR3_X1   g235(.A1(new_n434), .A2(G169gat), .A3(G176gat), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n419), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n432), .A2(KEYINPUT64), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n432), .A2(KEYINPUT64), .ZN(new_n440));
  OAI211_X1 g239(.A(KEYINPUT23), .B(new_n431), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n434), .B1(G169gat), .B2(G176gat), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n426), .A2(new_n441), .A3(new_n427), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n430), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n427), .A2(new_n428), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n446));
  OAI211_X1 g245(.A(KEYINPUT25), .B(new_n442), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n422), .A2(G183gat), .A3(G190gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n420), .A2(KEYINPUT24), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n448), .B1(new_n449), .B2(new_n424), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n437), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(KEYINPUT66), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n438), .A2(new_n444), .A3(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(KEYINPUT27), .B(G183gat), .ZN(new_n455));
  INV_X1    g254(.A(G190gat), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OR2_X1    g256(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n458));
  OR2_X1    g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n457), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  OR2_X1    g260(.A1(new_n433), .A2(KEYINPUT26), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n433), .A2(KEYINPUT26), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(new_n427), .A3(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n459), .A2(new_n420), .A3(new_n461), .A4(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n454), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n418), .B1(new_n466), .B2(new_n389), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n417), .B1(new_n454), .B2(new_n465), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n416), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n466), .A2(new_n418), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT29), .B1(new_n454), .B2(new_n465), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n470), .B(new_n388), .C1(new_n418), .C2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT75), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT76), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n467), .A2(new_n468), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n388), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT75), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n474), .A2(new_n475), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n478), .B1(new_n469), .B2(new_n472), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT75), .B1(new_n476), .B2(new_n388), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT76), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G8gat), .B(G36gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(G64gat), .B(G92gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n485), .B(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n487), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n474), .A2(new_n479), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT30), .ZN(new_n491));
  OR2_X1    g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(new_n491), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n488), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  AND2_X1   g293(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n495));
  NOR2_X1   g294(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n496));
  OAI21_X1  g295(.A(G120gat), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT70), .ZN(new_n498));
  XNOR2_X1  g297(.A(KEYINPUT69), .B(G113gat), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT70), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(new_n500), .A3(G120gat), .ZN(new_n501));
  INV_X1    g300(.A(G113gat), .ZN(new_n502));
  XOR2_X1   g301(.A(KEYINPUT68), .B(G120gat), .Z(new_n503));
  OAI211_X1 g302(.A(new_n498), .B(new_n501), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  XOR2_X1   g303(.A(G127gat), .B(G134gat), .Z(new_n505));
  NOR2_X1   g304(.A1(new_n505), .A2(KEYINPUT1), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT1), .B1(G113gat), .B2(G120gat), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n508), .B1(G113gat), .B2(G120gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n401), .B(new_n511), .C1(new_n377), .C2(new_n391), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT4), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n396), .B1(new_n399), .B2(new_n400), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n513), .B1(new_n514), .B2(new_n511), .ZN(new_n515));
  AOI22_X1  g314(.A1(new_n504), .A2(new_n506), .B1(new_n505), .B2(new_n509), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n377), .A2(KEYINPUT4), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n512), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(G225gat), .A2(G233gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(KEYINPUT84), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  OR2_X1    g320(.A1(new_n521), .A2(KEYINPUT39), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n377), .A2(new_n516), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n514), .A2(new_n511), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n523), .A2(new_n524), .A3(KEYINPUT85), .ZN(new_n525));
  OR3_X1    g324(.A1(new_n377), .A2(KEYINPUT85), .A3(new_n516), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n521), .B(KEYINPUT39), .C1(new_n527), .C2(new_n520), .ZN(new_n528));
  XNOR2_X1  g327(.A(G1gat), .B(G29gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(G85gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(KEYINPUT0), .B(G57gat), .ZN(new_n531));
  XOR2_X1   g330(.A(new_n530), .B(new_n531), .Z(new_n532));
  NAND3_X1  g331(.A1(new_n522), .A2(new_n528), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT40), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT40), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n522), .A2(new_n528), .A3(new_n535), .A4(new_n532), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n515), .A2(new_n517), .ZN(new_n537));
  INV_X1    g336(.A(new_n520), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n537), .A2(KEYINPUT5), .A3(new_n538), .A4(new_n512), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n512), .A2(new_n538), .A3(new_n515), .A4(new_n517), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT5), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n532), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n525), .A2(new_n526), .A3(new_n520), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n539), .A2(new_n542), .A3(new_n543), .A4(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT87), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n545), .A2(new_n546), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n534), .A2(new_n536), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n494), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n539), .A2(new_n542), .A3(new_n544), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT6), .B1(new_n552), .B2(new_n532), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n545), .A2(new_n546), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n553), .B1(new_n554), .B2(new_n547), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT88), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n545), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT6), .ZN(new_n559));
  OAI211_X1 g358(.A(KEYINPUT88), .B(new_n553), .C1(new_n554), .C2(new_n547), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT37), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n474), .A2(new_n561), .A3(new_n479), .ZN(new_n562));
  AOI21_X1  g361(.A(KEYINPUT38), .B1(new_n473), .B2(KEYINPUT37), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(new_n487), .A3(new_n563), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n557), .A2(new_n559), .A3(new_n560), .A4(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n561), .B1(new_n480), .B2(new_n483), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n562), .A2(new_n487), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT38), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(new_n490), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n415), .B(new_n551), .C1(new_n565), .C2(new_n569), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n490), .A2(new_n491), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n553), .A2(new_n545), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n571), .B1(new_n559), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT77), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n488), .A2(new_n492), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n489), .B1(new_n480), .B2(new_n483), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n490), .A2(new_n491), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT77), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n573), .A2(new_n575), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(new_n414), .ZN(new_n580));
  XNOR2_X1  g379(.A(G71gat), .B(G99gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT71), .ZN(new_n582));
  XNOR2_X1  g381(.A(G15gat), .B(G43gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n466), .A2(new_n516), .ZN(new_n586));
  NAND2_X1  g385(.A1(G227gat), .A2(G233gat), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n454), .A2(new_n511), .A3(new_n465), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT33), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n585), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT34), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n594), .B1(new_n590), .B2(KEYINPUT32), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n590), .A2(KEYINPUT32), .A3(new_n594), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n586), .A2(new_n589), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(new_n587), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT72), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n596), .A2(new_n597), .A3(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n600), .B1(new_n596), .B2(new_n597), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n593), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n603), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n605), .A2(new_n592), .A3(new_n601), .ZN(new_n606));
  AND3_X1   g405(.A1(new_n604), .A2(KEYINPUT36), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT36), .B1(new_n604), .B2(new_n606), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n570), .A2(new_n580), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n414), .B1(new_n604), .B2(new_n606), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(KEYINPUT35), .B1(new_n579), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n557), .A2(new_n559), .A3(new_n560), .ZN(new_n614));
  INV_X1    g413(.A(new_n494), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT35), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n614), .A2(new_n615), .A3(new_n616), .A4(new_n611), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n340), .B1(new_n610), .B2(new_n618), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n266), .A2(new_n301), .A3(new_n268), .A4(new_n269), .ZN(new_n620));
  NAND2_X1  g419(.A1(G229gat), .A2(G233gat), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n228), .A2(new_n317), .A3(new_n230), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT94), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT18), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G113gat), .B(G141gat), .ZN(new_n627));
  INV_X1    g426(.A(G197gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(KEYINPUT11), .B(G169gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  AND2_X1   g431(.A1(new_n626), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n624), .B1(new_n623), .B2(new_n625), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n620), .A2(KEYINPUT18), .A3(new_n621), .A4(new_n622), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n228), .A2(new_n230), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n301), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n637), .A2(KEYINPUT93), .A3(new_n622), .ZN(new_n638));
  OR3_X1    g437(.A1(new_n636), .A2(KEYINPUT93), .A3(new_n301), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n621), .B(KEYINPUT13), .Z(new_n640));
  NAND3_X1  g439(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n635), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n634), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n623), .A2(new_n625), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n644), .A2(new_n641), .A3(new_n635), .ZN(new_n645));
  INV_X1    g444(.A(new_n632), .ZN(new_n646));
  AOI22_X1  g445(.A1(new_n633), .A2(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  XOR2_X1   g446(.A(G120gat), .B(G148gat), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(G204gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(KEYINPUT103), .B(G176gat), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n649), .B(new_n650), .Z(new_n651));
  NAND3_X1  g450(.A1(new_n253), .A2(new_n306), .A3(new_n254), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT10), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n247), .A2(new_n248), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n307), .A2(new_n252), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n652), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n318), .A2(new_n289), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n255), .A2(KEYINPUT10), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(G230gat), .A2(G233gat), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n652), .A2(new_n655), .ZN(new_n662));
  INV_X1    g461(.A(new_n660), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n651), .B1(new_n661), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT104), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT102), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n659), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n656), .A2(KEYINPUT102), .A3(new_n658), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n668), .A2(new_n660), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n670), .A2(new_n664), .A3(new_n651), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n666), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n647), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n619), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n572), .A2(new_n559), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(G1gat), .ZN(G1324gat));
  INV_X1    g477(.A(KEYINPUT42), .ZN(new_n679));
  NOR2_X1   g478(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n619), .A2(new_n494), .A3(new_n673), .A4(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n297), .A2(new_n296), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n679), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n685));
  OR2_X1    g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n682), .A2(new_n679), .A3(new_n683), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n296), .B1(new_n674), .B2(new_n494), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n684), .A2(new_n685), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n686), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT106), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n686), .A2(new_n689), .A3(KEYINPUT106), .A4(new_n690), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(G1325gat));
  NAND2_X1  g494(.A1(new_n604), .A2(new_n606), .ZN(new_n696));
  AOI21_X1  g495(.A(G15gat), .B1(new_n674), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n609), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n698), .A2(G15gat), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n697), .B1(new_n674), .B2(new_n699), .ZN(G1326gat));
  NAND2_X1  g499(.A1(new_n674), .A2(new_n414), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(G22gat), .ZN(new_n702));
  XNOR2_X1  g501(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1327gat));
  NAND2_X1  g503(.A1(new_n610), .A2(new_n618), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n279), .A2(new_n338), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n706), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n710), .B1(new_n610), .B2(new_n618), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(KEYINPUT44), .ZN(new_n712));
  INV_X1    g511(.A(new_n334), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n673), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n709), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(G29gat), .B1(new_n717), .B2(new_n675), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n711), .A2(new_n715), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n719), .A2(G29gat), .A3(new_n675), .ZN(new_n720));
  XNOR2_X1  g519(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n718), .A2(new_n722), .ZN(G1328gat));
  OAI21_X1  g522(.A(G36gat), .B1(new_n717), .B2(new_n615), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n711), .A2(new_n208), .A3(new_n494), .A4(new_n715), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n725), .B1(new_n726), .B2(KEYINPUT46), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT46), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n727), .B1(KEYINPUT109), .B2(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n725), .A2(new_n726), .A3(KEYINPUT46), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n724), .A2(new_n729), .A3(new_n730), .ZN(G1329gat));
  NAND4_X1  g530(.A1(new_n709), .A2(new_n698), .A3(new_n712), .A4(new_n715), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(G43gat), .ZN(new_n733));
  INV_X1    g532(.A(G43gat), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n711), .A2(new_n734), .A3(new_n696), .A4(new_n715), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n733), .A2(KEYINPUT47), .A3(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT111), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n735), .B(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n733), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT47), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n737), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AOI211_X1 g541(.A(KEYINPUT111), .B(KEYINPUT47), .C1(new_n739), .C2(new_n733), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n736), .B1(new_n742), .B2(new_n743), .ZN(G1330gat));
  AOI21_X1  g543(.A(new_n218), .B1(new_n716), .B2(new_n414), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n711), .A2(new_n218), .A3(new_n414), .A4(new_n715), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT48), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  OR3_X1    g548(.A1(new_n745), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n745), .B2(new_n747), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(G1331gat));
  NAND4_X1  g551(.A1(new_n705), .A2(new_n339), .A3(new_n647), .A4(new_n672), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT113), .ZN(new_n754));
  OR2_X1    g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n676), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g559(.A1(new_n757), .A2(new_n615), .ZN(new_n761));
  NOR2_X1   g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  AND2_X1   g561(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n761), .B2(new_n762), .ZN(G1333gat));
  OAI21_X1  g564(.A(G71gat), .B1(new_n757), .B2(new_n609), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT50), .ZN(new_n767));
  INV_X1    g566(.A(G71gat), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n755), .A2(new_n768), .A3(new_n696), .A4(new_n756), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n766), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n767), .B1(new_n766), .B2(new_n769), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n770), .A2(new_n771), .ZN(G1334gat));
  NAND2_X1  g571(.A1(new_n758), .A2(new_n414), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(G78gat), .ZN(G1335gat));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n709), .A2(new_n712), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n647), .A2(new_n713), .ZN(new_n777));
  INV_X1    g576(.A(new_n672), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n775), .B1(new_n780), .B2(new_n675), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n776), .A2(KEYINPUT114), .A3(new_n676), .A4(new_n779), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n781), .A2(G85gat), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n777), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n705), .A2(new_n706), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT51), .B1(new_n711), .B2(new_n784), .ZN(new_n788));
  OR2_X1    g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n789), .A2(new_n672), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n790), .A2(new_n243), .A3(new_n676), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n783), .A2(new_n791), .ZN(G1336gat));
  NAND3_X1  g591(.A1(new_n776), .A2(new_n494), .A3(new_n779), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(G92gat), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n494), .A2(new_n244), .A3(new_n672), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(KEYINPUT115), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT52), .B1(new_n789), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT116), .ZN(new_n800));
  AOI211_X1 g599(.A(new_n800), .B(new_n786), .C1(new_n711), .C2(new_n784), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT51), .B1(new_n785), .B2(KEYINPUT116), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI22_X1  g602(.A1(new_n793), .A2(G92gat), .B1(new_n803), .B2(new_n796), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n798), .B1(new_n799), .B2(new_n804), .ZN(G1337gat));
  INV_X1    g604(.A(G99gat), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n780), .A2(new_n806), .A3(new_n609), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n790), .A2(new_n696), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n807), .B1(new_n808), .B2(new_n806), .ZN(G1338gat));
  NAND4_X1  g608(.A1(new_n709), .A2(new_n414), .A3(new_n712), .A4(new_n779), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(G106gat), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n415), .A2(G106gat), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n672), .B(new_n813), .C1(new_n787), .C2(new_n788), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n811), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  AOI211_X1 g614(.A(new_n710), .B(new_n777), .C1(new_n610), .C2(new_n618), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n786), .B1(new_n816), .B2(new_n800), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n785), .A2(KEYINPUT116), .A3(KEYINPUT51), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n778), .A2(new_n415), .A3(G106gat), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n812), .B1(new_n811), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT117), .B1(new_n815), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n811), .A2(new_n812), .A3(new_n814), .ZN(new_n824));
  AOI22_X1  g623(.A1(new_n803), .A2(new_n819), .B1(G106gat), .B2(new_n810), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n823), .B(new_n824), .C1(new_n825), .C2(new_n812), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n822), .A2(new_n826), .ZN(G1339gat));
  INV_X1    g626(.A(new_n634), .ZN(new_n828));
  INV_X1    g627(.A(new_n642), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n828), .A2(new_n829), .A3(new_n632), .A4(new_n626), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n621), .B1(new_n620), .B2(new_n622), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n640), .B1(new_n638), .B2(new_n639), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n631), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n830), .A2(new_n672), .A3(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT119), .ZN(new_n836));
  AND3_X1   g635(.A1(new_n656), .A2(KEYINPUT102), .A3(new_n658), .ZN(new_n837));
  AOI21_X1  g636(.A(KEYINPUT102), .B1(new_n656), .B2(new_n658), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n837), .A2(new_n838), .A3(new_n663), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n659), .A2(new_n660), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n836), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT54), .B1(new_n840), .B2(new_n836), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n659), .A2(new_n845), .A3(new_n660), .ZN(new_n846));
  INV_X1    g645(.A(new_n651), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n846), .A2(KEYINPUT120), .A3(new_n847), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n835), .B1(new_n844), .B2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n840), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n670), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n842), .B1(new_n856), .B2(new_n836), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n857), .A2(new_n852), .A3(KEYINPUT55), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n671), .B1(new_n854), .B2(new_n858), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n710), .B(new_n834), .C1(new_n859), .C2(new_n647), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n830), .A2(new_n833), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n706), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n860), .A2(new_n713), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n339), .A2(new_n647), .A3(new_n778), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(KEYINPUT118), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n339), .A2(new_n647), .A3(new_n866), .A4(new_n778), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT121), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT121), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n863), .A2(new_n868), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n612), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n494), .A2(new_n675), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n647), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(new_n499), .A3(new_n877), .ZN(new_n878));
  OR2_X1    g677(.A1(new_n875), .A2(KEYINPUT122), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n875), .A2(KEYINPUT122), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n647), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n878), .B1(new_n881), .B2(new_n502), .ZN(G1340gat));
  OR3_X1    g681(.A1(new_n875), .A2(new_n503), .A3(new_n778), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n778), .B1(new_n879), .B2(new_n880), .ZN(new_n884));
  INV_X1    g683(.A(G120gat), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(G1341gat));
  AOI21_X1  g685(.A(G127gat), .B1(new_n876), .B2(new_n334), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n713), .B1(new_n879), .B2(new_n880), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(new_n888), .B2(G127gat), .ZN(G1342gat));
  NOR3_X1   g688(.A1(new_n875), .A2(G134gat), .A3(new_n710), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT56), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n891), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n710), .B1(new_n879), .B2(new_n880), .ZN(new_n894));
  INV_X1    g693(.A(G134gat), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n892), .B(new_n893), .C1(new_n894), .C2(new_n895), .ZN(G1343gat));
  INV_X1    g695(.A(KEYINPUT57), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n863), .A2(new_n868), .A3(new_n871), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n871), .B1(new_n863), .B2(new_n868), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n897), .B(new_n414), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n698), .A2(new_n675), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n615), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n869), .A2(new_n414), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n903), .B2(KEYINPUT57), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n900), .A2(new_n904), .A3(new_n877), .ZN(new_n905));
  AOI21_X1  g704(.A(KEYINPUT58), .B1(new_n905), .B2(G141gat), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n414), .B(new_n901), .C1(new_n898), .C2(new_n899), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT123), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n870), .A2(new_n872), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n910), .A2(KEYINPUT123), .A3(new_n414), .A4(new_n901), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n647), .A2(G141gat), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n909), .A2(new_n911), .A3(new_n615), .A4(new_n912), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n906), .A2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT58), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n905), .A2(G141gat), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n415), .B1(new_n870), .B2(new_n872), .ZN(new_n917));
  INV_X1    g716(.A(new_n902), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n917), .A2(new_n918), .A3(new_n912), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n915), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(KEYINPUT124), .B1(new_n914), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n913), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT124), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n917), .A2(new_n918), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  AOI22_X1  g724(.A1(new_n925), .A2(new_n912), .B1(new_n905), .B2(G141gat), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n922), .B(new_n923), .C1(new_n915), .C2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n921), .A2(new_n927), .ZN(G1344gat));
  INV_X1    g727(.A(KEYINPUT59), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n917), .A2(new_n897), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n863), .A2(new_n864), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n931), .A2(new_n897), .A3(new_n414), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n930), .A2(new_n672), .A3(new_n918), .A4(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n929), .B1(new_n933), .B2(G148gat), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n900), .A2(new_n904), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n929), .B1(new_n935), .B2(new_n778), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n936), .A2(new_n350), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n909), .A2(new_n911), .A3(new_n615), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n672), .A2(new_n350), .ZN(new_n939));
  OAI22_X1  g738(.A1(new_n934), .A2(new_n937), .B1(new_n938), .B2(new_n939), .ZN(G1345gat));
  NAND2_X1  g739(.A1(new_n334), .A2(G155gat), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT125), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n935), .A2(new_n942), .ZN(new_n943));
  OR2_X1    g742(.A1(new_n938), .A2(new_n713), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n943), .B1(new_n944), .B2(new_n354), .ZN(G1346gat));
  OAI21_X1  g744(.A(G162gat), .B1(new_n935), .B2(new_n710), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n706), .A2(new_n355), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n946), .B1(new_n938), .B2(new_n947), .ZN(G1347gat));
  NOR2_X1   g747(.A1(new_n615), .A2(new_n676), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n873), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n950), .A2(new_n647), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(new_n431), .ZN(G1348gat));
  INV_X1    g751(.A(new_n950), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(new_n672), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(G176gat), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n439), .A2(new_n440), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n955), .B1(new_n954), .B2(new_n956), .ZN(G1349gat));
  NAND3_X1  g756(.A1(new_n953), .A2(new_n455), .A3(new_n334), .ZN(new_n958));
  OAI21_X1  g757(.A(G183gat), .B1(new_n950), .B2(new_n713), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT60), .ZN(G1350gat));
  NAND4_X1  g760(.A1(new_n953), .A2(KEYINPUT61), .A3(G190gat), .A4(new_n706), .ZN(new_n962));
  XOR2_X1   g761(.A(KEYINPUT61), .B(G190gat), .Z(new_n963));
  OAI21_X1  g762(.A(new_n963), .B1(new_n950), .B2(new_n710), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n962), .A2(new_n964), .ZN(G1351gat));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n609), .ZN(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n930), .A2(new_n932), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(G197gat), .B1(new_n968), .B2(new_n647), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n917), .A2(new_n967), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n971), .A2(new_n628), .A3(new_n877), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n969), .A2(new_n972), .ZN(G1352gat));
  NAND3_X1  g772(.A1(new_n930), .A2(new_n672), .A3(new_n932), .ZN(new_n974));
  OAI21_X1  g773(.A(G204gat), .B1(new_n974), .B2(new_n966), .ZN(new_n975));
  NOR3_X1   g774(.A1(new_n970), .A2(G204gat), .A3(new_n778), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT62), .ZN(new_n977));
  OR2_X1    g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n976), .A2(new_n977), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n975), .A2(new_n978), .A3(new_n979), .ZN(G1353gat));
  NAND4_X1  g779(.A1(new_n930), .A2(new_n334), .A3(new_n932), .A4(new_n967), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT127), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT63), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n981), .A2(G211gat), .A3(new_n984), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n982), .A2(new_n983), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND4_X1  g786(.A1(new_n917), .A2(new_n380), .A3(new_n334), .A4(new_n967), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n988), .B(KEYINPUT126), .ZN(new_n989));
  INV_X1    g788(.A(new_n986), .ZN(new_n990));
  NAND4_X1  g789(.A1(new_n981), .A2(G211gat), .A3(new_n984), .A4(new_n990), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n987), .A2(new_n989), .A3(new_n991), .ZN(G1354gat));
  OAI21_X1  g791(.A(G218gat), .B1(new_n968), .B2(new_n710), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n971), .A2(new_n381), .A3(new_n706), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n993), .A2(new_n994), .ZN(G1355gat));
endmodule


