//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 0 1 1 1 1 0 1 1 0 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n571, new_n572, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n594, new_n596, new_n597, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1122, new_n1123;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT67), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n454), .A2(G2106), .ZN(new_n460));
  NAND3_X1  g035(.A1(new_n457), .A2(KEYINPUT68), .A3(G567), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n462));
  INV_X1    g037(.A(G567), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n462), .B1(new_n456), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n460), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(G319));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n470), .A2(G137), .B1(G101), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n474), .B1(new_n469), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(G112), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(new_n481), .B2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n470), .A2(G136), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  XNOR2_X1  g059(.A(KEYINPUT3), .B(G2104), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  AOI211_X1 g062(.A(new_n482), .B(new_n484), .C1(G124), .C2(new_n487), .ZN(G162));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n489));
  NAND2_X1  g064(.A1(G126), .A2(G2105), .ZN(new_n490));
  OR2_X1    g065(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n491));
  NAND2_X1  g066(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G2105), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n489), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n490), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n499), .B1(new_n467), .B2(new_n468), .ZN(new_n500));
  INV_X1    g075(.A(G102), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(new_n494), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G2105), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n502), .A2(new_n504), .A3(G2104), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n500), .A2(new_n505), .A3(KEYINPUT69), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n507));
  INV_X1    g082(.A(G138), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n508), .A2(G2105), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n507), .B1(new_n485), .B2(new_n509), .ZN(new_n510));
  OAI211_X1 g085(.A(new_n509), .B(new_n507), .C1(new_n468), .C2(new_n467), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  OAI211_X1 g087(.A(new_n498), .B(new_n506), .C1(new_n510), .C2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(G164));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n516), .B2(KEYINPUT71), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT71), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n518), .A2(KEYINPUT5), .A3(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n520), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n521));
  INV_X1    g096(.A(G651), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT6), .B(G651), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(G543), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n525), .A2(G88), .B1(new_n527), .B2(G50), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(KEYINPUT72), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT72), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n523), .A2(new_n528), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n530), .A2(new_n532), .ZN(G166));
  AND2_X1   g108(.A1(new_n525), .A2(G89), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n520), .A2(G63), .A3(G651), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  INV_X1    g112(.A(G51), .ZN(new_n538));
  OAI211_X1 g113(.A(new_n535), .B(new_n537), .C1(new_n526), .C2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n534), .A2(new_n539), .ZN(G168));
  AOI22_X1  g115(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n541), .A2(new_n522), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n527), .A2(G52), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n520), .A2(G90), .A3(new_n524), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT73), .ZN(new_n545));
  AND3_X1   g120(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n545), .B1(new_n543), .B2(new_n544), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n542), .B1(new_n546), .B2(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  AOI22_X1  g124(.A1(new_n520), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(new_n522), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n525), .A2(G81), .B1(new_n527), .B2(G43), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  NAND2_X1  g134(.A1(new_n527), .A2(G53), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT74), .ZN(new_n563));
  INV_X1    g138(.A(new_n520), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n566), .A2(G651), .B1(new_n525), .B2(G91), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n561), .A2(new_n567), .ZN(G299));
  INV_X1    g143(.A(G168), .ZN(G286));
  INV_X1    g144(.A(G166), .ZN(G303));
  AOI22_X1  g145(.A1(new_n525), .A2(G87), .B1(new_n527), .B2(G49), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(G288));
  AOI22_X1  g148(.A1(new_n520), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n574));
  OR2_X1    g149(.A1(new_n574), .A2(new_n522), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n525), .A2(G86), .B1(new_n527), .B2(G48), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(G305));
  AOI22_X1  g152(.A1(new_n525), .A2(G85), .B1(new_n527), .B2(G47), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n522), .B2(new_n579), .ZN(G290));
  NAND2_X1  g155(.A1(G301), .A2(G868), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n525), .A2(G92), .ZN(new_n582));
  XOR2_X1   g157(.A(new_n582), .B(KEYINPUT10), .Z(new_n583));
  NAND2_X1  g158(.A1(G79), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G66), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n564), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n586), .A2(G651), .B1(G54), .B2(new_n527), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n581), .B1(new_n589), .B2(G868), .ZN(G284));
  OAI21_X1  g165(.A(new_n581), .B1(new_n589), .B2(G868), .ZN(G321));
  MUX2_X1   g166(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g167(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g168(.A(G559), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n589), .B1(new_n594), .B2(G860), .ZN(G148));
  NAND2_X1  g170(.A1(new_n589), .A2(new_n594), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(G868), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g173(.A(KEYINPUT75), .B(KEYINPUT11), .ZN(new_n599));
  XNOR2_X1  g174(.A(G323), .B(new_n599), .ZN(G282));
  NAND2_X1  g175(.A1(new_n485), .A2(new_n472), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT12), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT13), .ZN(new_n603));
  INV_X1    g178(.A(G2100), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n606));
  INV_X1    g181(.A(G111), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(G2105), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n487), .A2(G123), .ZN(new_n609));
  XOR2_X1   g184(.A(new_n609), .B(KEYINPUT76), .Z(new_n610));
  AOI211_X1 g185(.A(new_n608), .B(new_n610), .C1(G135), .C2(new_n470), .ZN(new_n611));
  INV_X1    g186(.A(G2096), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n605), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n603), .A2(new_n604), .ZN(new_n614));
  OAI211_X1 g189(.A(new_n613), .B(new_n614), .C1(new_n612), .C2(new_n611), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT77), .Z(G156));
  XOR2_X1   g191(.A(KEYINPUT15), .B(G2435), .Z(new_n617));
  XOR2_X1   g192(.A(KEYINPUT79), .B(G2438), .Z(new_n618));
  XOR2_X1   g193(.A(new_n617), .B(new_n618), .Z(new_n619));
  XNOR2_X1  g194(.A(G2427), .B(G2430), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(KEYINPUT14), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT80), .Z(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(new_n620), .B2(new_n619), .ZN(new_n624));
  XOR2_X1   g199(.A(G1341), .B(G1348), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2451), .B(G2454), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n626), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2443), .B(G2446), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n632), .A2(G14), .A3(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(G401));
  XOR2_X1   g210(.A(G2084), .B(G2090), .Z(new_n636));
  XNOR2_X1  g211(.A(G2067), .B(G2678), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G2072), .B(G2078), .Z(new_n639));
  NOR2_X1   g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT18), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n639), .B(KEYINPUT17), .ZN(new_n642));
  INV_X1    g217(.A(new_n636), .ZN(new_n643));
  INV_X1    g218(.A(new_n637), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n643), .A2(new_n639), .A3(new_n644), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(new_n638), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n641), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2096), .B(G2100), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(G227));
  XOR2_X1   g225(.A(G1971), .B(G1976), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT19), .ZN(new_n652));
  XOR2_X1   g227(.A(G1956), .B(G2474), .Z(new_n653));
  XOR2_X1   g228(.A(G1961), .B(G1966), .Z(new_n654));
  AND2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT20), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n653), .A2(new_n654), .ZN(new_n658));
  NOR3_X1   g233(.A1(new_n652), .A2(new_n655), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n659), .B1(new_n652), .B2(new_n658), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT81), .Z(new_n662));
  XNOR2_X1  g237(.A(G1981), .B(G1986), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT82), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n664), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1991), .B(G1996), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(G229));
  INV_X1    g245(.A(G29), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(G35), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(G162), .B2(new_n671), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT29), .Z(new_n674));
  INV_X1    g249(.A(G2090), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  INV_X1    g252(.A(G1348), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n589), .A2(G16), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(G4), .B2(G16), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n676), .B(new_n677), .C1(new_n678), .C2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(new_n678), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT91), .B(KEYINPUT24), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(G34), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n684), .A2(G29), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(G160), .B2(G29), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n686), .A2(G2084), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(G2084), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT30), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT93), .ZN(new_n690));
  AND3_X1   g265(.A1(new_n690), .A2(new_n689), .A3(G28), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n690), .B1(new_n689), .B2(G28), .ZN(new_n692));
  OAI221_X1 g267(.A(new_n671), .B1(new_n689), .B2(G28), .C1(new_n691), .C2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT31), .B(G11), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(new_n611), .B2(G29), .ZN(new_n696));
  NAND4_X1  g271(.A1(new_n682), .A2(new_n687), .A3(new_n688), .A4(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G21), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G168), .B2(new_n698), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n700), .A2(G1966), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n671), .A2(G26), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT28), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n487), .A2(G128), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n470), .A2(G140), .ZN(new_n705));
  OR2_X1    g280(.A1(G104), .A2(G2105), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n706), .B(G2104), .C1(G116), .C2(new_n494), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n704), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n703), .B1(new_n709), .B2(new_n671), .ZN(new_n710));
  INV_X1    g285(.A(G2067), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n700), .A2(G1966), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR4_X1   g289(.A1(new_n681), .A2(new_n697), .A3(new_n701), .A4(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n671), .A2(G32), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n470), .A2(G141), .B1(G105), .B2(new_n472), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n487), .A2(G129), .ZN(new_n718));
  NAND3_X1  g293(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT26), .Z(new_n720));
  NAND3_X1  g295(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT92), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n716), .B1(new_n723), .B2(new_n671), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT27), .ZN(new_n725));
  INV_X1    g300(.A(G1996), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(G5), .A2(G16), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT94), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G301), .B2(new_n698), .ZN(new_n730));
  INV_X1    g305(.A(G1961), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT95), .Z(new_n733));
  NOR2_X1   g308(.A1(new_n727), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(G16), .A2(G19), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(new_n554), .B2(G16), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT88), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G1341), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n671), .A2(G33), .ZN(new_n739));
  NAND2_X1  g314(.A1(G115), .A2(G2104), .ZN(new_n740));
  INV_X1    g315(.A(G127), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n740), .B1(new_n469), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n494), .B1(new_n742), .B2(KEYINPUT89), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(KEYINPUT89), .B2(new_n742), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n494), .A2(G103), .A3(G2104), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT25), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G139), .B2(new_n470), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT90), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n739), .B1(new_n749), .B2(new_n671), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n750), .A2(G2072), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n750), .A2(G2072), .ZN(new_n752));
  NOR3_X1   g327(.A1(new_n738), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n730), .A2(new_n731), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n671), .A2(G27), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G164), .B2(new_n671), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT96), .B(G2078), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n754), .B1(new_n758), .B2(KEYINPUT97), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n698), .A2(G20), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT23), .Z(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G299), .B2(G16), .ZN(new_n762));
  INV_X1    g337(.A(G1956), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  AOI211_X1 g339(.A(new_n759), .B(new_n764), .C1(KEYINPUT97), .C2(new_n758), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n715), .A2(new_n734), .A3(new_n753), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n698), .A2(G22), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G166), .B2(new_n698), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT85), .B(G1971), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n771), .A2(KEYINPUT86), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(KEYINPUT86), .ZN(new_n773));
  MUX2_X1   g348(.A(G6), .B(G305), .S(G16), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT32), .ZN(new_n775));
  INV_X1    g350(.A(G1981), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n698), .A2(G23), .ZN(new_n778));
  INV_X1    g353(.A(G288), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n778), .B1(new_n779), .B2(new_n698), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT33), .B(G1976), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n772), .A2(new_n773), .A3(new_n777), .A4(new_n782), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n783), .A2(KEYINPUT34), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(KEYINPUT34), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n671), .A2(G25), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT83), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n487), .A2(G119), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n470), .A2(G131), .ZN(new_n789));
  OR2_X1    g364(.A1(G95), .A2(G2105), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n790), .B(G2104), .C1(G107), .C2(new_n494), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n788), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n787), .B1(new_n793), .B2(new_n671), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT35), .B(G1991), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n698), .A2(G24), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT84), .Z(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G290), .B2(G16), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G1986), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n784), .A2(new_n785), .A3(new_n796), .A4(new_n800), .ZN(new_n801));
  AND2_X1   g376(.A1(KEYINPUT87), .A2(KEYINPUT36), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n766), .B1(new_n803), .B2(new_n804), .ZN(G311));
  INV_X1    g380(.A(G311), .ZN(G150));
  AND2_X1   g381(.A1(new_n525), .A2(G93), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n520), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n808), .A2(new_n522), .ZN(new_n809));
  AOI211_X1 g384(.A(new_n807), .B(new_n809), .C1(G55), .C2(new_n527), .ZN(new_n810));
  INV_X1    g385(.A(G860), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT37), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n594), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT99), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n814), .B(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n810), .B(new_n554), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n817), .B(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(KEYINPUT39), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT100), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n811), .B1(new_n821), .B2(KEYINPUT39), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n813), .B1(new_n823), .B2(new_n824), .ZN(G145));
  OAI21_X1  g400(.A(KEYINPUT101), .B1(new_n512), .B2(new_n510), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n509), .B1(new_n467), .B2(new_n468), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n827), .A2(KEYINPUT70), .A3(KEYINPUT4), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT101), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n828), .A2(new_n829), .A3(new_n511), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n500), .A2(new_n505), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n826), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n749), .B(new_n833), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n487), .A2(G130), .B1(new_n470), .B2(G142), .ZN(new_n835));
  NOR3_X1   g410(.A1(new_n494), .A2(KEYINPUT102), .A3(G118), .ZN(new_n836));
  OAI21_X1  g411(.A(KEYINPUT102), .B1(new_n494), .B2(G118), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n837), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n835), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT103), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(new_n602), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n834), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n722), .B(new_n708), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n792), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n842), .B(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(G162), .B(new_n478), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n611), .B(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(G37), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n847), .B2(new_n845), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g425(.A(G166), .B(G288), .ZN(new_n851));
  XOR2_X1   g426(.A(G290), .B(G305), .Z(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(KEYINPUT104), .B2(KEYINPUT42), .ZN(new_n854));
  NAND2_X1  g429(.A1(KEYINPUT104), .A2(KEYINPUT42), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n588), .B(G299), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT41), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n818), .B(new_n596), .Z(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n857), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n861), .B1(new_n862), .B2(new_n860), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n856), .B(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(G868), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n865), .B1(G868), .B2(new_n810), .ZN(G295));
  OAI21_X1  g441(.A(new_n865), .B1(G868), .B2(new_n810), .ZN(G331));
  AND2_X1   g442(.A1(G301), .A2(KEYINPUT105), .ZN(new_n868));
  OAI21_X1  g443(.A(G168), .B1(G301), .B2(KEYINPUT105), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n870), .A2(new_n818), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n818), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n872), .A2(new_n862), .A3(new_n873), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n870), .A2(new_n818), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(KEYINPUT106), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT106), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n871), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n853), .B(new_n874), .C1(new_n879), .C2(new_n859), .ZN(new_n880));
  AOI21_X1  g455(.A(G37), .B1(new_n880), .B2(KEYINPUT107), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n876), .A2(new_n878), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n858), .B1(new_n882), .B2(new_n871), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT107), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n883), .A2(new_n884), .A3(new_n853), .A4(new_n874), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n874), .B1(new_n879), .B2(new_n859), .ZN(new_n886));
  INV_X1    g461(.A(new_n853), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n881), .A2(new_n885), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT43), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n858), .B1(new_n871), .B2(new_n875), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT108), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n872), .A2(new_n862), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n894), .B1(new_n882), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n892), .A2(new_n893), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n887), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AND4_X1   g473(.A1(KEYINPUT43), .A2(new_n881), .A3(new_n898), .A4(new_n885), .ZN(new_n899));
  OAI21_X1  g474(.A(KEYINPUT44), .B1(new_n891), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n889), .A2(KEYINPUT43), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n881), .A2(new_n898), .A3(new_n885), .A4(new_n890), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n900), .A2(new_n905), .ZN(G397));
  INV_X1    g481(.A(G1384), .ZN(new_n907));
  AOI21_X1  g482(.A(KEYINPUT45), .B1(new_n833), .B2(new_n907), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n473), .A2(G40), .A3(new_n477), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(KEYINPUT109), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n708), .B(G2067), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n910), .A2(G1996), .ZN(new_n915));
  OAI221_X1 g490(.A(new_n914), .B1(KEYINPUT46), .B2(new_n915), .C1(new_n723), .C2(new_n911), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(KEYINPUT46), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT127), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(KEYINPUT47), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n914), .B(KEYINPUT110), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n915), .B1(new_n912), .B2(new_n722), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n922), .B1(new_n726), .B2(new_n722), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n924), .A2(new_n795), .A3(new_n793), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n709), .A2(new_n711), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n911), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n792), .B(new_n795), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT111), .ZN(new_n929));
  AOI211_X1 g504(.A(new_n921), .B(new_n923), .C1(new_n912), .C2(new_n929), .ZN(new_n930));
  NOR3_X1   g505(.A1(new_n910), .A2(G1986), .A3(G290), .ZN(new_n931));
  XOR2_X1   g506(.A(new_n931), .B(KEYINPUT48), .Z(new_n932));
  AOI211_X1 g507(.A(new_n920), .B(new_n927), .C1(new_n930), .C2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(KEYINPUT114), .B(G8), .ZN(new_n934));
  NOR2_X1   g509(.A1(G168), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n909), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n908), .A2(new_n936), .ZN(new_n937));
  AOI22_X1  g512(.A1(new_n828), .A2(new_n511), .B1(new_n831), .B2(new_n489), .ZN(new_n938));
  AOI21_X1  g513(.A(G1384), .B1(new_n938), .B2(new_n506), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(KEYINPUT45), .ZN(new_n940));
  AOI21_X1  g515(.A(G1966), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n513), .A2(new_n907), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT50), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT50), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n833), .A2(new_n944), .A3(new_n907), .ZN(new_n945));
  INV_X1    g520(.A(G2084), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n943), .A2(new_n945), .A3(new_n946), .A4(new_n909), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n935), .B1(new_n941), .B2(new_n948), .ZN(new_n949));
  XOR2_X1   g524(.A(KEYINPUT124), .B(KEYINPUT51), .Z(new_n950));
  INV_X1    g525(.A(G8), .ZN(new_n951));
  INV_X1    g526(.A(new_n908), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n952), .A2(new_n909), .A3(new_n940), .ZN(new_n953));
  INV_X1    g528(.A(G1966), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n951), .B1(new_n955), .B2(new_n947), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n949), .B(new_n950), .C1(new_n956), .C2(new_n935), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n943), .A2(new_n945), .A3(new_n909), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n731), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT45), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n942), .A2(new_n960), .ZN(new_n961));
  NOR3_X1   g536(.A1(new_n961), .A2(new_n908), .A3(new_n936), .ZN(new_n962));
  INV_X1    g537(.A(G2078), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(KEYINPUT53), .A3(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT112), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n965), .B1(new_n939), .B2(KEYINPUT45), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n942), .A2(KEYINPUT112), .A3(new_n960), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n833), .A2(KEYINPUT45), .A3(new_n907), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n966), .A2(new_n909), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n969), .A2(G2078), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n959), .B(new_n964), .C1(new_n970), .C2(KEYINPUT53), .ZN(new_n971));
  XNOR2_X1  g546(.A(G301), .B(KEYINPUT54), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n967), .A2(new_n968), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT45), .B1(new_n513), .B2(new_n907), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n909), .B1(new_n975), .B2(KEYINPUT112), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n963), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT53), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n978), .A2(new_n979), .B1(new_n731), .B2(new_n958), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n968), .A2(KEYINPUT53), .A3(new_n963), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n972), .B1(new_n937), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n935), .A2(KEYINPUT51), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n941), .A2(new_n948), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n984), .B1(new_n985), .B2(new_n934), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n957), .A2(new_n973), .A3(new_n983), .A4(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  OAI22_X1  g563(.A1(new_n977), .A2(G1971), .B1(G2090), .B2(new_n958), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n951), .B1(new_n989), .B2(KEYINPUT113), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n530), .A2(G8), .A3(new_n532), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(KEYINPUT55), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT113), .ZN(new_n994));
  OAI221_X1 g569(.A(new_n994), .B1(G2090), .B2(new_n958), .C1(new_n977), .C2(G1971), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n990), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n934), .ZN(new_n997));
  INV_X1    g572(.A(G1976), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n833), .A2(new_n907), .ZN(new_n999));
  OAI221_X1 g574(.A(new_n997), .B1(new_n998), .B2(G288), .C1(new_n936), .C2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT52), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1002), .B1(new_n779), .B2(G1976), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1001), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(G305), .A2(G1981), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT49), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n776), .B1(new_n575), .B2(new_n576), .ZN(new_n1007));
  OR3_X1    g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n936), .A2(new_n999), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1009), .A2(new_n934), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1006), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1008), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT115), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1008), .A2(new_n1010), .A3(KEYINPUT115), .A4(new_n1011), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1004), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n996), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G1971), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n909), .B1(new_n942), .B2(KEYINPUT50), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n944), .B1(new_n833), .B2(new_n907), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AOI22_X1  g596(.A1(new_n969), .A2(new_n1018), .B1(new_n1021), .B2(new_n675), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n992), .B1(new_n1022), .B2(new_n934), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT117), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n992), .B(KEYINPUT117), .C1(new_n1022), .C2(new_n934), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n988), .A2(new_n1017), .A3(KEYINPUT125), .A4(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT125), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1027), .A2(new_n996), .A3(new_n1016), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1029), .B1(new_n1030), .B2(new_n987), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  AOI22_X1  g607(.A1(new_n958), .A2(new_n678), .B1(new_n1009), .B2(new_n711), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT122), .B1(new_n1033), .B2(KEYINPUT60), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1033), .A2(KEYINPUT122), .A3(KEYINPUT60), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n589), .A3(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1033), .A2(KEYINPUT60), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1038), .B1(new_n1034), .B2(new_n588), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT123), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT123), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1037), .A2(new_n1039), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT61), .ZN(new_n1045));
  XNOR2_X1  g620(.A(G299), .B(KEYINPUT57), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n763), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  OAI211_X1 g624(.A(KEYINPUT119), .B(new_n763), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT120), .ZN(new_n1051));
  XOR2_X1   g626(.A(KEYINPUT56), .B(G2072), .Z(new_n1052));
  OAI21_X1  g627(.A(new_n1051), .B1(new_n969), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n974), .ZN(new_n1054));
  INV_X1    g629(.A(new_n976), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1052), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1054), .A2(new_n1055), .A3(KEYINPUT120), .A4(new_n1056), .ZN(new_n1057));
  AOI221_X4 g632(.A(new_n1046), .B1(new_n1049), .B2(new_n1050), .C1(new_n1053), .C2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1046), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1053), .A2(new_n1057), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1059), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1045), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT120), .B1(new_n977), .B2(new_n1056), .ZN(new_n1064));
  NOR4_X1   g639(.A1(new_n974), .A2(new_n976), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1061), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n1046), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1060), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1067), .A2(KEYINPUT61), .A3(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g644(.A(KEYINPUT58), .B(G1341), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1009), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1071), .B1(new_n977), .B2(new_n726), .ZN(new_n1072));
  OR3_X1    g647(.A1(new_n1072), .A2(KEYINPUT59), .A3(new_n553), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT59), .B1(new_n1072), .B2(new_n553), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1063), .A2(new_n1069), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT121), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1063), .A2(new_n1069), .A3(new_n1078), .A4(new_n1075), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1044), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1033), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n589), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1058), .B1(new_n1067), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1032), .B1(new_n1080), .B2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1016), .A2(new_n993), .A3(new_n995), .A4(new_n990), .ZN(new_n1085));
  NOR2_X1   g660(.A1(G288), .A2(G1976), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1086), .B(KEYINPUT116), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1087), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1010), .B1(new_n1088), .B2(new_n1005), .ZN(new_n1089));
  AND2_X1   g664(.A1(new_n1085), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(G301), .B1(new_n980), .B2(new_n964), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT62), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n949), .A2(new_n950), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n947), .B1(new_n962), .B2(G1966), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n935), .B1(new_n1094), .B2(G8), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n986), .B(new_n1092), .C1(new_n1093), .C2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1092), .B1(new_n957), .B2(new_n986), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1091), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1090), .B1(new_n1099), .B2(new_n1030), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n985), .A2(G286), .A3(new_n934), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1027), .A2(new_n996), .A3(new_n1016), .A4(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT63), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n993), .B1(new_n990), .B2(new_n995), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1101), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n1105), .A2(new_n1103), .A3(new_n1106), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1104), .A2(KEYINPUT118), .B1(new_n1017), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT118), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1102), .A2(new_n1109), .A3(new_n1103), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1100), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1084), .A2(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(G290), .B(G1986), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1113), .A2(new_n909), .A3(new_n908), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n930), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT126), .B1(new_n1112), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT126), .ZN(new_n1118));
  AOI211_X1 g693(.A(new_n1118), .B(new_n1115), .C1(new_n1084), .C2(new_n1111), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n933), .B1(new_n1117), .B2(new_n1119), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g695(.A1(G227), .A2(new_n465), .ZN(new_n1122));
  AND4_X1   g696(.A1(new_n634), .A2(new_n849), .A3(new_n669), .A4(new_n1122), .ZN(new_n1123));
  NAND2_X1  g697(.A1(new_n903), .A2(new_n1123), .ZN(G225));
  INV_X1    g698(.A(G225), .ZN(G308));
endmodule


