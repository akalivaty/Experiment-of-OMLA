//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 1 0 1 0 0 1 1 0 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 1 1 0 0 1 1 0 1 1 0 0 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G107), .A2(G264), .ZN(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n207), .B(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  OR2_X1    g0011(.A1(new_n211), .A2(KEYINPUT65), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G116), .A2(G270), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(KEYINPUT65), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  OAI22_X1  g0016(.A1(new_n201), .A2(new_n215), .B1(new_n203), .B2(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n217), .B1(G77), .B2(G244), .ZN(new_n218));
  NAND4_X1  g0018(.A1(new_n212), .A2(new_n213), .A3(new_n214), .A4(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G20), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AND2_X1   g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(KEYINPUT64), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT64), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G20), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n202), .A2(new_n203), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NOR3_X1   g0031(.A1(new_n228), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n220), .A2(G13), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n233), .B(G250), .C1(G257), .C2(G264), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(KEYINPUT0), .Z(new_n235));
  NOR4_X1   g0035(.A1(new_n222), .A2(new_n223), .A3(new_n232), .A4(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G226), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G238), .B(G244), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  INV_X1    g0042(.A(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT67), .B(G250), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n241), .B(new_n246), .ZN(G358));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G87), .B(G97), .Z(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  INV_X1    g0054(.A(KEYINPUT13), .ZN(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n256), .B1(G41), .B2(G45), .ZN(new_n257));
  INV_X1    g0057(.A(G274), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n215), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G232), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G1698), .ZN(new_n263));
  AND2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n261), .B(new_n263), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G97), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(G1), .A3(G13), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n259), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  AND3_X1   g0072(.A1(new_n270), .A2(G238), .A3(new_n257), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n255), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n270), .B1(new_n266), .B2(new_n267), .ZN(new_n276));
  NOR4_X1   g0076(.A1(new_n276), .A2(KEYINPUT13), .A3(new_n273), .A4(new_n259), .ZN(new_n277));
  OAI21_X1  g0077(.A(G169), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT14), .ZN(new_n279));
  INV_X1    g0079(.A(new_n275), .ZN(new_n280));
  INV_X1    g0080(.A(new_n277), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(G179), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT14), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n283), .B(G169), .C1(new_n275), .C2(new_n277), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n279), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT74), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  AND2_X1   g0088(.A1(new_n288), .A2(new_n231), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n228), .A2(G33), .ZN(new_n291));
  INV_X1    g0091(.A(G77), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G20), .A2(G33), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  OAI22_X1  g0094(.A1(new_n291), .A2(new_n292), .B1(new_n201), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n224), .A2(G68), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n290), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT11), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n289), .B1(G1), .B2(new_n224), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n297), .A2(new_n298), .B1(new_n203), .B2(new_n299), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n297), .A2(new_n298), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n296), .A2(new_n256), .A3(G13), .ZN(new_n302));
  XOR2_X1   g0102(.A(new_n302), .B(KEYINPUT12), .Z(new_n303));
  NOR3_X1   g0103(.A1(new_n300), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n279), .A2(KEYINPUT74), .A3(new_n282), .A4(new_n284), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n287), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n280), .A2(new_n281), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G200), .ZN(new_n309));
  INV_X1    g0109(.A(G190), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n304), .B(new_n309), .C1(new_n310), .C2(new_n308), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT75), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n307), .A2(new_n311), .A3(KEYINPUT75), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n215), .A2(G1698), .ZN(new_n317));
  OAI221_X1 g0117(.A(new_n317), .B1(G223), .B2(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G33), .A2(G87), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n271), .ZN(new_n321));
  INV_X1    g0121(.A(new_n259), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n270), .A2(new_n257), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n323), .A2(new_n262), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n321), .A2(new_n322), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G169), .ZN(new_n327));
  INV_X1    g0127(.A(G179), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n327), .B1(new_n328), .B2(new_n326), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT18), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT78), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT16), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n264), .A2(new_n265), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n228), .A2(new_n333), .A3(KEYINPUT7), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT3), .ZN(new_n335));
  INV_X1    g0135(.A(G33), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(KEYINPUT3), .A2(G33), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(new_n224), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT7), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n203), .B1(new_n334), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G58), .A2(G68), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT76), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(KEYINPUT76), .A2(G58), .A3(G68), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(new_n229), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G20), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n293), .A2(G159), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n332), .B1(new_n342), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n228), .A2(new_n333), .A3(new_n340), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n339), .A2(KEYINPUT7), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n352), .A2(new_n353), .A3(G68), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n347), .A2(G20), .B1(G159), .B2(new_n293), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(KEYINPUT16), .A3(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n351), .A2(new_n290), .A3(new_n356), .ZN(new_n357));
  XOR2_X1   g0157(.A(KEYINPUT8), .B(G58), .Z(new_n358));
  NAND2_X1  g0158(.A1(new_n299), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n256), .A2(G13), .A3(G20), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n359), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  AND3_X1   g0162(.A1(new_n357), .A2(KEYINPUT77), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT77), .B1(new_n357), .B2(new_n362), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n329), .B(new_n331), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n330), .A2(KEYINPUT78), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n357), .A2(new_n362), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT77), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n357), .A2(KEYINPUT77), .A3(new_n362), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n366), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n372), .A2(new_n329), .A3(new_n331), .A4(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n326), .A2(G200), .ZN(new_n375));
  XNOR2_X1  g0175(.A(KEYINPUT79), .B(G190), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n321), .A2(new_n322), .A3(new_n325), .A4(new_n376), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n357), .A2(new_n362), .A3(new_n375), .A4(new_n377), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n378), .B(KEYINPUT17), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n367), .A2(new_n374), .A3(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT80), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n367), .A2(new_n374), .A3(KEYINPUT80), .A4(new_n379), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g0184(.A(KEYINPUT15), .B(G87), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n291), .A2(new_n385), .B1(new_n292), .B2(new_n228), .ZN(new_n386));
  INV_X1    g0186(.A(new_n358), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n387), .A2(new_n294), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n290), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n361), .A2(new_n292), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n389), .B(new_n390), .C1(new_n292), .C2(new_n299), .ZN(new_n391));
  XNOR2_X1  g0191(.A(new_n391), .B(KEYINPUT70), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n333), .B1(G232), .B2(new_n260), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(new_n216), .B2(new_n260), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n337), .A2(new_n338), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n395), .B(new_n271), .C1(G107), .C2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G244), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n397), .B(new_n322), .C1(new_n398), .C2(new_n323), .ZN(new_n399));
  INV_X1    g0199(.A(G169), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OR2_X1    g0201(.A1(new_n399), .A2(G179), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n393), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n399), .A2(G200), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n392), .B(new_n404), .C1(new_n310), .C2(new_n399), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT71), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT71), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n403), .A2(new_n405), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G223), .A2(G1698), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n260), .A2(G222), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n396), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n413), .B(new_n271), .C1(G77), .C2(new_n396), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n270), .A2(G226), .A3(new_n257), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(new_n322), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT68), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT68), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n414), .A2(new_n418), .A3(new_n322), .A4(new_n415), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n400), .ZN(new_n422));
  XNOR2_X1  g0222(.A(KEYINPUT64), .B(G20), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n423), .A2(new_n336), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n424), .A2(new_n358), .B1(G150), .B2(new_n293), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n204), .A2(G20), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n289), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT69), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n299), .A2(G50), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n360), .A2(new_n201), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n430), .A2(new_n429), .A3(new_n431), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n428), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n422), .B(new_n434), .C1(G179), .C2(new_n421), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n433), .A2(new_n432), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT9), .B1(new_n437), .B2(new_n427), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT9), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n428), .B(new_n439), .C1(new_n432), .C2(new_n433), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n421), .A2(G200), .ZN(new_n442));
  AOI21_X1  g0242(.A(KEYINPUT72), .B1(new_n420), .B2(G190), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT72), .ZN(new_n444));
  AOI211_X1 g0244(.A(new_n444), .B(new_n310), .C1(new_n417), .C2(new_n419), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n441), .B(new_n442), .C1(new_n443), .C2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT10), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT73), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n447), .B1(new_n442), .B2(new_n448), .ZN(new_n449));
  OR2_X1    g0249(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n446), .A2(new_n449), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n436), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n316), .A2(new_n384), .A3(new_n410), .A4(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT81), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n446), .A2(new_n449), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n446), .A2(new_n449), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n435), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n458), .B1(new_n314), .B2(new_n315), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n459), .A2(KEYINPUT81), .A3(new_n410), .A4(new_n384), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n226), .A2(G20), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n224), .A2(KEYINPUT64), .ZN(new_n464));
  OAI211_X1 g0264(.A(G33), .B(G97), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT19), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n228), .A2(new_n396), .A3(G68), .ZN(new_n468));
  NOR4_X1   g0268(.A1(KEYINPUT82), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT82), .ZN(new_n470));
  NOR2_X1   g0270(.A1(G87), .A2(G97), .ZN(new_n471));
  INV_X1    g0271(.A(G107), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n267), .A2(new_n466), .ZN(new_n474));
  OAI22_X1  g0274(.A1(new_n469), .A2(new_n473), .B1(new_n423), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n467), .A2(new_n468), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT83), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT83), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n467), .A2(new_n475), .A3(new_n478), .A4(new_n468), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n477), .A2(new_n290), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n256), .A2(G33), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n360), .A2(new_n481), .A3(new_n231), .A4(new_n288), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n385), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n385), .A2(new_n361), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n480), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n398), .A2(G1698), .ZN(new_n488));
  OAI221_X1 g0288(.A(new_n488), .B1(G238), .B2(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G33), .A2(G116), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n270), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n256), .A2(G45), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n492), .A2(new_n258), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n270), .A2(G250), .A3(new_n492), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NOR3_X1   g0295(.A1(new_n491), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n328), .ZN(new_n497));
  OR2_X1    g0297(.A1(new_n496), .A2(G169), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n487), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(G200), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n491), .A2(new_n495), .ZN(new_n501));
  INV_X1    g0301(.A(new_n493), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NOR4_X1   g0303(.A1(new_n491), .A2(new_n310), .A3(new_n493), .A4(new_n495), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n483), .A2(G87), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n505), .A2(new_n486), .A3(new_n480), .A4(new_n506), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n499), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n225), .A2(new_n227), .A3(new_n472), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT23), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n224), .A2(G33), .A3(G116), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n472), .A2(KEYINPUT23), .A3(G20), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(KEYINPUT89), .A2(KEYINPUT24), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT22), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n225), .A2(new_n227), .B1(new_n337), .B2(new_n338), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n516), .B1(new_n517), .B2(G87), .ZN(new_n518));
  AND4_X1   g0318(.A1(new_n516), .A2(new_n228), .A3(new_n396), .A4(G87), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n514), .B(new_n515), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(KEYINPUT89), .A2(KEYINPUT24), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n228), .A2(new_n396), .A3(G87), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(KEYINPUT22), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n517), .A2(new_n516), .A3(G87), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n521), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n526), .A2(new_n514), .A3(new_n515), .A4(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n522), .A2(new_n290), .A3(new_n528), .ZN(new_n529));
  OR3_X1    g0329(.A1(new_n360), .A2(KEYINPUT25), .A3(G107), .ZN(new_n530));
  OAI21_X1  g0330(.A(KEYINPUT25), .B1(new_n360), .B2(G107), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n530), .B(new_n531), .C1(new_n472), .C2(new_n482), .ZN(new_n532));
  XNOR2_X1  g0332(.A(new_n532), .B(KEYINPUT90), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n210), .A2(new_n260), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n243), .A2(G1698), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n535), .B(new_n536), .C1(new_n264), .C2(new_n265), .ZN(new_n537));
  INV_X1    g0337(.A(G294), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT91), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT91), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G294), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n539), .A2(new_n541), .A3(G33), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT92), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n537), .A2(KEYINPUT92), .A3(new_n542), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n271), .A3(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(G45), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n548), .A2(G1), .ZN(new_n549));
  NOR2_X1   g0349(.A1(KEYINPUT5), .A2(G41), .ZN(new_n550));
  AND2_X1   g0350(.A1(KEYINPUT5), .A2(G41), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n549), .B(G274), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n549), .B1(new_n551), .B2(new_n550), .ZN(new_n553));
  AND2_X1   g0353(.A1(new_n553), .A2(new_n270), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(G264), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n547), .A2(new_n552), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n400), .ZN(new_n557));
  OR2_X1    g0357(.A1(new_n556), .A2(G179), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n534), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n547), .A2(G190), .A3(new_n552), .A4(new_n555), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n556), .A2(G200), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n529), .A2(new_n560), .A3(new_n533), .A4(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT93), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n562), .A2(new_n563), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n508), .B(new_n559), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n260), .A2(G264), .ZN(new_n567));
  NOR2_X1   g0367(.A1(G257), .A2(G1698), .ZN(new_n568));
  OAI22_X1  g0368(.A1(new_n567), .A2(new_n568), .B1(new_n264), .B2(new_n265), .ZN(new_n569));
  INV_X1    g0369(.A(G303), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n337), .A2(new_n570), .A3(new_n338), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n271), .A3(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n553), .A2(G270), .A3(new_n270), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n572), .A2(new_n552), .A3(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT84), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n572), .A2(new_n573), .A3(KEYINPUT84), .A4(new_n552), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n576), .A2(G169), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(G116), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n360), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n483), .B2(new_n579), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT85), .ZN(new_n582));
  NAND2_X1  g0382(.A1(G33), .A2(G283), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n336), .A2(G97), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n583), .B(new_n584), .C1(new_n463), .C2(new_n464), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n288), .A2(new_n231), .B1(G20), .B2(new_n579), .ZN(new_n586));
  AND3_X1   g0386(.A1(new_n585), .A2(KEYINPUT20), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(KEYINPUT20), .B1(new_n585), .B2(new_n586), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n581), .B(new_n582), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n585), .A2(new_n586), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT20), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n585), .A2(KEYINPUT20), .A3(new_n586), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n582), .B1(new_n595), .B2(new_n581), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n578), .B1(new_n590), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT21), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(KEYINPUT86), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n581), .B1(new_n587), .B2(new_n588), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT85), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n589), .ZN(new_n603));
  OR2_X1    g0403(.A1(new_n574), .A2(new_n328), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n576), .A2(new_n577), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n599), .A2(G169), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n597), .A2(new_n600), .B1(new_n603), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n576), .A2(G200), .A3(new_n577), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n609), .A2(new_n602), .A3(new_n589), .ZN(new_n610));
  INV_X1    g0410(.A(new_n376), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n611), .B1(new_n576), .B2(new_n577), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(KEYINPUT87), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n609), .A2(new_n602), .A3(new_n589), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT87), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n615), .A2(new_n616), .A3(new_n612), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n608), .B1(new_n614), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT88), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n608), .B(KEYINPUT88), .C1(new_n614), .C2(new_n617), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT6), .ZN(new_n623));
  INV_X1    g0423(.A(G97), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n624), .A2(new_n472), .ZN(new_n625));
  NOR2_X1   g0425(.A1(G97), .A2(G107), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n472), .A2(KEYINPUT6), .A3(G97), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n228), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n294), .A2(new_n292), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n334), .A2(new_n341), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n630), .B(new_n632), .C1(new_n633), .C2(new_n472), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n634), .A2(new_n290), .B1(new_n624), .B2(new_n361), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT4), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n636), .A2(G1698), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n637), .B(G244), .C1(new_n265), .C2(new_n264), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n398), .B1(new_n337), .B2(new_n338), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n638), .B(new_n583), .C1(new_n639), .C2(KEYINPUT4), .ZN(new_n640));
  OAI21_X1  g0440(.A(G250), .B1(new_n264), .B2(new_n265), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n260), .B1(new_n641), .B2(KEYINPUT4), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n271), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n554), .A2(G257), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(new_n552), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(G200), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n483), .A2(G97), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n643), .A2(G190), .A3(new_n552), .A4(new_n644), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n635), .A2(new_n646), .A3(new_n647), .A4(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n361), .A2(new_n624), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n472), .B1(new_n334), .B2(new_n341), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n651), .A2(new_n631), .A3(new_n629), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n650), .B(new_n647), .C1(new_n652), .C2(new_n289), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n645), .A2(new_n400), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n643), .A2(new_n328), .A3(new_n552), .A4(new_n644), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n649), .A2(new_n656), .ZN(new_n657));
  NOR4_X1   g0457(.A1(new_n462), .A2(new_n566), .A3(new_n622), .A4(new_n657), .ZN(G372));
  NAND2_X1  g0458(.A1(new_n329), .A2(new_n368), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n659), .B(new_n330), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n311), .A2(new_n393), .A3(new_n401), .A4(new_n402), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n307), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n661), .B1(new_n663), .B2(new_n379), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n456), .A2(new_n457), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n435), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n562), .B(new_n563), .ZN(new_n668));
  INV_X1    g0468(.A(new_n657), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n608), .A2(new_n559), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n668), .A2(new_n669), .A3(new_n508), .A4(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n499), .ZN(new_n672));
  INV_X1    g0472(.A(new_n656), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n673), .A2(new_n499), .A3(new_n507), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n673), .A2(new_n499), .A3(new_n507), .A4(KEYINPUT26), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n672), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n671), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n667), .B1(new_n462), .B2(new_n680), .ZN(G369));
  INV_X1    g0481(.A(G13), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n423), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n256), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(G213), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G343), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n603), .A2(new_n689), .ZN(new_n690));
  MUX2_X1   g0490(.A(new_n622), .B(new_n608), .S(new_n690), .Z(new_n691));
  XOR2_X1   g0491(.A(new_n691), .B(KEYINPUT94), .Z(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G330), .ZN(new_n693));
  INV_X1    g0493(.A(new_n559), .ZN(new_n694));
  INV_X1    g0494(.A(new_n689), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n534), .A2(new_n689), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n668), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n696), .B1(new_n698), .B2(new_n694), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n693), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n699), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n608), .A2(new_n689), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n696), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT95), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n704), .A2(KEYINPUT95), .A3(new_n696), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n701), .A2(new_n709), .ZN(G399));
  INV_X1    g0510(.A(new_n233), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT96), .ZN(new_n712));
  OR3_X1    g0512(.A1(new_n711), .A2(new_n712), .A3(G41), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n712), .B1(new_n711), .B2(G41), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OR3_X1    g0515(.A1(new_n469), .A2(new_n473), .A3(G116), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n715), .A2(new_n717), .A3(G1), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n230), .B2(new_n715), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT28), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n689), .B1(new_n671), .B2(new_n678), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT29), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n657), .A2(KEYINPUT99), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT99), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n649), .A2(new_n725), .A3(new_n656), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n727), .A2(new_n668), .A3(new_n508), .A4(new_n670), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n499), .A2(KEYINPUT98), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n499), .A2(KEYINPUT98), .ZN(new_n730));
  AOI22_X1  g0530(.A1(new_n676), .A2(new_n677), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n689), .B1(new_n728), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n723), .B1(new_n722), .B2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT30), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n645), .A2(new_n604), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n496), .A2(new_n555), .A3(new_n547), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n738), .A2(KEYINPUT97), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n736), .A2(new_n737), .ZN(new_n740));
  INV_X1    g0540(.A(new_n645), .ZN(new_n741));
  NOR4_X1   g0541(.A1(new_n741), .A2(new_n605), .A3(G179), .A4(new_n496), .ZN(new_n742));
  AOI22_X1  g0542(.A1(new_n740), .A2(KEYINPUT30), .B1(new_n742), .B2(new_n556), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n738), .A2(KEYINPUT97), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n739), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n745), .A2(new_n689), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n620), .A2(new_n621), .ZN(new_n747));
  INV_X1    g0547(.A(new_n566), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n747), .A2(new_n748), .A3(new_n669), .A4(new_n695), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n746), .B1(new_n749), .B2(KEYINPUT31), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT31), .ZN(new_n751));
  AOI211_X1 g0551(.A(new_n751), .B(new_n695), .C1(new_n743), .C2(new_n738), .ZN(new_n752));
  OAI21_X1  g0552(.A(G330), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  AND2_X1   g0553(.A1(new_n734), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n720), .B1(new_n754), .B2(G1), .ZN(G364));
  NAND2_X1  g0555(.A1(new_n683), .A2(G45), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n715), .A2(G1), .A3(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n758), .B1(new_n692), .B2(G330), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n759), .B1(G330), .B2(new_n692), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n711), .A2(new_n396), .ZN(new_n761));
  INV_X1    g0561(.A(new_n230), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(new_n548), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n761), .B(new_n763), .C1(new_n250), .C2(new_n548), .ZN(new_n764));
  INV_X1    g0564(.A(G355), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n396), .A2(new_n233), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n764), .B1(G116), .B2(new_n233), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G13), .A2(G33), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n231), .B1(G20), .B2(new_n400), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n767), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n423), .A2(new_n310), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT100), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n775), .A2(G179), .A3(G200), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G159), .ZN(new_n777));
  XOR2_X1   g0577(.A(new_n777), .B(KEYINPUT32), .Z(new_n778));
  NOR3_X1   g0578(.A1(new_n775), .A2(G179), .A3(new_n500), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n228), .A2(new_n328), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n781), .A2(new_n500), .A3(new_n376), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n780), .A2(new_n472), .B1(new_n782), .B2(new_n202), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n781), .A2(G200), .A3(new_n376), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n781), .A2(new_n310), .A3(G200), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n201), .A2(new_n784), .B1(new_n785), .B2(new_n203), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n500), .A2(G179), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n787), .A2(G20), .A3(G190), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G87), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n310), .A2(G179), .A3(G200), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n228), .A2(new_n791), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n790), .B(new_n396), .C1(new_n624), .C2(new_n792), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n783), .A2(new_n786), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n781), .A2(new_n500), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(G190), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n778), .B(new_n794), .C1(new_n292), .C2(new_n797), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n798), .B(KEYINPUT101), .Z(new_n799));
  NAND2_X1  g0599(.A1(new_n539), .A2(new_n541), .ZN(new_n800));
  INV_X1    g0600(.A(G326), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n333), .B1(new_n800), .B2(new_n792), .C1(new_n784), .C2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n782), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G322), .ZN(new_n804));
  XNOR2_X1  g0604(.A(KEYINPUT103), .B(KEYINPUT33), .ZN(new_n805));
  INV_X1    g0605(.A(G317), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n805), .B(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G311), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n804), .B1(new_n785), .B2(new_n807), .C1(new_n797), .C2(new_n808), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n802), .B(new_n809), .C1(G283), .C2(new_n779), .ZN(new_n810));
  INV_X1    g0610(.A(G329), .ZN(new_n811));
  XOR2_X1   g0611(.A(new_n776), .B(KEYINPUT102), .Z(new_n812));
  OAI221_X1 g0612(.A(new_n810), .B1(new_n570), .B2(new_n788), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n799), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n757), .B1(new_n814), .B2(new_n771), .ZN(new_n815));
  INV_X1    g0615(.A(new_n770), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n773), .B(new_n815), .C1(new_n692), .C2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n760), .A2(new_n817), .ZN(G396));
  NOR2_X1   g0618(.A1(new_n403), .A2(new_n689), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n405), .B1(new_n392), .B2(new_n695), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n819), .B1(new_n403), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(new_n721), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n753), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n757), .ZN(new_n825));
  INV_X1    g0625(.A(G132), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n396), .B1(new_n812), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT106), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n827), .A2(new_n828), .ZN(new_n830));
  INV_X1    g0630(.A(new_n785), .ZN(new_n831));
  AOI22_X1  g0631(.A1(G143), .A2(new_n803), .B1(new_n831), .B2(G150), .ZN(new_n832));
  INV_X1    g0632(.A(G137), .ZN(new_n833));
  INV_X1    g0633(.A(G159), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n832), .B1(new_n833), .B2(new_n784), .C1(new_n834), .C2(new_n797), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT34), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n779), .A2(G68), .ZN(new_n838));
  INV_X1    g0638(.A(new_n792), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(G58), .ZN(new_n840));
  AND3_X1   g0640(.A1(new_n837), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n830), .B(new_n841), .C1(new_n836), .C2(new_n835), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n829), .B(new_n842), .C1(G50), .C2(new_n789), .ZN(new_n843));
  INV_X1    g0643(.A(new_n812), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n844), .A2(G311), .B1(G97), .B2(new_n839), .ZN(new_n845));
  INV_X1    g0645(.A(new_n784), .ZN(new_n846));
  AOI22_X1  g0646(.A1(G116), .A2(new_n796), .B1(new_n846), .B2(G303), .ZN(new_n847));
  INV_X1    g0647(.A(G283), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n847), .B1(new_n848), .B2(new_n785), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT104), .Z(new_n850));
  OAI221_X1 g0650(.A(new_n333), .B1(new_n472), .B2(new_n788), .C1(new_n782), .C2(new_n538), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(new_n779), .B2(G87), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n845), .A2(new_n850), .A3(new_n852), .ZN(new_n853));
  XOR2_X1   g0653(.A(new_n853), .B(KEYINPUT105), .Z(new_n854));
  OAI21_X1  g0654(.A(new_n771), .B1(new_n843), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n822), .A2(new_n768), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n771), .A2(new_n768), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n292), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n855), .A2(new_n758), .A3(new_n856), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n825), .A2(new_n859), .ZN(G384));
  NAND2_X1  g0660(.A1(new_n305), .A2(new_n689), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n312), .B(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n862), .A2(new_n822), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n354), .A2(new_n355), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n332), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n865), .A2(new_n290), .A3(new_n356), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n687), .B1(new_n866), .B2(new_n362), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n380), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n329), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n869), .A2(new_n687), .B1(new_n362), .B2(new_n866), .ZN(new_n870));
  INV_X1    g0670(.A(new_n378), .ZN(new_n871));
  OAI21_X1  g0671(.A(KEYINPUT37), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n687), .ZN(new_n873));
  OAI22_X1  g0673(.A1(new_n363), .A2(new_n364), .B1(new_n329), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT37), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n874), .A2(new_n875), .A3(new_n378), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n868), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT38), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n868), .A2(KEYINPUT38), .A3(new_n877), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n746), .A2(KEYINPUT31), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n863), .B(new_n882), .C1(new_n750), .C2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT40), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n660), .A2(new_n379), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n687), .B1(new_n370), .B2(new_n371), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n659), .A2(new_n378), .ZN(new_n890));
  OAI21_X1  g0690(.A(KEYINPUT37), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n876), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n879), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n885), .B1(new_n894), .B2(new_n881), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n895), .B(new_n863), .C1(new_n750), .C2(new_n883), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n886), .A2(new_n896), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n750), .A2(new_n883), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n461), .A2(new_n898), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n897), .B(new_n899), .Z(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(G330), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n901), .B(KEYINPUT109), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n880), .A2(KEYINPUT39), .A3(new_n881), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT39), .ZN(new_n904));
  AOI221_X4 g0704(.A(new_n879), .B1(new_n872), .B2(new_n876), .C1(new_n380), .C2(new_n867), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT38), .B1(new_n889), .B2(new_n892), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n307), .A2(new_n689), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n903), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n821), .A2(new_n679), .A3(new_n695), .ZN(new_n910));
  INV_X1    g0710(.A(new_n819), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n862), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n912), .A2(new_n882), .A3(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n660), .A2(new_n873), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n909), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(KEYINPUT108), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT108), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n909), .A2(new_n914), .A3(new_n919), .A4(new_n916), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n666), .B1(new_n461), .B2(new_n733), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n921), .B(new_n922), .Z(new_n923));
  XNOR2_X1  g0723(.A(new_n902), .B(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n256), .B2(new_n683), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n627), .A2(new_n628), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n579), .B1(new_n926), .B2(KEYINPUT35), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n228), .A2(new_n231), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n927), .B(new_n928), .C1(KEYINPUT35), .C2(new_n926), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT36), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n762), .A2(G77), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n345), .A2(new_n346), .ZN(new_n932));
  OAI22_X1  g0732(.A1(new_n931), .A2(new_n932), .B1(G50), .B2(new_n203), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n933), .A2(G1), .A3(new_n682), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT107), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n925), .A2(new_n930), .A3(new_n935), .ZN(G367));
  NAND3_X1  g0736(.A1(new_n480), .A2(new_n486), .A3(new_n506), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n689), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n508), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n499), .A2(new_n938), .ZN(new_n940));
  OAI21_X1  g0740(.A(KEYINPUT110), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(KEYINPUT110), .B2(new_n940), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n689), .A2(new_n653), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n727), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n673), .A2(new_n689), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  OR3_X1    g0748(.A1(new_n704), .A2(KEYINPUT42), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n656), .B1(new_n945), .B2(new_n559), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n695), .ZN(new_n951));
  OAI21_X1  g0751(.A(KEYINPUT42), .B1(new_n704), .B2(new_n948), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n949), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n943), .B(new_n953), .C1(new_n701), .C2(new_n948), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n953), .A2(new_n943), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n700), .A2(new_n956), .A3(new_n947), .ZN(new_n957));
  AND3_X1   g0757(.A1(new_n954), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n955), .B1(new_n954), .B2(new_n957), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n715), .B(KEYINPUT41), .Z(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n948), .B1(new_n707), .B2(new_n708), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n963), .B(KEYINPUT45), .Z(new_n964));
  NAND3_X1  g0764(.A1(new_n707), .A2(new_n708), .A3(new_n948), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n965), .A2(KEYINPUT44), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(KEYINPUT44), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n700), .B1(new_n964), .B2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT111), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n704), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n692), .A2(G330), .A3(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n971), .B1(new_n692), .B2(G330), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n973), .A2(new_n974), .B1(new_n702), .B2(new_n703), .ZN(new_n975));
  INV_X1    g0775(.A(new_n974), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n702), .A2(new_n703), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n976), .A2(new_n977), .A3(new_n972), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n963), .B(KEYINPUT45), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n980), .A2(new_n701), .A3(new_n967), .A4(new_n966), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n969), .A2(new_n979), .A3(new_n754), .A4(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n962), .B1(new_n982), .B2(new_n754), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n756), .A2(G1), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n960), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G283), .A2(new_n796), .B1(new_n846), .B2(G311), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n800), .B2(new_n785), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n789), .A2(G116), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT46), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n396), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n990), .B1(new_n989), .B2(new_n988), .C1(new_n570), .C2(new_n782), .ZN(new_n991));
  XOR2_X1   g0791(.A(KEYINPUT112), .B(G317), .Z(new_n992));
  AOI21_X1  g0792(.A(new_n991), .B1(new_n776), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n624), .B2(new_n780), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n987), .B(new_n994), .C1(G107), .C2(new_n839), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n831), .A2(G159), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n839), .A2(G68), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n333), .B1(new_n789), .B2(G58), .ZN(new_n998));
  INV_X1    g0798(.A(new_n776), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n997), .B(new_n998), .C1(new_n999), .C2(new_n833), .ZN(new_n1000));
  INV_X1    g0800(.A(G143), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n780), .A2(new_n292), .B1(new_n1001), .B2(new_n784), .ZN(new_n1002));
  INV_X1    g0802(.A(G150), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n797), .A2(new_n201), .B1(new_n1003), .B2(new_n782), .ZN(new_n1004));
  NOR3_X1   g0804(.A1(new_n1000), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n995), .B1(new_n996), .B2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT47), .Z(new_n1007));
  AOI21_X1  g0807(.A(new_n757), .B1(new_n1007), .B2(new_n771), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n761), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n772), .B1(new_n233), .B2(new_n385), .C1(new_n246), .C2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1008), .B(new_n1010), .C1(new_n816), .C2(new_n942), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n985), .A2(new_n1011), .ZN(G387));
  OR2_X1    g0812(.A1(new_n979), .A2(new_n754), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n715), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n979), .A2(new_n754), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n333), .B1(new_n780), .B2(new_n579), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G303), .A2(new_n796), .B1(new_n846), .B2(G322), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n808), .B2(new_n785), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(new_n803), .B2(new_n992), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT48), .Z(new_n1021));
  OAI221_X1 g0821(.A(new_n1021), .B1(new_n848), .B2(new_n792), .C1(new_n800), .C2(new_n788), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT49), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1017), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1024), .B1(new_n1023), .B2(new_n1022), .C1(new_n801), .C2(new_n999), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n797), .A2(new_n203), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n792), .A2(new_n385), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n396), .B1(new_n788), .B2(new_n292), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1027), .B(new_n1028), .C1(new_n776), .C2(G150), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G159), .A2(new_n846), .B1(new_n831), .B2(new_n358), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n779), .A2(G97), .B1(G50), .B2(new_n803), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1025), .B1(new_n1026), .B2(new_n1032), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n241), .A2(new_n548), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT113), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1009), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n358), .A2(new_n201), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1037), .A2(KEYINPUT50), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(G68), .A2(G77), .ZN(new_n1039));
  AOI21_X1  g0839(.A(G45), .B1(new_n1037), .B2(KEYINPUT50), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n717), .A2(new_n1038), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1036), .B(new_n1041), .C1(new_n1035), .C2(new_n1034), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(G107), .B2(new_n233), .C1(new_n717), .C2(new_n766), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n1033), .A2(new_n771), .B1(new_n772), .B2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1044), .B(new_n758), .C1(new_n702), .C2(new_n816), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(new_n979), .B2(new_n984), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1016), .A2(new_n1047), .ZN(G393));
  NOR2_X1   g0848(.A1(new_n792), .A2(new_n292), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n396), .B1(new_n203), .B2(new_n788), .C1(new_n797), .C2(new_n387), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(G50), .C2(new_n831), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n1003), .A2(new_n784), .B1(new_n782), .B2(new_n834), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT51), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1051), .B(new_n1053), .C1(new_n209), .C2(new_n780), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n999), .A2(new_n1001), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n788), .A2(new_n848), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n333), .B1(new_n579), .B2(new_n792), .C1(new_n797), .C2(new_n538), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(G303), .B2(new_n831), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n808), .A2(new_n782), .B1(new_n784), .B2(new_n806), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT52), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G107), .A2(new_n779), .B1(new_n776), .B2(G322), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1058), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n1054), .A2(new_n1055), .B1(new_n1056), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n757), .B1(new_n1063), .B2(new_n771), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n772), .B1(new_n624), .B2(new_n233), .C1(new_n253), .C2(new_n1009), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1064), .B(new_n1065), .C1(new_n816), .C2(new_n947), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n969), .A2(new_n981), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n984), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n715), .B1(new_n1067), .B2(new_n1015), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1069), .B1(new_n982), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(G390));
  NAND2_X1  g0872(.A1(new_n789), .A2(G150), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n1073), .A2(KEYINPUT53), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n396), .B1(new_n792), .B2(new_n834), .C1(new_n1073), .C2(KEYINPUT53), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(G132), .B2(new_n803), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n779), .A2(G50), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n831), .A2(G137), .ZN(new_n1078));
  XOR2_X1   g0878(.A(KEYINPUT54), .B(G143), .Z(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT117), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n796), .A2(new_n1080), .B1(new_n846), .B2(G128), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .A4(new_n1081), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1074), .B(new_n1082), .C1(new_n844), .C2(G125), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n396), .B(new_n1049), .C1(new_n796), .C2(G97), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n790), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G116), .A2(new_n803), .B1(new_n846), .B2(G283), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n838), .B(new_n1086), .C1(new_n472), .C2(new_n785), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n1085), .B(new_n1087), .C1(new_n844), .C2(G294), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n1083), .A2(new_n1088), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n1089), .A2(new_n771), .B1(new_n387), .B2(new_n857), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n903), .A2(new_n907), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n758), .B(new_n1090), .C1(new_n1092), .C2(new_n769), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n821), .A2(G330), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n913), .B(new_n1094), .C1(new_n750), .C2(new_n752), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n908), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n819), .B1(new_n721), .B2(new_n821), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1096), .B1(new_n1097), .B2(new_n862), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n728), .A2(new_n731), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n820), .A2(new_n403), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1099), .A2(new_n695), .A3(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n862), .B1(new_n1101), .B2(new_n911), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1096), .B1(new_n905), .B2(new_n906), .ZN(new_n1103));
  OAI21_X1  g0903(.A(KEYINPUT114), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n908), .B1(new_n894), .B2(new_n881), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT114), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n819), .B1(new_n732), .B2(new_n1100), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1105), .B(new_n1106), .C1(new_n1107), .C2(new_n862), .ZN(new_n1108));
  AOI221_X4 g0908(.A(new_n1095), .B1(new_n1091), .B2(new_n1098), .C1(new_n1104), .C2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n913), .B(new_n1094), .C1(new_n750), .C2(new_n883), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1104), .A2(new_n1108), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1091), .A2(new_n1098), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1109), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1093), .B1(new_n1115), .B2(new_n1068), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT116), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n461), .A2(new_n898), .A3(G330), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n922), .A2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1094), .B1(new_n750), .B2(new_n752), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n862), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n1110), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n912), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1094), .B1(new_n750), .B2(new_n883), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n862), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1126), .A2(new_n1107), .A3(new_n1095), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1120), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1095), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1112), .A2(new_n1113), .A3(new_n1129), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n1104), .A2(new_n1108), .B1(new_n1091), .B2(new_n1098), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1130), .B1(new_n1131), .B2(new_n1111), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1128), .A2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(KEYINPUT115), .B1(new_n1133), .B2(new_n1014), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT115), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1135), .B(new_n715), .C1(new_n1128), .C2(new_n1132), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n1126), .A2(new_n1107), .A3(new_n1095), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1097), .B1(new_n1122), .B2(new_n1110), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n922), .B(new_n1119), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1115), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1118), .B1(new_n1137), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1014), .B1(new_n1115), .B2(new_n1140), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n1135), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1133), .A2(KEYINPUT115), .A3(new_n1014), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1144), .A2(new_n1118), .A3(new_n1141), .A4(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1117), .B1(new_n1142), .B2(new_n1147), .ZN(G378));
  NOR2_X1   g0948(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n922), .B(new_n1119), .C1(new_n1115), .C2(new_n1149), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n886), .A2(KEYINPUT122), .A3(G330), .A4(new_n896), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n921), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n452), .B(KEYINPUT55), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n434), .A2(new_n873), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n458), .B(KEYINPUT55), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1155), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1156), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT122), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n886), .A2(G330), .A3(new_n896), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1165), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1151), .A2(new_n920), .A3(new_n918), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n1153), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1168), .B1(new_n1153), .B2(new_n1169), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1150), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT57), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1168), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1169), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1151), .B1(new_n920), .B2(new_n918), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1175), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1153), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1180), .A2(KEYINPUT57), .A3(new_n1150), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1174), .A2(new_n1181), .A3(new_n1014), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n484), .A2(new_n796), .B1(new_n803), .B2(G107), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n624), .B2(new_n785), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n779), .A2(G58), .ZN(new_n1185));
  AOI211_X1 g0985(.A(G41), .B(new_n396), .C1(new_n789), .C2(G77), .ZN(new_n1186));
  OR2_X1    g0986(.A1(new_n1186), .A2(KEYINPUT118), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(KEYINPUT118), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1185), .A2(new_n997), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1184), .B(new_n1189), .C1(new_n844), .C2(G283), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n579), .B2(new_n784), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT58), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n201), .B1(new_n264), .B2(G41), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(G128), .A2(new_n803), .B1(new_n1080), .B2(new_n789), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n1194), .B(KEYINPUT119), .Z(new_n1195));
  OAI22_X1  g0995(.A1(new_n785), .A2(new_n826), .B1(new_n1003), .B2(new_n792), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(G125), .B2(new_n846), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1195), .B(new_n1197), .C1(new_n833), .C2(new_n797), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT59), .Z(new_n1199));
  AOI21_X1  g0999(.A(G41), .B1(new_n776), .B2(G124), .ZN(new_n1200));
  AOI21_X1  g1000(.A(G33), .B1(new_n779), .B2(G159), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1192), .A2(new_n1193), .A3(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT120), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n757), .B1(new_n1204), .B2(new_n771), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1165), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1205), .B1(new_n1206), .B2(new_n769), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(new_n201), .B2(new_n857), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n1180), .B2(new_n984), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1182), .A2(new_n1209), .ZN(G375));
  NAND2_X1  g1010(.A1(new_n1149), .A2(new_n1120), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1211), .A2(new_n961), .A3(new_n1140), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G150), .A2(new_n796), .B1(new_n831), .B2(new_n1080), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n833), .B2(new_n782), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n333), .B1(new_n839), .B2(G50), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1185), .B(new_n1215), .C1(new_n826), .C2(new_n784), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1214), .B(new_n1216), .C1(new_n844), .C2(G128), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n834), .B2(new_n788), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n333), .B1(new_n624), .B2(new_n788), .C1(new_n797), .C2(new_n472), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G77), .B2(new_n779), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n579), .A2(new_n785), .B1(new_n782), .B2(new_n848), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1027), .B(new_n1221), .C1(G294), .C2(new_n846), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1220), .B(new_n1222), .C1(new_n812), .C2(new_n570), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1218), .A2(new_n1223), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1224), .A2(new_n771), .B1(new_n203), .B2(new_n857), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n862), .A2(new_n768), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n1225), .A2(new_n758), .A3(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1149), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1227), .B1(new_n1228), .B2(new_n984), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1212), .A2(new_n1229), .ZN(G381));
  AND3_X1   g1030(.A1(new_n985), .A2(new_n1011), .A3(new_n1071), .ZN(new_n1231));
  INV_X1    g1031(.A(G396), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1016), .A2(new_n1232), .A3(new_n1047), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1144), .A2(new_n1141), .A3(new_n1145), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n1117), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(G375), .A2(new_n1236), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(G381), .A2(G384), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1231), .A2(new_n1234), .A3(new_n1237), .A4(new_n1238), .ZN(G407));
  NAND2_X1  g1039(.A1(new_n688), .A2(G213), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1237), .A2(new_n1241), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1242), .B(KEYINPUT123), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1243), .A2(G213), .A3(G407), .ZN(G409));
  NAND2_X1  g1044(.A1(G393), .A2(G396), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1233), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1071), .B1(new_n985), .B2(new_n1011), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1247), .B1(new_n1231), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(G387), .A2(G390), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n985), .A2(new_n1011), .A3(new_n1071), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1250), .A2(new_n1251), .A3(new_n1246), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1249), .A2(new_n1252), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(new_n1253), .B(KEYINPUT126), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT61), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1180), .A2(new_n961), .A3(new_n1150), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1236), .B1(new_n1209), .B2(new_n1256), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(G378), .A2(KEYINPUT124), .A3(new_n1209), .A4(new_n1182), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT124), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1235), .A2(KEYINPUT116), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1116), .B1(new_n1260), .B2(new_n1146), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1259), .B1(G375), .B2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1257), .B1(new_n1258), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT60), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1014), .B(new_n1140), .C1(new_n1211), .C2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(KEYINPUT60), .B1(new_n1149), .B2(new_n1120), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1229), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1267), .A2(new_n859), .A3(new_n825), .ZN(new_n1268));
  OAI211_X1 g1068(.A(G384), .B(new_n1229), .C1(new_n1265), .C2(new_n1266), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NOR3_X1   g1070(.A1(new_n1263), .A2(new_n1241), .A3(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT62), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1255), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1257), .ZN(new_n1274));
  AND2_X1   g1074(.A1(new_n1182), .A2(new_n1209), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT124), .B1(new_n1275), .B2(G378), .ZN(new_n1276));
  NOR3_X1   g1076(.A1(G375), .A2(new_n1261), .A3(new_n1259), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1274), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1270), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1278), .A2(new_n1240), .A3(new_n1279), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1270), .A2(G2897), .A3(new_n1241), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1270), .B1(G2897), .B2(new_n1241), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1283), .B1(new_n1263), .B2(new_n1241), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT62), .B1(new_n1280), .B2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1254), .B1(new_n1273), .B2(new_n1285), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1249), .A2(new_n1252), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n1255), .B(new_n1287), .C1(new_n1271), .C2(KEYINPUT63), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT63), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1289), .B1(new_n1280), .B2(new_n1284), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT125), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(new_n1288), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1283), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1293), .B1(new_n1278), .B2(new_n1240), .ZN(new_n1294));
  OAI21_X1  g1094(.A(KEYINPUT63), .B1(new_n1294), .B2(new_n1271), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1249), .A2(new_n1252), .A3(new_n1255), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1296), .B1(new_n1280), .B2(new_n1289), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT125), .B1(new_n1295), .B2(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1286), .B1(new_n1292), .B2(new_n1298), .ZN(G405));
  INV_X1    g1099(.A(new_n1236), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(G375), .A2(new_n1300), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1301), .B(KEYINPUT127), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1258), .A2(new_n1262), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  XNOR2_X1  g1104(.A(new_n1304), .B(new_n1279), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(new_n1305), .B(new_n1253), .ZN(G402));
endmodule


