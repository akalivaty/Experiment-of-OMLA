//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 1 0 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 0 1 1 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 1 0 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n803, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1051, new_n1052, new_n1053;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  INV_X1    g001(.A(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(KEYINPUT83), .B(KEYINPUT31), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G228gat), .ZN(new_n208));
  INV_X1    g007(.A(G233gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G218gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G211gat), .ZN(new_n212));
  INV_X1    g011(.A(G211gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G218gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT73), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G197gat), .B(G204gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(G211gat), .B(G218gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n218), .B1(new_n219), .B2(KEYINPUT73), .ZN(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT72), .B(G211gat), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT22), .B1(new_n221), .B2(G218gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n217), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT29), .ZN(new_n224));
  AND2_X1   g023(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n226));
  OAI21_X1  g025(.A(G218gat), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT22), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n215), .A2(new_n216), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n219), .A2(KEYINPUT73), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n229), .A2(new_n230), .A3(new_n231), .A4(new_n218), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n223), .A2(new_n224), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(G155gat), .A2(G162gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT2), .ZN(new_n237));
  OR2_X1    g036(.A1(G141gat), .A2(G148gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(G141gat), .A2(G148gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n237), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT79), .ZN(new_n241));
  XNOR2_X1  g040(.A(G155gat), .B(G162gat), .ZN(new_n242));
  AND3_X1   g041(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n242), .B1(new_n240), .B2(new_n241), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n235), .A2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n234), .B1(new_n243), .B2(new_n244), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT80), .ZN(new_n248));
  XNOR2_X1  g047(.A(G141gat), .B(G148gat), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT2), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n250), .B1(G155gat), .B2(G162gat), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n241), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n242), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT80), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n256), .A2(new_n257), .A3(new_n234), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT29), .B1(new_n248), .B2(new_n258), .ZN(new_n259));
  AND3_X1   g058(.A1(new_n223), .A2(KEYINPUT74), .A3(new_n232), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT74), .B1(new_n223), .B2(new_n232), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n210), .B(new_n246), .C1(new_n259), .C2(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n256), .B1(new_n233), .B2(new_n234), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n257), .B1(new_n256), .B2(new_n234), .ZN(new_n265));
  AOI211_X1 g064(.A(KEYINPUT80), .B(KEYINPUT3), .C1(new_n254), .C2(new_n255), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n224), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n232), .ZN(new_n268));
  INV_X1    g067(.A(G197gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(G204gat), .ZN(new_n270));
  INV_X1    g069(.A(G204gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(G197gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n273), .B1(new_n216), .B2(new_n215), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n231), .B1(new_n274), .B2(new_n229), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n268), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n264), .B1(new_n267), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n263), .B1(new_n278), .B2(new_n210), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n207), .B1(new_n279), .B2(G22gat), .ZN(new_n280));
  INV_X1    g079(.A(G22gat), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n263), .B(new_n281), .C1(new_n278), .C2(new_n210), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT84), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n246), .B1(new_n259), .B2(new_n276), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n284), .B1(new_n208), .B2(new_n209), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT84), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n285), .A2(new_n286), .A3(new_n281), .A4(new_n263), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n280), .A2(new_n283), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT85), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n280), .A2(new_n283), .A3(KEYINPUT85), .A4(new_n287), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n279), .A2(G22gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(new_n282), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(new_n207), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G127gat), .B(G134gat), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G113gat), .B(G120gat), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n298), .B1(KEYINPUT1), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n299), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT1), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(new_n302), .A3(new_n297), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n254), .A2(KEYINPUT3), .A3(new_n255), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n304), .B(new_n305), .C1(new_n265), .C2(new_n266), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT4), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n307), .B1(new_n245), .B2(new_n304), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n300), .A2(new_n303), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n309), .A2(new_n256), .A3(KEYINPUT4), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT5), .ZN(new_n312));
  NAND2_X1  g111(.A1(G225gat), .A2(G233gat), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n306), .A2(new_n311), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n305), .A2(new_n304), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n315), .B1(new_n248), .B2(new_n258), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n308), .A2(new_n310), .ZN(new_n317));
  INV_X1    g116(.A(new_n313), .ZN(new_n318));
  NOR3_X1   g117(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n256), .B(new_n304), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT5), .B1(new_n320), .B2(new_n313), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n314), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G1gat), .B(G29gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n323), .B(KEYINPUT0), .ZN(new_n324));
  XNOR2_X1  g123(.A(G57gat), .B(G85gat), .ZN(new_n325));
  XOR2_X1   g124(.A(new_n324), .B(new_n325), .Z(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n322), .A2(new_n327), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n314), .B(new_n326), .C1(new_n319), .C2(new_n321), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT81), .B(KEYINPUT6), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT82), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n328), .A2(KEYINPUT82), .A3(new_n329), .A4(new_n330), .ZN(new_n334));
  INV_X1    g133(.A(new_n330), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n322), .A2(new_n327), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n333), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT68), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g139(.A(KEYINPUT68), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AND2_X1   g141(.A1(G169gat), .A2(G176gat), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT26), .ZN(new_n344));
  NOR2_X1   g143(.A1(G169gat), .A2(G176gat), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(G183gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT27), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT27), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(G183gat), .ZN(new_n351));
  INV_X1    g150(.A(G190gat), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n349), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G183gat), .A2(G190gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT27), .B(G183gat), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT28), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n357), .A2(KEYINPUT67), .A3(new_n358), .A4(new_n352), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n347), .A2(new_n355), .A3(new_n356), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT23), .ZN(new_n361));
  INV_X1    g160(.A(new_n343), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT25), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT23), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n364), .B1(G169gat), .B2(G176gat), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n361), .A2(new_n362), .A3(new_n363), .A4(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n367), .B1(G183gat), .B2(G190gat), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OR2_X1    g169(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n361), .A2(new_n362), .A3(new_n365), .ZN(new_n372));
  AND2_X1   g171(.A1(G183gat), .A2(G190gat), .ZN(new_n373));
  OR2_X1    g172(.A1(KEYINPUT64), .A2(KEYINPUT24), .ZN(new_n374));
  NAND2_X1  g173(.A1(KEYINPUT64), .A2(KEYINPUT24), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n348), .A2(new_n352), .A3(KEYINPUT66), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT66), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n378), .B1(G183gat), .B2(G190gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n367), .B(KEYINPUT65), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n372), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n360), .B(new_n371), .C1(new_n383), .C2(new_n363), .ZN(new_n384));
  INV_X1    g183(.A(G226gat), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n385), .A2(new_n209), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n386), .A2(KEYINPUT29), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n366), .A2(new_n370), .ZN(new_n389));
  INV_X1    g188(.A(new_n372), .ZN(new_n390));
  AND2_X1   g189(.A1(KEYINPUT64), .A2(KEYINPUT24), .ZN(new_n391));
  NOR2_X1   g190(.A1(KEYINPUT64), .A2(KEYINPUT24), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n356), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n393), .A2(new_n379), .A3(new_n377), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT65), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n367), .B(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n390), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n389), .B1(new_n397), .B2(KEYINPUT25), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n388), .B1(new_n398), .B2(new_n360), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n262), .B1(new_n387), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n388), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n386), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n398), .A2(new_n360), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n402), .A2(new_n404), .A3(new_n277), .ZN(new_n405));
  XOR2_X1   g204(.A(G8gat), .B(G36gat), .Z(new_n406));
  XOR2_X1   g205(.A(G64gat), .B(G92gat), .Z(new_n407));
  XOR2_X1   g206(.A(new_n406), .B(new_n407), .Z(new_n408));
  XNOR2_X1  g207(.A(new_n408), .B(KEYINPUT75), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n400), .A2(new_n405), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT76), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n408), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n413), .B1(new_n400), .B2(new_n405), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT30), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n405), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT74), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n418), .B1(new_n268), .B2(new_n275), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n223), .A2(KEYINPUT74), .A3(new_n232), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n421), .B1(new_n402), .B2(new_n404), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n408), .B1(new_n417), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT77), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT30), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n414), .A2(KEYINPUT77), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT78), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT78), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n425), .A2(new_n427), .A3(new_n430), .A4(new_n426), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n416), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n384), .A2(new_n304), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n398), .A2(new_n309), .A3(new_n360), .ZN(new_n434));
  NAND2_X1  g233(.A1(G227gat), .A2(G233gat), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT34), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT34), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n433), .A2(new_n434), .A3(new_n438), .A4(new_n435), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G15gat), .B(G43gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(G71gat), .B(G99gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n435), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n384), .A2(new_n304), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n309), .B1(new_n398), .B2(new_n360), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  XOR2_X1   g246(.A(KEYINPUT69), .B(KEYINPUT33), .Z(new_n448));
  AOI21_X1  g247(.A(new_n443), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n440), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n448), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n433), .A2(new_n434), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n451), .B1(new_n452), .B2(new_n444), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n437), .B(new_n439), .C1(new_n453), .C2(new_n443), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n447), .A2(KEYINPUT32), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n456), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n450), .A2(new_n454), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n296), .A2(new_n337), .A3(new_n432), .A4(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT35), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n290), .A2(new_n291), .B1(new_n294), .B2(new_n207), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n464), .A2(new_n460), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n412), .A2(new_n415), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n400), .A2(new_n405), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT77), .B1(new_n467), .B2(new_n408), .ZN(new_n468));
  AOI211_X1 g267(.A(new_n424), .B(new_n413), .C1(new_n400), .C2(new_n405), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n430), .B1(new_n470), .B2(new_n426), .ZN(new_n471));
  INV_X1    g270(.A(new_n431), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n466), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n336), .A2(KEYINPUT87), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT87), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n322), .A2(new_n475), .A3(new_n327), .A4(new_n335), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n331), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT35), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT71), .B1(new_n457), .B2(new_n459), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT70), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n483), .B1(new_n457), .B2(new_n459), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT36), .ZN(new_n485));
  OAI22_X1  g284(.A1(KEYINPUT70), .A2(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT71), .ZN(new_n487));
  INV_X1    g286(.A(new_n459), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n458), .B1(new_n450), .B2(new_n454), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n490), .A2(new_n483), .A3(KEYINPUT36), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n432), .A2(new_n337), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n486), .A2(new_n491), .B1(new_n492), .B2(new_n464), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT40), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n318), .B1(new_n316), .B2(new_n317), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n320), .A2(new_n313), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n495), .A2(KEYINPUT39), .A3(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n326), .B1(new_n495), .B2(KEYINPUT39), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n494), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n328), .ZN(new_n500));
  NOR3_X1   g299(.A1(new_n497), .A2(new_n498), .A3(new_n494), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n473), .A2(new_n502), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n331), .A2(new_n474), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n387), .A2(new_n399), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n421), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n506), .B(KEYINPUT37), .C1(new_n277), .C2(new_n505), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n507), .A2(KEYINPUT86), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(KEYINPUT86), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT37), .B1(new_n400), .B2(new_n405), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT38), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n409), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n508), .A2(new_n509), .A3(new_n511), .A4(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT37), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n413), .B1(new_n467), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT38), .B1(new_n516), .B2(new_n510), .ZN(new_n517));
  AND2_X1   g316(.A1(new_n517), .A2(new_n470), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n504), .A2(new_n514), .A3(new_n518), .A4(new_n476), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n503), .A2(new_n296), .A3(new_n519), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n463), .A2(new_n481), .B1(new_n493), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G113gat), .B(G141gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n522), .B(new_n523), .ZN(new_n524));
  XOR2_X1   g323(.A(G169gat), .B(G197gat), .Z(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(KEYINPUT12), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT93), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(G8gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(G15gat), .B(G22gat), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n530), .B1(new_n531), .B2(G1gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n281), .A2(G15gat), .ZN(new_n533));
  INV_X1    g332(.A(G15gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(G22gat), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT16), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n533), .B(new_n535), .C1(new_n536), .C2(G1gat), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n532), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT92), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n531), .B(new_n540), .C1(new_n536), .C2(G1gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n537), .A2(KEYINPUT92), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n533), .A2(new_n535), .ZN(new_n543));
  INV_X1    g342(.A(G1gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n543), .A2(new_n529), .A3(new_n544), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n541), .A2(new_n542), .A3(new_n532), .A4(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n539), .B1(new_n546), .B2(G8gat), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(G29gat), .ZN(new_n549));
  INV_X1    g348(.A(G36gat), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n549), .A2(new_n550), .A3(KEYINPUT14), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT14), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n552), .B1(G29gat), .B2(G36gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(G29gat), .A2(G36gat), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n551), .A2(new_n553), .A3(KEYINPUT89), .A4(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT15), .ZN(new_n556));
  OR2_X1    g355(.A1(G43gat), .A2(G50gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(G43gat), .A2(G50gat), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n555), .A2(new_n559), .ZN(new_n561));
  AND3_X1   g360(.A1(new_n551), .A2(new_n553), .A3(new_n554), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n558), .A2(new_n556), .ZN(new_n563));
  XOR2_X1   g362(.A(KEYINPUT90), .B(G43gat), .Z(new_n564));
  AOI21_X1  g363(.A(new_n563), .B1(new_n564), .B2(new_n203), .ZN(new_n565));
  AOI22_X1  g364(.A1(new_n560), .A2(new_n561), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n548), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n555), .B(new_n559), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n562), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n547), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n567), .A2(KEYINPUT94), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(G229gat), .A2(G233gat), .ZN(new_n573));
  XOR2_X1   g372(.A(new_n573), .B(KEYINPUT13), .Z(new_n574));
  INV_X1    g373(.A(new_n571), .ZN(new_n575));
  OAI21_X1  g374(.A(KEYINPUT94), .B1(new_n547), .B2(new_n570), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n572), .A2(new_n574), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n570), .A2(KEYINPUT17), .ZN(new_n579));
  NOR3_X1   g378(.A1(new_n570), .A2(KEYINPUT91), .A3(KEYINPUT17), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT91), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT17), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n581), .B1(new_n566), .B2(new_n582), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n547), .B(new_n579), .C1(new_n580), .C2(new_n583), .ZN(new_n584));
  OAI211_X1 g383(.A(KEYINPUT18), .B(new_n573), .C1(new_n547), .C2(new_n570), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n578), .A2(new_n587), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n548), .A2(new_n566), .B1(G229gat), .B2(G233gat), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT18), .B1(new_n584), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n528), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n584), .A2(new_n589), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT18), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n594), .A2(new_n587), .A3(new_n578), .A4(new_n527), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT95), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n591), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n596), .B1(new_n591), .B2(new_n595), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n521), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G134gat), .B(G162gat), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT41), .ZN(new_n603));
  INV_X1    g402(.A(G232gat), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n603), .B1(new_n604), .B2(new_n209), .ZN(new_n605));
  XOR2_X1   g404(.A(new_n602), .B(new_n605), .Z(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(G99gat), .B(G106gat), .Z(new_n608));
  XNOR2_X1  g407(.A(KEYINPUT100), .B(KEYINPUT7), .ZN(new_n609));
  INV_X1    g408(.A(G85gat), .ZN(new_n610));
  INV_X1    g409(.A(G92gat), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G99gat), .A2(G106gat), .ZN(new_n613));
  AOI22_X1  g412(.A1(KEYINPUT8), .A2(new_n613), .B1(new_n610), .B2(new_n611), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NOR3_X1   g414(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n608), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OR3_X1    g416(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n618));
  INV_X1    g417(.A(new_n608), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n618), .A2(new_n619), .A3(new_n612), .A4(new_n614), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n579), .B(new_n621), .C1(new_n580), .C2(new_n583), .ZN(new_n622));
  XOR2_X1   g421(.A(G190gat), .B(G218gat), .Z(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NOR3_X1   g423(.A1(new_n603), .A2(new_n604), .A3(new_n209), .ZN(new_n625));
  INV_X1    g424(.A(new_n621), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n625), .B1(new_n626), .B2(new_n566), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n622), .A2(new_n624), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n624), .B1(new_n622), .B2(new_n627), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n607), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n630), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n632), .A2(new_n606), .A3(new_n628), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT97), .ZN(new_n636));
  OAI21_X1  g435(.A(KEYINPUT96), .B1(G71gat), .B2(G78gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(G57gat), .B(G64gat), .ZN(new_n638));
  AOI21_X1  g437(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AND2_X1   g439(.A1(G71gat), .A2(G78gat), .ZN(new_n641));
  NOR2_X1   g440(.A1(G71gat), .A2(G78gat), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  OR2_X1    g443(.A1(new_n641), .A2(new_n642), .ZN(new_n645));
  OR2_X1    g444(.A1(G57gat), .A2(G64gat), .ZN(new_n646));
  NAND2_X1  g445(.A1(G57gat), .A2(G64gat), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n646), .B(new_n647), .C1(new_n641), .C2(KEYINPUT9), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n645), .B1(new_n648), .B2(new_n637), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n636), .B1(new_n644), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n640), .A2(new_n643), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n648), .A2(new_n645), .A3(new_n637), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n651), .A2(new_n652), .A3(KEYINPUT97), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT21), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n547), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(KEYINPUT99), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT99), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n659), .B(new_n547), .C1(new_n655), .C2(new_n656), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n650), .A2(new_n656), .A3(new_n653), .ZN(new_n661));
  AND2_X1   g460(.A1(G231gat), .A2(G233gat), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(G127gat), .B(G155gat), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n664), .B(KEYINPUT20), .Z(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n661), .A2(new_n662), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n663), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n666), .B1(new_n663), .B2(new_n667), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n658), .B(new_n660), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n670), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n658), .A2(new_n660), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n672), .A2(new_n673), .A3(new_n668), .ZN(new_n674));
  XNOR2_X1  g473(.A(G183gat), .B(G211gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n675), .B(new_n676), .Z(new_n677));
  AND3_X1   g476(.A1(new_n671), .A2(new_n674), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n677), .B1(new_n671), .B2(new_n674), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n635), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(G120gat), .B(G148gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(G176gat), .B(G204gat), .ZN(new_n683));
  XOR2_X1   g482(.A(new_n682), .B(new_n683), .Z(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(G230gat), .A2(G233gat), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  XOR2_X1   g486(.A(KEYINPUT101), .B(KEYINPUT10), .Z(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n617), .A2(new_n620), .A3(new_n651), .A4(new_n652), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  AOI22_X1  g490(.A1(new_n650), .A2(new_n653), .B1(new_n617), .B2(new_n620), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n689), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  AND3_X1   g492(.A1(new_n617), .A2(new_n620), .A3(KEYINPUT10), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n654), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n687), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n691), .A2(new_n692), .A3(new_n686), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n685), .B1(new_n698), .B2(KEYINPUT102), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT102), .ZN(new_n700));
  OAI211_X1 g499(.A(new_n700), .B(new_n684), .C1(new_n696), .C2(new_n697), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n681), .A2(new_n703), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n601), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n337), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(G1gat), .ZN(G1324gat));
  NAND3_X1  g507(.A1(new_n601), .A2(new_n473), .A3(new_n704), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n709), .A2(G8gat), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT16), .B(G8gat), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT42), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n713), .B1(KEYINPUT42), .B2(new_n712), .ZN(G1325gat));
  NAND3_X1  g513(.A1(new_n705), .A2(new_n534), .A3(new_n461), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n482), .A2(KEYINPUT70), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n485), .B1(new_n460), .B2(KEYINPUT70), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n491), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n705), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n715), .B1(new_n720), .B2(new_n534), .ZN(G1326gat));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n464), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT43), .B(G22gat), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1327gat));
  NOR3_X1   g523(.A1(new_n492), .A2(new_n464), .A3(new_n460), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n481), .B1(new_n725), .B2(new_n478), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n492), .A2(new_n464), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n520), .A2(new_n718), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n591), .A2(new_n595), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(KEYINPUT95), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n597), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n678), .A2(new_n679), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n702), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(new_n634), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n729), .A2(new_n732), .A3(new_n736), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n737), .A2(G29gat), .A3(new_n337), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n738), .B(KEYINPUT45), .Z(new_n739));
  AOI21_X1  g538(.A(KEYINPUT44), .B1(new_n729), .B2(new_n635), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n741));
  AOI211_X1 g540(.A(new_n741), .B(new_n634), .C1(new_n726), .C2(new_n728), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n730), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n735), .A2(new_n744), .ZN(new_n745));
  AND3_X1   g544(.A1(new_n743), .A2(new_n706), .A3(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n739), .B1(new_n549), .B2(new_n746), .ZN(G1328gat));
  NOR3_X1   g546(.A1(new_n737), .A2(G36gat), .A3(new_n432), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT46), .ZN(new_n749));
  AND3_X1   g548(.A1(new_n743), .A2(new_n473), .A3(new_n745), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n550), .B2(new_n750), .ZN(G1329gat));
  NOR2_X1   g550(.A1(new_n718), .A2(new_n564), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n743), .A2(new_n745), .A3(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n564), .B1(new_n737), .B2(new_n460), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(KEYINPUT47), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT47), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n753), .A2(new_n757), .A3(new_n754), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(G1330gat));
  NOR2_X1   g558(.A1(new_n296), .A2(new_n203), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n743), .A2(new_n745), .A3(new_n760), .ZN(new_n761));
  XNOR2_X1  g560(.A(KEYINPUT104), .B(KEYINPUT48), .ZN(new_n762));
  OR2_X1    g561(.A1(new_n737), .A2(KEYINPUT103), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n296), .B1(new_n737), .B2(KEYINPUT103), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n761), .B(new_n762), .C1(new_n765), .C2(G50gat), .ZN(new_n766));
  INV_X1    g565(.A(new_n762), .ZN(new_n767));
  INV_X1    g566(.A(new_n761), .ZN(new_n768));
  AOI21_X1  g567(.A(G50gat), .B1(new_n763), .B2(new_n764), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n766), .A2(new_n770), .ZN(G1331gat));
  NOR3_X1   g570(.A1(new_n681), .A2(new_n730), .A3(new_n702), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n729), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(KEYINPUT105), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT105), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n729), .A2(new_n775), .A3(new_n772), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n777), .A2(new_n337), .ZN(new_n778));
  XNOR2_X1  g577(.A(KEYINPUT106), .B(G57gat), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n778), .B(new_n779), .ZN(G1332gat));
  NOR2_X1   g579(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT108), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n432), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n774), .A2(new_n776), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT107), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n785), .A2(KEYINPUT107), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n783), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OR2_X1    g588(.A1(new_n785), .A2(KEYINPUT107), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n790), .A2(new_n782), .A3(new_n786), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(new_n791), .ZN(G1333gat));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n793));
  INV_X1    g592(.A(G71gat), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n774), .A2(new_n776), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n794), .B1(new_n795), .B2(new_n719), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n777), .A2(G71gat), .A3(new_n460), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n793), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n795), .A2(new_n794), .A3(new_n461), .ZN(new_n799));
  OAI21_X1  g598(.A(G71gat), .B1(new_n777), .B2(new_n718), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n799), .A2(new_n800), .A3(KEYINPUT50), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n801), .ZN(G1334gat));
  NAND2_X1  g601(.A1(new_n795), .A2(new_n464), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g603(.A1(new_n733), .A2(new_n730), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n520), .A2(new_n718), .A3(new_n727), .ZN(new_n806));
  AOI22_X1  g605(.A1(new_n462), .A2(KEYINPUT35), .B1(new_n465), .B2(new_n480), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n635), .B(new_n805), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(KEYINPUT51), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n729), .A2(new_n810), .A3(new_n635), .A4(new_n805), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n812), .A2(new_n610), .A3(new_n706), .A4(new_n703), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n733), .A2(new_n730), .A3(new_n702), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n743), .A2(new_n706), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n813), .B1(new_n815), .B2(new_n610), .ZN(G1336gat));
  NOR3_X1   g615(.A1(new_n432), .A2(G92gat), .A3(new_n702), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n812), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n741), .B1(new_n521), .B2(new_n634), .ZN(new_n820));
  OAI211_X1 g619(.A(KEYINPUT44), .B(new_n635), .C1(new_n806), .C2(new_n807), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n820), .A2(new_n473), .A3(new_n821), .A4(new_n814), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(G92gat), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n818), .A2(new_n819), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n810), .A2(KEYINPUT109), .ZN(new_n825));
  XOR2_X1   g624(.A(new_n808), .B(new_n825), .Z(new_n826));
  AOI22_X1  g625(.A1(new_n826), .A2(new_n817), .B1(G92gat), .B2(new_n822), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n824), .B1(new_n827), .B2(new_n819), .ZN(G1337gat));
  NAND3_X1  g627(.A1(new_n743), .A2(new_n719), .A3(new_n814), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(G99gat), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n460), .A2(G99gat), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n812), .A2(new_n703), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(G1338gat));
  NOR3_X1   g632(.A1(new_n296), .A2(G106gat), .A3(new_n702), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n809), .A2(new_n811), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(KEYINPUT110), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT110), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n809), .A2(new_n837), .A3(new_n811), .A4(new_n834), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT53), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(G106gat), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n820), .A2(new_n464), .A3(new_n821), .A4(new_n814), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n841), .B2(KEYINPUT111), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT111), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n743), .A2(new_n843), .A3(new_n464), .A4(new_n814), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n839), .A2(new_n845), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n808), .A2(KEYINPUT109), .A3(new_n810), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n808), .B1(KEYINPUT109), .B2(new_n810), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n834), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n841), .A2(G106gat), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT53), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n846), .A2(new_n852), .ZN(G1339gat));
  NAND4_X1  g652(.A1(new_n733), .A2(new_n744), .A3(new_n634), .A4(new_n702), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT112), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n680), .A2(KEYINPUT112), .A3(new_n744), .A4(new_n702), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n574), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n575), .A2(new_n576), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n548), .A2(KEYINPUT94), .A3(new_n566), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n573), .B1(new_n584), .B2(new_n567), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n863), .B1(new_n864), .B2(KEYINPUT113), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT113), .ZN(new_n866));
  AOI211_X1 g665(.A(new_n866), .B(new_n573), .C1(new_n584), .C2(new_n567), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n526), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n595), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT54), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n684), .B1(new_n696), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n654), .A2(new_n621), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n688), .B1(new_n873), .B2(new_n690), .ZN(new_n874));
  INV_X1    g673(.A(new_n695), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n686), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n693), .A2(new_n695), .A3(new_n687), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(new_n877), .A3(KEYINPUT54), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n872), .A2(new_n878), .A3(KEYINPUT55), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n698), .A2(new_n684), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n872), .A2(new_n878), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT55), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n870), .A2(new_n635), .A3(new_n882), .A4(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n868), .A2(new_n595), .A3(new_n701), .A4(new_n699), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n888), .A2(KEYINPUT114), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n882), .A2(new_n730), .A3(new_n885), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(KEYINPUT114), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n887), .B1(new_n892), .B2(new_n634), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n859), .B1(new_n893), .B2(new_n733), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n894), .A2(new_n706), .A3(new_n432), .A4(new_n465), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT116), .ZN(new_n896));
  INV_X1    g695(.A(G113gat), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n896), .A2(new_n897), .A3(new_n730), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT115), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n706), .A2(new_n432), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n891), .A2(new_n890), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n635), .B1(new_n902), .B2(new_n889), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n734), .B1(new_n903), .B2(new_n887), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n901), .B1(new_n904), .B2(new_n859), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n905), .A2(KEYINPUT115), .A3(new_n465), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n900), .A2(new_n906), .A3(new_n732), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n898), .B1(new_n897), .B2(new_n907), .ZN(G1340gat));
  INV_X1    g707(.A(G120gat), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n896), .A2(new_n909), .A3(new_n703), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n900), .A2(new_n906), .A3(new_n703), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT117), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n911), .A2(new_n912), .A3(G120gat), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n912), .B1(new_n911), .B2(G120gat), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n910), .B1(new_n913), .B2(new_n914), .ZN(G1341gat));
  NAND3_X1  g714(.A1(new_n900), .A2(new_n906), .A3(new_n733), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(G127gat), .ZN(new_n917));
  OR2_X1    g716(.A1(new_n734), .A2(G127gat), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n895), .B2(new_n918), .ZN(G1342gat));
  INV_X1    g718(.A(KEYINPUT56), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n634), .A2(G134gat), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n905), .A2(new_n465), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT118), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n922), .A2(KEYINPUT118), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n920), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(new_n925), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(KEYINPUT56), .A3(new_n923), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n900), .A2(new_n906), .A3(new_n635), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(G134gat), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n926), .A2(new_n928), .A3(new_n930), .ZN(G1343gat));
  NOR2_X1   g730(.A1(new_n719), .A2(new_n901), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT119), .ZN(new_n933));
  AOI21_X1  g732(.A(KEYINPUT55), .B1(new_n883), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n872), .A2(new_n878), .A3(KEYINPUT119), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n881), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AOI22_X1  g735(.A1(new_n936), .A2(new_n732), .B1(new_n870), .B2(new_n703), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n886), .B1(new_n937), .B2(new_n635), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n858), .B1(new_n938), .B2(new_n734), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n464), .A2(KEYINPUT57), .ZN(new_n940));
  OAI21_X1  g739(.A(KEYINPUT120), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT120), .ZN(new_n942));
  INV_X1    g741(.A(new_n940), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n934), .A2(new_n935), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(new_n882), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n888), .B1(new_n945), .B2(new_n600), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(new_n634), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n733), .B1(new_n947), .B2(new_n886), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n942), .B(new_n943), .C1(new_n948), .C2(new_n858), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n941), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(KEYINPUT57), .B1(new_n894), .B2(new_n464), .ZN(new_n951));
  OAI211_X1 g750(.A(new_n732), .B(new_n932), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(G141gat), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n718), .A2(new_n464), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n905), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n600), .A2(G141gat), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT58), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n953), .A2(new_n958), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n730), .B(new_n932), .C1(new_n950), .C2(new_n951), .ZN(new_n960));
  AOI22_X1  g759(.A1(new_n960), .A2(G141gat), .B1(new_n956), .B2(new_n957), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT58), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(G1344gat));
  XOR2_X1   g762(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n964));
  AOI211_X1 g763(.A(G148gat), .B(new_n964), .C1(new_n956), .C2(new_n703), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n703), .B(new_n932), .C1(new_n950), .C2(new_n951), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT59), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n938), .A2(new_n734), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n704), .A2(new_n600), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g770(.A(KEYINPUT57), .B1(new_n971), .B2(new_n464), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n940), .B1(new_n904), .B2(new_n859), .ZN(new_n973));
  OR2_X1    g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n702), .A2(new_n964), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n975), .B1(new_n932), .B2(KEYINPUT122), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n976), .B1(KEYINPUT122), .B2(new_n932), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n968), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n965), .B1(new_n979), .B2(G148gat), .ZN(G1345gat));
  OAI21_X1  g779(.A(new_n932), .B1(new_n950), .B2(new_n951), .ZN(new_n981));
  OAI21_X1  g780(.A(G155gat), .B1(new_n981), .B2(new_n734), .ZN(new_n982));
  INV_X1    g781(.A(G155gat), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n956), .A2(new_n983), .A3(new_n733), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n982), .A2(new_n984), .ZN(G1346gat));
  INV_X1    g784(.A(G162gat), .ZN(new_n986));
  NOR3_X1   g785(.A1(new_n981), .A2(new_n986), .A3(new_n634), .ZN(new_n987));
  AOI21_X1  g786(.A(G162gat), .B1(new_n956), .B2(new_n635), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n987), .A2(new_n988), .ZN(G1347gat));
  NOR2_X1   g788(.A1(new_n706), .A2(new_n432), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(new_n461), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n296), .B1(new_n991), .B2(KEYINPUT123), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n992), .B1(KEYINPUT123), .B2(new_n991), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n993), .A2(new_n894), .ZN(new_n994));
  INV_X1    g793(.A(G169gat), .ZN(new_n995));
  NOR3_X1   g794(.A1(new_n994), .A2(new_n995), .A3(new_n600), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n706), .B1(new_n904), .B2(new_n859), .ZN(new_n997));
  NOR3_X1   g796(.A1(new_n464), .A2(new_n432), .A3(new_n460), .ZN(new_n998));
  AND2_X1   g797(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n999), .A2(new_n730), .ZN(new_n1000));
  AOI21_X1  g799(.A(new_n996), .B1(new_n1000), .B2(new_n995), .ZN(G1348gat));
  INV_X1    g800(.A(G176gat), .ZN(new_n1002));
  NOR3_X1   g801(.A1(new_n994), .A2(new_n1002), .A3(new_n702), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n997), .A2(new_n998), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n1002), .B1(new_n1004), .B2(new_n702), .ZN(new_n1005));
  OR2_X1    g804(.A1(new_n1005), .A2(KEYINPUT124), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1005), .A2(KEYINPUT124), .ZN(new_n1007));
  AOI21_X1  g806(.A(new_n1003), .B1(new_n1006), .B2(new_n1007), .ZN(G1349gat));
  NAND3_X1  g807(.A1(new_n999), .A2(new_n357), .A3(new_n733), .ZN(new_n1009));
  OAI21_X1  g808(.A(G183gat), .B1(new_n994), .B2(new_n734), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g810(.A(KEYINPUT125), .ZN(new_n1012));
  NAND3_X1  g811(.A1(new_n1011), .A2(new_n1012), .A3(KEYINPUT60), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n1012), .A2(KEYINPUT60), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n1009), .A2(new_n1014), .A3(new_n1010), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1013), .A2(new_n1015), .ZN(G1350gat));
  NAND3_X1  g815(.A1(new_n999), .A2(new_n352), .A3(new_n635), .ZN(new_n1017));
  OAI21_X1  g816(.A(G190gat), .B1(new_n994), .B2(new_n634), .ZN(new_n1018));
  AND2_X1   g817(.A1(new_n1018), .A2(KEYINPUT61), .ZN(new_n1019));
  NOR2_X1   g818(.A1(new_n1018), .A2(KEYINPUT61), .ZN(new_n1020));
  OAI21_X1  g819(.A(new_n1017), .B1(new_n1019), .B2(new_n1020), .ZN(G1351gat));
  AND3_X1   g820(.A1(new_n894), .A2(new_n337), .A3(new_n955), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n1022), .A2(new_n473), .ZN(new_n1023));
  INV_X1    g822(.A(new_n1023), .ZN(new_n1024));
  AOI21_X1  g823(.A(G197gat), .B1(new_n1024), .B2(new_n730), .ZN(new_n1025));
  AND2_X1   g824(.A1(new_n718), .A2(new_n990), .ZN(new_n1026));
  AND2_X1   g825(.A1(new_n974), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g826(.A1(new_n600), .A2(new_n269), .ZN(new_n1028));
  AOI21_X1  g827(.A(new_n1025), .B1(new_n1027), .B2(new_n1028), .ZN(G1352gat));
  NAND3_X1  g828(.A1(new_n974), .A2(new_n703), .A3(new_n1026), .ZN(new_n1030));
  NAND2_X1  g829(.A1(new_n1030), .A2(G204gat), .ZN(new_n1031));
  NAND4_X1  g830(.A1(new_n1022), .A2(new_n271), .A3(new_n473), .A4(new_n703), .ZN(new_n1032));
  NAND2_X1  g831(.A1(new_n1032), .A2(KEYINPUT62), .ZN(new_n1033));
  OR2_X1    g832(.A1(new_n1032), .A2(KEYINPUT62), .ZN(new_n1034));
  NAND3_X1  g833(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .ZN(G1353gat));
  OAI211_X1 g834(.A(new_n733), .B(new_n1026), .C1(new_n972), .C2(new_n973), .ZN(new_n1036));
  NAND2_X1  g835(.A1(new_n1036), .A2(G211gat), .ZN(new_n1037));
  INV_X1    g836(.A(KEYINPUT127), .ZN(new_n1038));
  INV_X1    g837(.A(KEYINPUT63), .ZN(new_n1039));
  NAND3_X1  g838(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g839(.A(KEYINPUT126), .ZN(new_n1041));
  NOR2_X1   g840(.A1(new_n734), .A2(new_n221), .ZN(new_n1042));
  INV_X1    g841(.A(new_n1042), .ZN(new_n1043));
  OAI21_X1  g842(.A(new_n1041), .B1(new_n1023), .B2(new_n1043), .ZN(new_n1044));
  NAND4_X1  g843(.A1(new_n1022), .A2(KEYINPUT126), .A3(new_n473), .A4(new_n1042), .ZN(new_n1045));
  NAND2_X1  g844(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g845(.A1(new_n1036), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1047));
  NAND2_X1  g846(.A1(new_n1047), .A2(KEYINPUT127), .ZN(new_n1048));
  AOI21_X1  g847(.A(KEYINPUT63), .B1(new_n1036), .B2(G211gat), .ZN(new_n1049));
  OAI211_X1 g848(.A(new_n1040), .B(new_n1046), .C1(new_n1048), .C2(new_n1049), .ZN(G1354gat));
  NAND3_X1  g849(.A1(new_n974), .A2(new_n635), .A3(new_n1026), .ZN(new_n1051));
  NAND2_X1  g850(.A1(new_n1051), .A2(G218gat), .ZN(new_n1052));
  NAND3_X1  g851(.A1(new_n1024), .A2(new_n211), .A3(new_n635), .ZN(new_n1053));
  NAND2_X1  g852(.A1(new_n1052), .A2(new_n1053), .ZN(G1355gat));
endmodule


