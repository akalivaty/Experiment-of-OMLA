//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 1 0 1 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 1 0 1 0 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 1 0 0 1 1 0 1 1 0 1 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000;
  INV_X1    g000(.A(G137), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT66), .B1(new_n187), .B2(G134), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT66), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G137), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(G137), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT11), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT65), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n188), .B(new_n191), .C1(new_n192), .C2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(KEYINPUT11), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n187), .A2(G134), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(KEYINPUT11), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n197), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(G131), .B1(new_n195), .B2(new_n200), .ZN(new_n201));
  AND2_X1   g015(.A1(new_n188), .A2(new_n191), .ZN(new_n202));
  OAI22_X1  g016(.A1(KEYINPUT65), .A2(new_n193), .B1(new_n190), .B2(G137), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(new_n194), .ZN(new_n204));
  INV_X1    g018(.A(G131), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n197), .A2(new_n198), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n202), .A2(new_n204), .A3(new_n205), .A4(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT67), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n201), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  OAI211_X1 g023(.A(KEYINPUT67), .B(G131), .C1(new_n195), .C2(new_n200), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT0), .B(G128), .ZN(new_n212));
  XNOR2_X1  g026(.A(G143), .B(G146), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G143), .ZN(new_n216));
  INV_X1    g030(.A(G143), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G146), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AND2_X1   g033(.A1(KEYINPUT0), .A2(G128), .ZN(new_n220));
  NOR2_X1   g034(.A1(KEYINPUT0), .A2(G128), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n219), .A2(new_n222), .A3(KEYINPUT64), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n213), .A2(new_n220), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n214), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n209), .A2(new_n210), .A3(new_n225), .ZN(new_n226));
  XOR2_X1   g040(.A(G116), .B(G119), .Z(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT2), .B(G113), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n227), .B(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT1), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n216), .A2(new_n218), .A3(new_n231), .A4(G128), .ZN(new_n232));
  INV_X1    g046(.A(G128), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n233), .B1(new_n216), .B2(KEYINPUT1), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n232), .B1(new_n234), .B2(new_n213), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT68), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n187), .A2(G134), .ZN(new_n237));
  OAI21_X1  g051(.A(G131), .B1(new_n192), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n232), .B(new_n239), .C1(new_n234), .C2(new_n213), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n236), .A2(new_n207), .A3(new_n238), .A4(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n226), .A2(new_n230), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT28), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n226), .A2(KEYINPUT69), .A3(new_n230), .A4(new_n241), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n226), .A2(new_n241), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n229), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n246), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n244), .B1(new_n250), .B2(KEYINPUT28), .ZN(new_n251));
  NOR2_X1   g065(.A1(G237), .A2(G953), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G210), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n253), .B(KEYINPUT27), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT26), .B(G101), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n254), .B(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT29), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(G902), .B1(new_n251), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n226), .A2(KEYINPUT30), .A3(new_n241), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n207), .A2(new_n238), .A3(new_n235), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT30), .B1(new_n226), .B2(new_n264), .ZN(new_n265));
  NOR3_X1   g079(.A1(new_n263), .A2(new_n265), .A3(new_n230), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n246), .A2(new_n247), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n257), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n258), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n226), .A2(new_n264), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n229), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n246), .A2(new_n247), .A3(new_n271), .ZN(new_n272));
  AOI211_X1 g086(.A(new_n257), .B(new_n244), .C1(new_n272), .C2(KEYINPUT28), .ZN(new_n273));
  OAI22_X1  g087(.A1(new_n260), .A2(new_n261), .B1(new_n269), .B2(new_n273), .ZN(new_n274));
  AOI211_X1 g088(.A(KEYINPUT71), .B(G902), .C1(new_n251), .C2(new_n259), .ZN(new_n275));
  OAI21_X1  g089(.A(G472), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT72), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n278), .B(G472), .C1(new_n274), .C2(new_n275), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT30), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n270), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(new_n229), .A3(new_n262), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n282), .A2(new_n246), .A3(new_n247), .A4(new_n256), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT31), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n267), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n286), .A2(KEYINPUT31), .A3(new_n256), .A4(new_n282), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n272), .A2(KEYINPUT28), .ZN(new_n288));
  INV_X1    g102(.A(new_n244), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI22_X1  g104(.A1(new_n285), .A2(new_n287), .B1(new_n290), .B2(new_n257), .ZN(new_n291));
  NOR2_X1   g105(.A1(G472), .A2(G902), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n292), .B(KEYINPUT70), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT32), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n285), .A2(new_n287), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n290), .A2(new_n257), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT32), .ZN(new_n298));
  INV_X1    g112(.A(new_n293), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n277), .A2(new_n279), .A3(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT9), .B(G234), .ZN(new_n303));
  OAI21_X1  g117(.A(G221), .B1(new_n303), .B2(G902), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G469), .ZN(new_n306));
  INV_X1    g120(.A(G902), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G104), .ZN(new_n309));
  OAI21_X1  g123(.A(KEYINPUT3), .B1(new_n309), .B2(G107), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT3), .ZN(new_n311));
  INV_X1    g125(.A(G107), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n312), .A3(G104), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n309), .A2(G107), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n310), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G101), .ZN(new_n316));
  INV_X1    g130(.A(G101), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n310), .A2(new_n313), .A3(new_n317), .A4(new_n314), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n316), .A2(KEYINPUT4), .A3(new_n318), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n216), .A2(new_n218), .A3(new_n220), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n219), .A2(new_n222), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n320), .B1(new_n321), .B2(new_n211), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT4), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n315), .A2(new_n323), .A3(G101), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n319), .A2(new_n223), .A3(new_n322), .A4(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n309), .A2(G107), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n312), .A2(G104), .ZN(new_n327));
  OAI21_X1  g141(.A(G101), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n318), .A2(new_n328), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n236), .A2(KEYINPUT10), .A3(new_n329), .A4(new_n240), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n209), .A2(new_n210), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT81), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT80), .B(KEYINPUT10), .ZN(new_n334));
  INV_X1    g148(.A(new_n232), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT1), .B1(new_n217), .B2(G146), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT79), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT79), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n216), .A2(new_n338), .A3(KEYINPUT1), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n337), .A2(G128), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n335), .B1(new_n340), .B2(new_n219), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n318), .A2(new_n328), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n334), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT81), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n209), .A2(new_n344), .A3(new_n210), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n331), .A2(new_n333), .A3(new_n343), .A4(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n343), .A2(new_n325), .A3(new_n330), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT84), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n343), .A2(new_n325), .A3(new_n330), .A4(KEYINPUT84), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n209), .A2(new_n210), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n346), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(G110), .B(G140), .ZN(new_n354));
  INV_X1    g168(.A(G953), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n355), .A2(G227), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n354), .B(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n336), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n219), .B1(new_n359), .B2(new_n233), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n342), .A2(new_n360), .A3(new_n232), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n361), .B1(new_n341), .B2(new_n342), .ZN(new_n362));
  XNOR2_X1  g176(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n362), .A2(new_n210), .A3(new_n209), .A4(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT83), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT83), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n351), .A2(new_n366), .A3(new_n362), .A4(new_n363), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT12), .ZN(new_n368));
  INV_X1    g182(.A(new_n362), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n368), .B1(new_n369), .B2(new_n332), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n365), .A2(new_n367), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n357), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n372), .A3(new_n346), .ZN(new_n373));
  AOI21_X1  g187(.A(G902), .B1(new_n358), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n308), .B1(new_n374), .B2(new_n306), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n347), .A2(new_n348), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(new_n351), .A3(new_n350), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(new_n372), .A3(new_n346), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n371), .A2(new_n346), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  OAI211_X1 g194(.A(G469), .B(new_n378), .C1(new_n380), .C2(new_n372), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n305), .B1(new_n375), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(G214), .B1(G237), .B2(G902), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n229), .A2(new_n319), .A3(new_n324), .ZN(new_n384));
  OR2_X1    g198(.A1(new_n227), .A2(new_n228), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT5), .ZN(new_n386));
  INV_X1    g200(.A(G119), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n387), .A3(G116), .ZN(new_n388));
  OAI211_X1 g202(.A(G113), .B(new_n388), .C1(new_n227), .C2(new_n386), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n329), .A2(new_n385), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n384), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(G110), .B(G122), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n384), .A2(new_n392), .A3(new_n390), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(KEYINPUT6), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT6), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n391), .A2(new_n397), .A3(new_n393), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n214), .A2(new_n223), .A3(G125), .A4(new_n224), .ZN(new_n399));
  INV_X1    g213(.A(G125), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n235), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n355), .A2(G224), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n402), .B(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n396), .A2(new_n398), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT85), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n396), .A2(KEYINPUT85), .A3(new_n398), .A4(new_n404), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n403), .A2(KEYINPUT7), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n402), .B(new_n409), .ZN(new_n410));
  XOR2_X1   g224(.A(new_n392), .B(KEYINPUT8), .Z(new_n411));
  NAND2_X1  g225(.A1(new_n389), .A2(new_n385), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n342), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n411), .B1(new_n413), .B2(new_n390), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(G902), .B1(new_n415), .B2(new_n395), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n407), .A2(new_n408), .A3(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(G210), .B1(G237), .B2(G902), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(KEYINPUT86), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n407), .A2(new_n418), .A3(new_n408), .A4(new_n416), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n382), .A2(new_n383), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G478), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n424), .A2(KEYINPUT15), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G116), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G122), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT89), .B(G122), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n428), .B1(new_n429), .B2(new_n427), .ZN(new_n430));
  OR2_X1    g244(.A1(new_n430), .A2(new_n312), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n233), .A2(G143), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT13), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n217), .A2(G128), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n217), .A2(KEYINPUT90), .A3(KEYINPUT13), .A4(G128), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT90), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT13), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n437), .B1(new_n434), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n435), .A2(new_n436), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(G134), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT91), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n434), .A2(new_n432), .A3(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n442), .B1(new_n434), .B2(new_n432), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n190), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n430), .A2(new_n312), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n431), .A2(new_n441), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT14), .B1(new_n429), .B2(new_n427), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n430), .A2(new_n449), .A3(G107), .ZN(new_n450));
  OAI221_X1 g264(.A(new_n428), .B1(KEYINPUT14), .B2(new_n312), .C1(new_n429), .C2(new_n427), .ZN(new_n451));
  INV_X1    g265(.A(new_n445), .ZN(new_n452));
  AOI21_X1  g266(.A(G134), .B1(new_n452), .B2(new_n443), .ZN(new_n453));
  NOR3_X1   g267(.A1(new_n444), .A2(new_n190), .A3(new_n445), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n450), .B(new_n451), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n448), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G217), .ZN(new_n457));
  NOR3_X1   g271(.A1(new_n303), .A2(new_n457), .A3(G953), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n456), .B(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n426), .B1(new_n460), .B2(new_n307), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n456), .A2(new_n459), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n458), .B1(new_n448), .B2(new_n455), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n307), .B(new_n426), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(G113), .B(G122), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(new_n309), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n252), .A2(G214), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n217), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n252), .A2(G143), .A3(G214), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(KEYINPUT18), .A3(G131), .ZN(new_n473));
  XNOR2_X1  g287(.A(G125), .B(G140), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(new_n215), .ZN(new_n475));
  NAND2_X1  g289(.A1(KEYINPUT18), .A2(G131), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n470), .A2(new_n471), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n473), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n472), .A2(G131), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n470), .A2(new_n205), .A3(new_n471), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n481), .A2(KEYINPUT17), .ZN(new_n482));
  INV_X1    g296(.A(G140), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(G125), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n400), .A2(G140), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n485), .A3(KEYINPUT16), .ZN(new_n486));
  OR3_X1    g300(.A1(new_n400), .A2(KEYINPUT16), .A3(G140), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n486), .A2(G146), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(G146), .B1(new_n486), .B2(new_n487), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT17), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n490), .B1(new_n491), .B2(new_n479), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n468), .B(new_n478), .C1(new_n482), .C2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n478), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n474), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT19), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n496), .B(KEYINPUT88), .C1(new_n497), .C2(new_n474), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n498), .B1(KEYINPUT88), .B2(new_n496), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n215), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n488), .B1(new_n479), .B2(new_n480), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n494), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n493), .B1(new_n502), .B2(new_n468), .ZN(new_n503));
  NOR2_X1   g317(.A1(G475), .A2(G902), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT20), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT20), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n503), .A2(new_n507), .A3(new_n504), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(G234), .A2(G237), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n510), .A2(G952), .A3(new_n355), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n510), .A2(G902), .A3(G953), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT21), .B(G898), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n478), .B1(new_n482), .B2(new_n492), .ZN(new_n516));
  INV_X1    g330(.A(new_n468), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(G902), .B1(new_n518), .B2(new_n493), .ZN(new_n519));
  INV_X1    g333(.A(G475), .ZN(new_n520));
  OR2_X1    g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n466), .A2(new_n509), .A3(new_n515), .A4(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n423), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n457), .B1(G234), .B2(new_n307), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n233), .A2(G119), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n387), .A2(G128), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT73), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT73), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n526), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(KEYINPUT24), .B(G110), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n529), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT74), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n526), .A2(new_n527), .A3(new_n535), .A4(KEYINPUT23), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(KEYINPUT23), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT23), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT74), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n537), .A2(new_n539), .A3(G119), .A4(new_n233), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n536), .A2(new_n540), .A3(G110), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n534), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n490), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT22), .B(G137), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(G221), .A2(G234), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT76), .B1(new_n547), .B2(G953), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT76), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n549), .A2(new_n355), .A3(G221), .A4(G234), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT77), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n551), .B1(new_n548), .B2(new_n550), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n546), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n554), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n556), .A2(new_n545), .A3(new_n552), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n533), .B1(new_n529), .B2(new_n531), .ZN(new_n559));
  AOI21_X1  g373(.A(G110), .B1(new_n536), .B2(new_n540), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT75), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n486), .A2(new_n487), .A3(G146), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n474), .A2(new_n215), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n561), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n526), .A2(new_n527), .A3(new_n530), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n530), .B1(new_n526), .B2(new_n527), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n532), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n536), .A2(new_n540), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n569), .B1(new_n570), .B2(G110), .ZN(new_n571));
  INV_X1    g385(.A(new_n565), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT75), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n544), .B(new_n558), .C1(new_n566), .C2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT78), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n558), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n555), .A2(new_n557), .A3(KEYINPUT78), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n562), .B1(new_n561), .B2(new_n565), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n571), .A2(KEYINPUT75), .A3(new_n572), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n543), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n574), .B(new_n307), .C1(new_n578), .C2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT25), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n544), .B1(new_n566), .B2(new_n573), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n576), .A2(new_n577), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n587), .A2(KEYINPUT25), .A3(new_n307), .A4(new_n574), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n525), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n587), .A2(new_n574), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n524), .A2(G902), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n589), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n302), .A2(new_n523), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(G101), .ZN(G3));
  INV_X1    g409(.A(new_n508), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n507), .B1(new_n503), .B2(new_n504), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n521), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n460), .A2(new_n307), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n424), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT33), .ZN(new_n601));
  OAI22_X1  g415(.A1(new_n462), .A2(new_n463), .B1(KEYINPUT93), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n424), .A2(G902), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT93), .B(KEYINPUT33), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n602), .B(new_n603), .C1(new_n460), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n598), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT94), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n598), .A2(KEYINPUT94), .A3(new_n606), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n383), .B1(new_n421), .B2(KEYINPUT92), .ZN(new_n612));
  INV_X1    g426(.A(new_n418), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n417), .A2(new_n613), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n421), .A2(KEYINPUT92), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n612), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n611), .A2(new_n616), .A3(new_n515), .ZN(new_n617));
  OAI21_X1  g431(.A(G472), .B1(new_n291), .B2(G902), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n297), .A2(new_n299), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n375), .A2(new_n381), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n304), .ZN(new_n623));
  INV_X1    g437(.A(new_n593), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n617), .A2(new_n621), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT95), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT34), .B(G104), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G6));
  INV_X1    g443(.A(new_n466), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n521), .A2(KEYINPUT96), .ZN(new_n631));
  OR3_X1    g445(.A1(new_n519), .A2(KEYINPUT96), .A3(new_n520), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n631), .A2(new_n509), .A3(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n616), .A2(new_n515), .A3(new_n630), .A4(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n635), .A2(new_n621), .A3(new_n625), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT98), .B(G107), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT97), .B(KEYINPUT35), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  INV_X1    g454(.A(KEYINPUT36), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n578), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT99), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n581), .A2(new_n643), .ZN(new_n644));
  AOI211_X1 g458(.A(KEYINPUT99), .B(new_n543), .C1(new_n579), .C2(new_n580), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n585), .A2(KEYINPUT99), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n581), .A2(new_n643), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n586), .A2(KEYINPUT36), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n592), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n589), .B1(KEYINPUT100), .B2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT100), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n651), .A2(new_n654), .A3(new_n592), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n522), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n656), .A2(new_n618), .A3(new_n619), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(new_n423), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT37), .B(G110), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G12));
  NAND3_X1  g474(.A1(new_n631), .A2(new_n509), .A3(new_n632), .ZN(new_n661));
  INV_X1    g475(.A(G900), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n512), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n511), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n661), .A2(new_n466), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n652), .A2(KEYINPUT100), .ZN(new_n668));
  INV_X1    g482(.A(new_n589), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n668), .A2(new_n669), .A3(new_n655), .ZN(new_n670));
  AND4_X1   g484(.A1(new_n382), .A2(new_n616), .A3(new_n667), .A4(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n302), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G128), .ZN(G30));
  NAND2_X1  g487(.A1(new_n286), .A2(new_n282), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n256), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n675), .B(new_n307), .C1(new_n250), .C2(new_n256), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(G472), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n301), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT101), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n665), .B(KEYINPUT39), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n382), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(new_n682), .B(KEYINPUT40), .Z(new_n683));
  AND2_X1   g497(.A1(new_n420), .A2(new_n421), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT38), .ZN(new_n685));
  INV_X1    g499(.A(new_n383), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n598), .A2(new_n630), .ZN(new_n687));
  NOR4_X1   g501(.A1(new_n685), .A2(new_n686), .A3(new_n670), .A4(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n680), .A2(new_n683), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G143), .ZN(G45));
  NOR2_X1   g504(.A1(new_n607), .A2(new_n666), .ZN(new_n691));
  AND4_X1   g505(.A1(new_n382), .A2(new_n616), .A3(new_n670), .A4(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n302), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G146), .ZN(G48));
  AND3_X1   g508(.A1(new_n371), .A2(new_n372), .A3(new_n346), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n372), .B1(new_n377), .B2(new_n346), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n307), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(G469), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n374), .A2(new_n306), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n698), .A2(new_n304), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(KEYINPUT102), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT102), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n698), .A2(new_n699), .A3(new_n702), .A4(new_n304), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n701), .A2(new_n593), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n302), .A2(new_n617), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT103), .ZN(new_n706));
  XOR2_X1   g520(.A(KEYINPUT41), .B(G113), .Z(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G15));
  NAND3_X1  g522(.A1(new_n701), .A2(new_n593), .A3(new_n703), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n634), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n710), .A2(KEYINPUT104), .A3(new_n302), .ZN(new_n711));
  AOI21_X1  g525(.A(KEYINPUT104), .B1(new_n710), .B2(new_n302), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(new_n427), .ZN(G18));
  AND4_X1   g528(.A1(new_n616), .A2(new_n701), .A3(new_n656), .A4(new_n703), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n302), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  NAND3_X1  g531(.A1(new_n701), .A2(new_n616), .A3(new_n703), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n295), .B1(new_n251), .B2(new_n256), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n299), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n687), .A2(new_n514), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n720), .A2(new_n721), .A3(new_n618), .A4(new_n593), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g537(.A(new_n723), .B(G122), .Z(G24));
  AND3_X1   g538(.A1(new_n701), .A2(new_n616), .A3(new_n703), .ZN(new_n725));
  AND4_X1   g539(.A1(new_n618), .A2(new_n691), .A3(new_n720), .A4(new_n670), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g541(.A(KEYINPUT105), .B(G125), .Z(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G27));
  NOR3_X1   g543(.A1(new_n422), .A2(new_n305), .A3(new_n686), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT106), .B1(new_n379), .B2(new_n357), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT106), .ZN(new_n732));
  AOI211_X1 g546(.A(new_n732), .B(new_n372), .C1(new_n371), .C2(new_n346), .ZN(new_n733));
  OAI211_X1 g547(.A(G469), .B(new_n378), .C1(new_n731), .C2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n375), .A2(new_n734), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n730), .A2(new_n593), .A3(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n302), .A2(new_n691), .A3(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT42), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n302), .A2(KEYINPUT42), .A3(new_n691), .A4(new_n736), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G131), .ZN(G33));
  NAND3_X1  g556(.A1(new_n302), .A2(new_n667), .A3(new_n736), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G134), .ZN(G36));
  OAI21_X1  g558(.A(new_n378), .B1(new_n380), .B2(new_n372), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT45), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n306), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI211_X1 g561(.A(KEYINPUT45), .B(new_n378), .C1(new_n731), .C2(new_n733), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n308), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(KEYINPUT107), .B1(new_n749), .B2(KEYINPUT46), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n750), .B1(new_n306), .B2(new_n374), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n749), .A2(KEYINPUT107), .A3(KEYINPUT46), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n751), .A2(KEYINPUT108), .A3(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n749), .A2(KEYINPUT46), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(KEYINPUT109), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(KEYINPUT108), .B1(new_n751), .B2(new_n752), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n304), .B(new_n681), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n600), .A2(new_n605), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n759), .A2(new_n598), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT43), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(KEYINPUT110), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT111), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n654), .B1(new_n651), .B2(new_n592), .ZN(new_n764));
  INV_X1    g578(.A(new_n592), .ZN(new_n765));
  AOI211_X1 g579(.A(KEYINPUT100), .B(new_n765), .C1(new_n646), .C2(new_n650), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n764), .A2(new_n766), .A3(new_n589), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n763), .B1(new_n621), .B2(new_n767), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n762), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n620), .A2(KEYINPUT111), .A3(new_n670), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT44), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n758), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n762), .A2(KEYINPUT44), .A3(new_n770), .A4(new_n768), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n773), .A2(KEYINPUT112), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n684), .A2(new_n383), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n775), .B1(new_n773), .B2(KEYINPUT112), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n774), .A2(KEYINPUT113), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT113), .B1(new_n774), .B2(new_n776), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n772), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G137), .ZN(G39));
  OAI21_X1  g594(.A(new_n304), .B1(new_n756), .B2(new_n757), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT47), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI211_X1 g597(.A(KEYINPUT47), .B(new_n304), .C1(new_n756), .C2(new_n757), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n302), .ZN(new_n786));
  NOR4_X1   g600(.A1(new_n775), .A2(new_n593), .A3(new_n607), .A4(new_n666), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G140), .ZN(G42));
  INV_X1    g603(.A(G952), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n761), .A2(new_n511), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n720), .A2(new_n618), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n792), .A2(new_n593), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  AOI211_X1 g609(.A(new_n790), .B(G953), .C1(new_n795), .C2(new_n725), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n701), .A2(new_n703), .ZN(new_n797));
  NOR4_X1   g611(.A1(new_n797), .A2(new_n624), .A3(new_n664), .A4(new_n775), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n679), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n611), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n786), .A2(new_n624), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n761), .A2(new_n511), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n803), .A2(new_n797), .A3(new_n775), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT117), .ZN(new_n806));
  NOR2_X1   g620(.A1(KEYINPUT118), .A2(KEYINPUT48), .ZN(new_n807));
  AND2_X1   g621(.A1(KEYINPUT118), .A2(KEYINPUT48), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  AOI211_X1 g623(.A(new_n801), .B(new_n809), .C1(new_n806), .C2(new_n807), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n799), .A2(new_n521), .A3(new_n509), .A4(new_n759), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n804), .A2(new_n670), .A3(new_n792), .ZN(new_n812));
  INV_X1    g626(.A(new_n685), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n797), .A2(new_n813), .A3(new_n383), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT50), .B1(new_n795), .B2(new_n814), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n795), .A2(KEYINPUT50), .A3(new_n814), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n811), .B(new_n812), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n698), .A2(new_n699), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n305), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n783), .A2(new_n784), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n794), .A2(new_n775), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n817), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n822), .A2(KEYINPUT51), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(KEYINPUT51), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n810), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n670), .A2(new_n633), .A3(new_n466), .A4(new_n665), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n826), .A2(new_n623), .A3(new_n775), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n302), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n726), .A2(new_n735), .A3(new_n730), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n743), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n830), .B1(new_n739), .B2(new_n740), .ZN(new_n831));
  AND4_X1   g645(.A1(new_n593), .A2(new_n721), .A3(new_n720), .A4(new_n618), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n656), .A2(new_n619), .A3(new_n618), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n422), .A2(new_n383), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n623), .A2(new_n834), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n725), .A2(new_n832), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n759), .A2(new_n598), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n837), .B1(new_n598), .B2(new_n630), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n838), .A2(new_n834), .A3(new_n514), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n839), .A2(new_n625), .A3(new_n621), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n836), .A2(new_n705), .A3(new_n716), .A4(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n594), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n302), .A2(new_n635), .A3(new_n704), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT104), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n831), .A2(new_n843), .A3(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n666), .A2(new_n305), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n735), .A2(new_n767), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n849), .B1(new_n301), .B2(new_n677), .ZN(new_n850));
  AOI211_X1 g664(.A(new_n687), .B(new_n612), .C1(new_n614), .C2(new_n615), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n302), .A2(new_n692), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n302), .A2(new_n671), .B1(new_n725), .B2(new_n726), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n852), .A2(KEYINPUT52), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT52), .B1(new_n852), .B2(new_n853), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT53), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT116), .B1(new_n847), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT53), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n850), .A2(new_n851), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n672), .A2(new_n693), .A3(new_n859), .A4(new_n727), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT52), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n852), .A2(KEYINPUT52), .A3(new_n853), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n858), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n839), .A2(new_n625), .A3(new_n621), .ZN(new_n865));
  OAI22_X1  g679(.A1(new_n718), .A2(new_n722), .B1(new_n657), .B2(new_n423), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n867), .A2(new_n594), .A3(new_n705), .A4(new_n716), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(new_n713), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT116), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n864), .A2(new_n869), .A3(new_n870), .A4(new_n831), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT115), .B1(new_n854), .B2(new_n855), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT115), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n862), .A2(new_n873), .A3(new_n863), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n872), .A2(new_n874), .A3(new_n869), .A4(new_n831), .ZN(new_n875));
  AOI22_X1  g689(.A1(new_n857), .A2(new_n871), .B1(new_n875), .B2(new_n858), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n875), .A2(KEYINPUT53), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT53), .B1(new_n862), .B2(new_n863), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n880), .A2(new_n869), .A3(new_n831), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n879), .A2(new_n881), .A3(KEYINPUT54), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  OAI22_X1  g697(.A1(new_n825), .A2(new_n883), .B1(G952), .B2(G953), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT49), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n818), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n818), .A2(new_n885), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n760), .A2(new_n593), .A3(new_n304), .A4(new_n383), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n679), .A2(new_n685), .A3(new_n889), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT114), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n884), .A2(new_n891), .ZN(G75));
  NOR2_X1   g706(.A1(new_n355), .A2(G952), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT120), .Z(new_n894));
  NOR2_X1   g708(.A1(new_n876), .A2(new_n307), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n895), .A2(new_n419), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n396), .A2(new_n398), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(new_n404), .ZN(new_n898));
  XOR2_X1   g712(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n899));
  XNOR2_X1  g713(.A(new_n898), .B(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT56), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n894), .B1(new_n896), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n895), .A2(G210), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n900), .B1(new_n904), .B2(new_n901), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n903), .A2(new_n905), .ZN(G51));
  NAND2_X1  g720(.A1(new_n857), .A2(new_n871), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n875), .A2(new_n858), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n909), .A2(KEYINPUT54), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n876), .A2(new_n877), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n308), .B(KEYINPUT57), .Z(new_n913));
  OAI22_X1  g727(.A1(new_n912), .A2(new_n913), .B1(new_n696), .B2(new_n695), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n895), .A2(new_n748), .A3(new_n747), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n893), .B1(new_n914), .B2(new_n915), .ZN(G54));
  INV_X1    g730(.A(KEYINPUT121), .ZN(new_n917));
  AND4_X1   g731(.A1(KEYINPUT58), .A2(new_n909), .A3(G475), .A4(G902), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n917), .B1(new_n918), .B2(new_n503), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n893), .B1(new_n918), .B2(new_n503), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n895), .A2(KEYINPUT58), .A3(G475), .ZN(new_n921));
  INV_X1    g735(.A(new_n503), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n921), .A2(KEYINPUT121), .A3(new_n922), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n919), .A2(new_n920), .A3(new_n923), .ZN(G60));
  OAI21_X1  g738(.A(new_n602), .B1(new_n460), .B2(new_n604), .ZN(new_n925));
  NAND2_X1  g739(.A1(G478), .A2(G902), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT59), .Z(new_n927));
  NOR2_X1   g741(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n928), .B1(new_n910), .B2(new_n911), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n929), .A2(KEYINPUT122), .A3(new_n894), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT122), .ZN(new_n931));
  INV_X1    g745(.A(new_n928), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n909), .A2(KEYINPUT54), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n932), .B1(new_n933), .B2(new_n878), .ZN(new_n934));
  INV_X1    g748(.A(new_n894), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n931), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n878), .A2(new_n882), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n925), .B1(new_n937), .B2(new_n927), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n930), .A2(new_n936), .A3(new_n938), .ZN(G63));
  NAND2_X1  g753(.A1(G217), .A2(G902), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT60), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n909), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n935), .B1(new_n943), .B2(new_n590), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT123), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n941), .B1(new_n907), .B2(new_n908), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n945), .B1(new_n946), .B2(new_n651), .ZN(new_n947));
  INV_X1    g761(.A(new_n651), .ZN(new_n948));
  NOR4_X1   g762(.A1(new_n876), .A2(KEYINPUT123), .A3(new_n948), .A4(new_n941), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n944), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT124), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n951), .B(new_n894), .C1(new_n946), .C2(new_n591), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n950), .A2(new_n954), .ZN(new_n955));
  OAI221_X1 g769(.A(new_n944), .B1(new_n951), .B2(KEYINPUT61), .C1(new_n947), .C2(new_n949), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(G66));
  NAND2_X1  g771(.A1(G224), .A2(G953), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n513), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n959), .B1(new_n869), .B2(new_n355), .ZN(new_n960));
  INV_X1    g774(.A(G898), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n897), .B1(new_n961), .B2(G953), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n960), .B(new_n962), .Z(G69));
  AND2_X1   g777(.A1(new_n853), .A2(new_n693), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n964), .A2(new_n741), .A3(new_n743), .ZN(new_n965));
  INV_X1    g779(.A(new_n758), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n802), .A2(new_n851), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n779), .A2(new_n788), .A3(new_n968), .A4(new_n355), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n263), .A2(new_n265), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(new_n499), .ZN(new_n971));
  NAND2_X1  g785(.A1(G900), .A2(G953), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n689), .A2(new_n964), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT62), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n689), .A2(KEYINPUT62), .A3(new_n964), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n682), .A2(new_n775), .A3(new_n838), .ZN(new_n979));
  AOI22_X1  g793(.A1(new_n977), .A2(new_n978), .B1(new_n802), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n779), .A2(new_n788), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n971), .B1(new_n981), .B2(new_n355), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n974), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n355), .B1(G227), .B2(G900), .ZN(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n983), .B(new_n985), .ZN(G72));
  NAND4_X1  g800(.A1(new_n779), .A2(new_n788), .A3(new_n869), .A4(new_n980), .ZN(new_n987));
  XOR2_X1   g801(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n988));
  NAND2_X1  g802(.A1(G472), .A2(G902), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n988), .B(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n675), .B1(new_n987), .B2(new_n990), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT126), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n674), .A2(new_n256), .ZN(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n994), .A2(new_n675), .A3(new_n990), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n995), .B(KEYINPUT127), .Z(new_n996));
  NAND3_X1  g810(.A1(new_n879), .A2(new_n881), .A3(new_n996), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n779), .A2(new_n788), .A3(new_n968), .A4(new_n869), .ZN(new_n998));
  AND2_X1   g812(.A1(new_n998), .A2(new_n990), .ZN(new_n999));
  OAI221_X1 g813(.A(new_n997), .B1(G952), .B2(new_n355), .C1(new_n999), .C2(new_n994), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n992), .A2(new_n1000), .ZN(G57));
endmodule


