//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 0 1 0 0 1 0 0 0 0 1 1 1 1 0 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1269, new_n1270, new_n1271, new_n1272, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  XOR2_X1   g0010(.A(KEYINPUT64), .B(G244), .Z(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G77), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G116), .A2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n216));
  NAND4_X1  g0016(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT65), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n210), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  OR2_X1    g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT66), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT67), .Z(new_n224));
  NOR2_X1   g0024(.A1(G58), .A2(G68), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G50), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR3_X1   g0028(.A1(new_n227), .A2(new_n208), .A3(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n210), .A2(G13), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n230), .B(G250), .C1(G257), .C2(G264), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT0), .Z(new_n232));
  NOR4_X1   g0032(.A1(new_n222), .A2(new_n224), .A3(new_n229), .A4(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  INV_X1    g0048(.A(G274), .ZN(new_n249));
  AND2_X1   g0049(.A1(G1), .A2(G13), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G41), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT68), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT68), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G41), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n252), .B(new_n207), .C1(new_n257), .C2(G45), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT69), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n250), .A2(new_n251), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n260), .A2(G226), .A3(new_n261), .ZN(new_n262));
  AND3_X1   g0062(.A1(new_n258), .A2(new_n259), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n259), .B1(new_n258), .B2(new_n262), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AND2_X1   g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  OAI21_X1  g0067(.A(KEYINPUT70), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT3), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT70), .ZN(new_n272));
  NAND2_X1  g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n268), .A2(new_n274), .A3(G222), .A4(new_n275), .ZN(new_n276));
  NAND4_X1  g0076(.A1(new_n268), .A2(new_n274), .A3(G223), .A4(G1698), .ZN(new_n277));
  NOR3_X1   g0077(.A1(new_n266), .A2(new_n267), .A3(KEYINPUT70), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n272), .B1(new_n271), .B2(new_n273), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G77), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n276), .B(new_n277), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n260), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n265), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G200), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n207), .A2(G20), .ZN(new_n288));
  NAND3_X1  g0088(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n288), .A2(new_n289), .A3(G50), .A4(new_n228), .ZN(new_n290));
  INV_X1    g0090(.A(G13), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(G1), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G20), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n290), .B1(G50), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n204), .A2(G20), .ZN(new_n295));
  INV_X1    g0095(.A(G150), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G20), .A2(G33), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n208), .A2(G33), .ZN(new_n299));
  XNOR2_X1  g0099(.A(KEYINPUT8), .B(G58), .ZN(new_n300));
  OAI221_X1 g0100(.A(new_n295), .B1(new_n296), .B2(new_n298), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n289), .A2(new_n228), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n294), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT9), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n303), .B(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n265), .A2(G190), .A3(new_n284), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NOR3_X1   g0107(.A1(new_n287), .A2(new_n307), .A3(KEYINPUT10), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT73), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n305), .A2(KEYINPUT73), .A3(new_n306), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n311), .A2(new_n312), .A3(new_n286), .ZN(new_n313));
  AND3_X1   g0113(.A1(new_n313), .A2(KEYINPUT74), .A3(KEYINPUT10), .ZN(new_n314));
  AOI21_X1  g0114(.A(KEYINPUT74), .B1(new_n313), .B2(KEYINPUT10), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n309), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n268), .A2(new_n274), .A3(G232), .A4(G1698), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n268), .A2(new_n274), .A3(G226), .A4(new_n275), .ZN(new_n318));
  INV_X1    g0118(.A(G97), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n317), .B(new_n318), .C1(new_n270), .C2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n283), .ZN(new_n321));
  INV_X1    g0121(.A(new_n258), .ZN(new_n322));
  AND2_X1   g0122(.A1(new_n260), .A2(new_n261), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n322), .B1(G238), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT13), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n321), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n325), .B1(new_n321), .B2(new_n324), .ZN(new_n328));
  OAI21_X1  g0128(.A(G200), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n328), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n330), .A2(G190), .A3(new_n326), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n297), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n281), .B2(new_n299), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n333), .A2(new_n302), .ZN(new_n334));
  OR2_X1    g0134(.A1(new_n334), .A2(KEYINPUT11), .ZN(new_n335));
  NOR3_X1   g0135(.A1(new_n291), .A2(new_n208), .A3(G1), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n203), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n337), .B(KEYINPUT12), .ZN(new_n338));
  INV_X1    g0138(.A(new_n302), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT72), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n339), .A2(new_n340), .A3(new_n293), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT72), .B1(new_n336), .B2(new_n302), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n341), .A2(new_n342), .A3(G68), .A4(new_n288), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n334), .A2(KEYINPUT11), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n335), .A2(new_n338), .A3(new_n343), .A4(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  AND3_X1   g0146(.A1(new_n329), .A2(new_n331), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n323), .A2(new_n212), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n258), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n280), .A2(G232), .A3(new_n275), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n280), .A2(G238), .A3(G1698), .ZN(new_n351));
  INV_X1    g0151(.A(G107), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n350), .B(new_n351), .C1(new_n352), .C2(new_n280), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n349), .B1(new_n353), .B2(new_n283), .ZN(new_n354));
  INV_X1    g0154(.A(G179), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n300), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n357), .A2(new_n297), .B1(G20), .B2(G77), .ZN(new_n358));
  OR2_X1    g0158(.A1(new_n358), .A2(KEYINPUT71), .ZN(new_n359));
  INV_X1    g0159(.A(new_n299), .ZN(new_n360));
  XOR2_X1   g0160(.A(KEYINPUT15), .B(G87), .Z(new_n361));
  AOI22_X1  g0161(.A1(new_n358), .A2(KEYINPUT71), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n339), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n341), .A2(new_n342), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n288), .A2(G77), .ZN(new_n365));
  OAI22_X1  g0165(.A1(new_n364), .A2(new_n365), .B1(G77), .B2(new_n293), .ZN(new_n366));
  OR2_X1    g0166(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n356), .B(new_n367), .C1(G169), .C2(new_n354), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n354), .A2(G190), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n363), .A2(new_n366), .ZN(new_n370));
  INV_X1    g0170(.A(G200), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n369), .B(new_n370), .C1(new_n371), .C2(new_n354), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(G169), .B1(new_n327), .B2(new_n328), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT14), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n330), .A2(G179), .A3(new_n326), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT14), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n377), .B(G169), .C1(new_n327), .C2(new_n328), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n375), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  AOI211_X1 g0179(.A(new_n347), .B(new_n373), .C1(new_n345), .C2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(G169), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n303), .B1(new_n285), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n265), .A2(new_n355), .A3(new_n284), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n293), .A2(new_n300), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n302), .B1(new_n207), .B2(G20), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n386), .B1(new_n387), .B2(new_n300), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  AND2_X1   g0189(.A1(G58), .A2(G68), .ZN(new_n390));
  OAI21_X1  g0190(.A(G20), .B1(new_n390), .B2(new_n225), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT75), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n297), .A2(G159), .ZN(new_n394));
  OAI211_X1 g0194(.A(KEYINPUT75), .B(G20), .C1(new_n390), .C2(new_n225), .ZN(new_n395));
  AND3_X1   g0195(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  NOR4_X1   g0197(.A1(new_n266), .A2(new_n267), .A3(new_n397), .A4(G20), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n208), .B1(new_n278), .B2(new_n279), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n398), .B1(new_n399), .B2(new_n397), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n396), .B1(new_n400), .B2(new_n203), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT16), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n266), .A2(new_n267), .ZN(new_n404));
  AOI21_X1  g0204(.A(KEYINPUT7), .B1(new_n404), .B2(new_n208), .ZN(new_n405));
  OAI21_X1  g0205(.A(G68), .B1(new_n405), .B2(new_n398), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n396), .A2(new_n406), .A3(KEYINPUT16), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n407), .A2(new_n302), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n389), .B1(new_n403), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n323), .A2(G232), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n258), .ZN(new_n411));
  XNOR2_X1  g0211(.A(KEYINPUT3), .B(G33), .ZN(new_n412));
  OR2_X1    g0212(.A1(G223), .A2(G1698), .ZN(new_n413));
  OR2_X1    g0213(.A1(new_n275), .A2(G226), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(G33), .A2(G87), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n260), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n411), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(G179), .ZN(new_n419));
  OAI21_X1  g0219(.A(G169), .B1(new_n411), .B2(new_n417), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT18), .B1(new_n409), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n424));
  INV_X1    g0224(.A(new_n398), .ZN(new_n425));
  AOI21_X1  g0225(.A(G20), .B1(new_n268), .B2(new_n274), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n425), .B1(new_n426), .B2(KEYINPUT7), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n424), .B1(new_n427), .B2(G68), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n302), .B(new_n407), .C1(new_n428), .C2(KEYINPUT16), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n388), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT18), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n430), .A2(new_n431), .A3(new_n421), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n423), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n415), .A2(new_n416), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n283), .ZN(new_n435));
  INV_X1    g0235(.A(G190), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n435), .A2(new_n436), .A3(new_n258), .A4(new_n410), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(new_n418), .B2(G200), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n427), .A2(G68), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT16), .B1(new_n439), .B2(new_n396), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n407), .A2(new_n302), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n438), .B(new_n388), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT76), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT76), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n429), .A2(new_n444), .A3(new_n388), .A4(new_n438), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n443), .A2(KEYINPUT17), .A3(new_n445), .ZN(new_n446));
  XNOR2_X1  g0246(.A(KEYINPUT77), .B(KEYINPUT17), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n409), .A2(new_n438), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n433), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  AND4_X1   g0249(.A1(new_n316), .A2(new_n380), .A3(new_n385), .A4(new_n449), .ZN(new_n450));
  AND2_X1   g0250(.A1(G264), .A2(G1698), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(new_n266), .B2(new_n267), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT83), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n412), .A2(KEYINPUT83), .A3(new_n451), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n412), .A2(G257), .A3(new_n275), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  XNOR2_X1  g0257(.A(KEYINPUT84), .B(G303), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n458), .B1(new_n268), .B2(new_n274), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n283), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT5), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n255), .A2(G41), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n253), .A2(KEYINPUT68), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n207), .B(G45), .C1(new_n461), .C2(G41), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n283), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(KEYINPUT5), .B1(new_n254), .B2(new_n256), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(new_n465), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n467), .A2(G270), .B1(new_n469), .B2(new_n252), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n460), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n207), .A2(G33), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n341), .A2(new_n342), .A3(G116), .A4(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(G116), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n292), .A2(G20), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G283), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n476), .B(new_n208), .C1(G33), .C2(new_n319), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n477), .B(new_n302), .C1(new_n208), .C2(G116), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT20), .ZN(new_n479));
  AND2_X1   g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n478), .A2(new_n479), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n473), .B(new_n475), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n471), .A2(G169), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT21), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT86), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT86), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n483), .A2(new_n487), .A3(new_n484), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  AOI211_X1 g0289(.A(new_n484), .B(new_n381), .C1(new_n460), .C2(new_n470), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n460), .A2(new_n470), .A3(G179), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n482), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT85), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI211_X1 g0295(.A(KEYINPUT85), .B(new_n482), .C1(new_n490), .C2(new_n492), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n482), .B1(new_n471), .B2(G200), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n460), .A2(new_n470), .A3(G190), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n489), .A2(new_n495), .A3(new_n496), .A4(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n476), .ZN(new_n501));
  OAI211_X1 g0301(.A(G244), .B(new_n275), .C1(new_n266), .C2(new_n267), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT4), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n268), .A2(new_n274), .A3(G250), .A4(G1698), .ZN(new_n505));
  AND2_X1   g0305(.A1(KEYINPUT4), .A2(G244), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n268), .A2(new_n274), .A3(new_n275), .A4(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n504), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n283), .ZN(new_n509));
  OAI211_X1 g0309(.A(G257), .B(new_n260), .C1(new_n468), .C2(new_n465), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n464), .A2(new_n252), .A3(new_n466), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT78), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT78), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n509), .A2(new_n514), .A3(new_n355), .A4(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT79), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n510), .A2(KEYINPUT78), .A3(new_n511), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT78), .B1(new_n510), .B2(new_n511), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n521), .A2(KEYINPUT79), .A3(new_n355), .A4(new_n509), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n352), .A2(KEYINPUT6), .A3(G97), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n319), .A2(new_n352), .ZN(new_n525));
  NOR2_X1   g0325(.A1(G97), .A2(G107), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n524), .B1(new_n527), .B2(KEYINPUT6), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n528), .A2(G20), .B1(G77), .B2(new_n297), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n400), .B2(new_n352), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n302), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n336), .A2(new_n319), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n339), .A2(new_n293), .A3(new_n472), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n532), .B1(new_n533), .B2(new_n319), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n512), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n509), .A2(new_n536), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n531), .A2(new_n535), .B1(new_n381), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n523), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g0339(.A(G244), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT80), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n270), .A2(new_n474), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n275), .A2(G238), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n543), .B1(new_n412), .B2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n412), .A2(KEYINPUT80), .A3(G244), .A4(G1698), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n542), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n283), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n207), .A2(new_n249), .A3(G45), .ZN(new_n549));
  INV_X1    g0349(.A(G250), .ZN(new_n550));
  INV_X1    g0350(.A(G45), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n550), .B1(new_n551), .B2(G1), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n260), .A2(new_n549), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(KEYINPUT81), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT81), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n548), .A2(new_n556), .A3(new_n553), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n555), .A2(new_n355), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n556), .B1(new_n548), .B2(new_n553), .ZN(new_n559));
  INV_X1    g0359(.A(new_n553), .ZN(new_n560));
  AOI211_X1 g0360(.A(KEYINPUT81), .B(new_n560), .C1(new_n547), .C2(new_n283), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n381), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n412), .A2(new_n208), .A3(G68), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n299), .A2(new_n319), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n563), .B1(KEYINPUT19), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n566), .A2(KEYINPUT82), .A3(new_n208), .ZN(new_n567));
  AOI21_X1  g0367(.A(KEYINPUT82), .B1(new_n566), .B2(new_n208), .ZN(new_n568));
  NOR3_X1   g0368(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n569));
  NOR3_X1   g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n302), .B1(new_n565), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n361), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n336), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n571), .B(new_n573), .C1(new_n572), .C2(new_n533), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n558), .A2(new_n562), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n555), .A2(G190), .A3(new_n557), .ZN(new_n576));
  OAI21_X1  g0376(.A(G200), .B1(new_n559), .B2(new_n561), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n571), .A2(new_n573), .ZN(new_n578));
  INV_X1    g0378(.A(G87), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n533), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n576), .A2(new_n577), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n534), .B1(new_n530), .B2(new_n302), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n509), .A2(new_n514), .A3(new_n515), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(G200), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n583), .B(new_n585), .C1(new_n436), .C2(new_n537), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n539), .A2(new_n575), .A3(new_n582), .A4(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n208), .B(G87), .C1(new_n266), .C2(new_n267), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT22), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n268), .A2(new_n274), .ZN(new_n590));
  OR3_X1    g0390(.A1(new_n579), .A2(KEYINPUT22), .A3(G20), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT23), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n593), .A2(new_n352), .A3(G20), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT87), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n593), .B2(new_n352), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n598));
  OAI22_X1  g0398(.A1(new_n594), .A2(new_n595), .B1(new_n598), .B2(G20), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n592), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT88), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT88), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n592), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n602), .A2(KEYINPUT24), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n603), .B1(new_n592), .B2(new_n600), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT24), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n339), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n336), .A2(new_n352), .ZN(new_n610));
  XOR2_X1   g0410(.A(KEYINPUT89), .B(KEYINPUT25), .Z(new_n611));
  XNOR2_X1  g0411(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n533), .A2(new_n352), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  OAI211_X1 g0415(.A(G257), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n275), .A2(G250), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n271), .B2(new_n273), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n616), .B1(new_n618), .B2(KEYINPUT90), .ZN(new_n619));
  NAND2_X1  g0419(.A1(G33), .A2(G294), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n550), .A2(G1698), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n266), .B2(new_n267), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT90), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n620), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n283), .B1(new_n619), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n467), .A2(G264), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(new_n511), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(KEYINPUT91), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n622), .A2(new_n623), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n412), .A2(KEYINPUT90), .A3(new_n621), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n629), .A2(new_n630), .A3(new_n620), .A4(new_n616), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n631), .A2(new_n283), .B1(G264), .B2(new_n467), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT91), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(new_n633), .A3(new_n511), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n628), .A2(new_n634), .A3(G169), .ZN(new_n635));
  INV_X1    g0435(.A(new_n627), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(G179), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n615), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n614), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n640), .B1(new_n605), .B2(new_n608), .ZN(new_n641));
  AOI21_X1  g0441(.A(G190), .B1(new_n628), .B2(new_n634), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n636), .A2(G200), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n639), .A2(new_n644), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n500), .A2(new_n587), .A3(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n450), .A2(new_n646), .ZN(G372));
  NAND2_X1  g0447(.A1(new_n379), .A2(new_n345), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n648), .B1(new_n347), .B2(new_n368), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n446), .A2(new_n448), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n433), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n313), .A2(KEYINPUT10), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT74), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n313), .A2(KEYINPUT74), .A3(KEYINPUT10), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n308), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n385), .B1(new_n651), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n316), .A2(new_n380), .A3(new_n385), .A4(new_n449), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT93), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n554), .A2(new_n381), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n558), .A2(new_n574), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n554), .A2(G200), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n576), .A2(new_n581), .A3(new_n663), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n662), .A2(new_n664), .A3(new_n523), .A4(new_n538), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n662), .B1(new_n665), .B2(KEYINPUT26), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT26), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n575), .A2(new_n582), .ZN(new_n668));
  INV_X1    g0468(.A(new_n539), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n660), .B1(new_n666), .B2(new_n670), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n662), .A2(new_n664), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n672), .A2(new_n667), .A3(new_n669), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n575), .A2(new_n582), .ZN(new_n674));
  OAI21_X1  g0474(.A(KEYINPUT26), .B1(new_n674), .B2(new_n539), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n673), .A2(new_n675), .A3(KEYINPUT93), .A4(new_n662), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n672), .A2(new_n644), .A3(new_n539), .A4(new_n586), .ZN(new_n677));
  INV_X1    g0477(.A(new_n482), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n471), .A2(KEYINPUT21), .A3(G169), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n678), .B1(new_n679), .B2(new_n491), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n680), .B1(new_n486), .B2(new_n488), .ZN(new_n681));
  AOI21_X1  g0481(.A(KEYINPUT92), .B1(new_n681), .B2(new_n639), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n681), .A2(KEYINPUT92), .A3(new_n639), .ZN(new_n684));
  AOI22_X1  g0484(.A1(new_n671), .A2(new_n676), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n658), .B1(new_n659), .B2(new_n685), .ZN(G369));
  AND3_X1   g0486(.A1(new_n483), .A2(new_n487), .A3(new_n484), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n487), .B1(new_n483), .B2(new_n484), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n496), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n680), .A2(KEYINPUT85), .ZN(new_n690));
  INV_X1    g0490(.A(new_n499), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT94), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n292), .A2(new_n208), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(new_n696), .A3(G213), .ZN(new_n697));
  INV_X1    g0497(.A(G343), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n678), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT94), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n701), .B1(new_n500), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n693), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n681), .A2(new_n701), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(G330), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n639), .B(new_n644), .C1(new_n641), .C2(new_n700), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT95), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n641), .B1(new_n635), .B2(new_n637), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n699), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n708), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n709), .B1(new_n708), .B2(new_n711), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n707), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n489), .A2(new_n495), .A3(new_n496), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n718), .B(new_n700), .C1(new_n713), .C2(new_n714), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n710), .A2(new_n700), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n717), .A2(new_n722), .ZN(G399));
  INV_X1    g0523(.A(new_n230), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n257), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n569), .A2(new_n474), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n726), .A2(G1), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(new_n227), .B2(new_n726), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT28), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT29), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(new_n685), .B2(new_n699), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n700), .A2(KEYINPUT29), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n668), .A2(new_n667), .A3(new_n669), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n665), .A2(KEYINPUT26), .ZN(new_n736));
  AND3_X1   g0536(.A1(new_n735), .A2(new_n662), .A3(new_n736), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n644), .A2(new_n539), .A3(new_n586), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n738), .B(new_n672), .C1(new_n718), .C2(new_n710), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n734), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n587), .ZN(new_n742));
  INV_X1    g0542(.A(new_n645), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n692), .A2(new_n742), .A3(new_n743), .A4(new_n700), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n632), .A2(new_n509), .A3(new_n536), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n491), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n559), .A2(new_n561), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n746), .A2(KEYINPUT30), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(G179), .B1(new_n548), .B2(new_n553), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n584), .A2(new_n471), .A3(new_n749), .A4(new_n627), .ZN(new_n750));
  AOI21_X1  g0550(.A(KEYINPUT30), .B1(new_n746), .B2(new_n747), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT96), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n748), .B(new_n750), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  AOI211_X1 g0553(.A(KEYINPUT96), .B(KEYINPUT30), .C1(new_n746), .C2(new_n747), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n699), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT31), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n748), .A2(new_n750), .ZN(new_n758));
  OAI211_X1 g0558(.A(KEYINPUT31), .B(new_n699), .C1(new_n758), .C2(new_n751), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n744), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n733), .A2(new_n741), .B1(G330), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n731), .B1(new_n761), .B2(G1), .ZN(G364));
  NOR2_X1   g0562(.A1(new_n291), .A2(G20), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n207), .B1(new_n763), .B2(G45), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n726), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n280), .A2(G355), .A3(new_n230), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n724), .A2(new_n412), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(G45), .B2(new_n227), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n244), .A2(new_n551), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n766), .B1(G116), .B2(new_n230), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT97), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G13), .A2(G33), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT98), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(new_n208), .ZN(new_n776));
  XOR2_X1   g0576(.A(new_n776), .B(KEYINPUT99), .Z(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n228), .B1(G20), .B2(new_n381), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n772), .A2(new_n773), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n208), .A2(G179), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G190), .A2(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n785), .A2(KEYINPUT100), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(KEYINPUT100), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  XNOR2_X1  g0589(.A(KEYINPUT101), .B(G159), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n792), .A2(KEYINPUT32), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(KEYINPUT32), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n436), .A2(G179), .A3(G200), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n208), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT102), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(G97), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n793), .A2(new_n794), .A3(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n208), .A2(new_n355), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G200), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n436), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(G190), .ZN(new_n803));
  AOI22_X1  g0603(.A1(G50), .A2(new_n802), .B1(new_n803), .B2(G68), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n800), .A2(G190), .A3(new_n371), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n800), .A2(new_n784), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n806), .A2(G58), .B1(new_n808), .B2(G77), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n783), .A2(G190), .A3(G200), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n783), .A2(new_n436), .A3(G200), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n811), .A2(G87), .B1(new_n813), .B2(G107), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n804), .A2(new_n280), .A3(new_n809), .A4(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G317), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(KEYINPUT33), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n816), .A2(KEYINPUT33), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n803), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n811), .A2(G303), .ZN(new_n820));
  INV_X1    g0620(.A(G294), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n819), .B(new_n820), .C1(new_n821), .C2(new_n796), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n789), .A2(G329), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n806), .A2(G322), .B1(new_n808), .B2(G311), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n802), .A2(G326), .B1(new_n813), .B2(G283), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n823), .A2(new_n590), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n799), .A2(new_n815), .B1(new_n822), .B2(new_n826), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n765), .B(new_n782), .C1(new_n779), .C2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n706), .B2(new_n777), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n707), .A2(new_n765), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n706), .A2(G330), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(G396));
  NAND2_X1  g0632(.A1(new_n367), .A2(new_n699), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n368), .A2(new_n372), .A3(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT104), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n368), .A2(new_n372), .A3(KEYINPUT104), .A4(new_n833), .ZN(new_n837));
  OR2_X1    g0637(.A1(new_n368), .A2(new_n700), .ZN(new_n838));
  AND3_X1   g0638(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n685), .B2(new_n699), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n671), .A2(new_n676), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n683), .A2(new_n684), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n699), .B1(new_n836), .B2(new_n837), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n760), .A2(G330), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT105), .ZN(new_n849));
  INV_X1    g0649(.A(new_n765), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(new_n846), .B2(new_n847), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  OR2_X1    g0652(.A1(new_n775), .A2(new_n779), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n850), .B1(G77), .B2(new_n853), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n796), .A2(new_n202), .B1(new_n812), .B2(new_n203), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n404), .B(new_n855), .C1(G50), .C2(new_n811), .ZN(new_n856));
  INV_X1    g0656(.A(G132), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n806), .A2(G143), .B1(new_n808), .B2(new_n791), .ZN(new_n858));
  INV_X1    g0658(.A(new_n803), .ZN(new_n859));
  INV_X1    g0659(.A(G137), .ZN(new_n860));
  INV_X1    g0660(.A(new_n802), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n858), .B1(new_n859), .B2(new_n296), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT34), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n856), .B1(new_n857), .B2(new_n788), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n862), .A2(new_n863), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n802), .A2(G303), .B1(new_n808), .B2(G116), .ZN(new_n866));
  INV_X1    g0666(.A(G283), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n866), .B1(new_n867), .B2(new_n859), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n868), .B(KEYINPUT103), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n789), .A2(G311), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n280), .B1(G294), .B2(new_n806), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n812), .A2(new_n579), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(G107), .B2(new_n811), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n870), .A2(new_n798), .A3(new_n871), .A4(new_n873), .ZN(new_n874));
  OAI22_X1  g0674(.A1(new_n864), .A2(new_n865), .B1(new_n869), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n854), .B1(new_n875), .B2(new_n779), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n877));
  INV_X1    g0677(.A(new_n775), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n852), .A2(new_n879), .ZN(G384));
  OR2_X1    g0680(.A1(new_n528), .A2(KEYINPUT35), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n528), .A2(KEYINPUT35), .ZN(new_n882));
  NOR3_X1   g0682(.A1(new_n228), .A2(new_n208), .A3(new_n474), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  XOR2_X1   g0684(.A(new_n884), .B(KEYINPUT36), .Z(new_n885));
  OR3_X1    g0685(.A1(new_n227), .A2(new_n281), .A3(new_n390), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n201), .A2(G68), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n207), .B(G13), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT38), .ZN(new_n890));
  INV_X1    g0690(.A(new_n697), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n396), .A2(new_n406), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT106), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT16), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n396), .A2(new_n406), .A3(KEYINPUT106), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n441), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n891), .B1(new_n896), .B2(new_n389), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n423), .A2(new_n432), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n897), .B1(new_n650), .B2(new_n898), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n443), .A2(new_n445), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n429), .A2(new_n388), .B1(new_n420), .B2(new_n419), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n697), .B1(new_n429), .B2(new_n388), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n901), .A2(new_n902), .A3(KEYINPUT37), .ZN(new_n903));
  OAI22_X1  g0703(.A1(new_n896), .A2(new_n389), .B1(new_n421), .B2(new_n891), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n904), .A2(new_n443), .A3(new_n445), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n900), .A2(new_n903), .B1(new_n905), .B2(KEYINPUT37), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n890), .B1(new_n899), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(KEYINPUT37), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n901), .A2(KEYINPUT37), .ZN(new_n909));
  INV_X1    g0709(.A(new_n902), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n909), .A2(new_n443), .A3(new_n445), .A4(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n912), .B(KEYINPUT38), .C1(new_n449), .C2(new_n897), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT107), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n907), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  OAI211_X1 g0715(.A(KEYINPUT107), .B(new_n890), .C1(new_n899), .C2(new_n906), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n915), .A2(KEYINPUT39), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n910), .B1(new_n650), .B2(new_n898), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n442), .B1(new_n409), .B2(new_n422), .ZN(new_n919));
  OAI21_X1  g0719(.A(KEYINPUT37), .B1(new_n919), .B2(new_n902), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n890), .B(new_n911), .C1(new_n918), .C2(new_n920), .ZN(new_n921));
  XOR2_X1   g0721(.A(KEYINPUT108), .B(KEYINPUT39), .Z(new_n922));
  NAND3_X1  g0722(.A1(new_n921), .A2(new_n913), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n917), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n379), .A2(new_n345), .A3(new_n700), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n915), .A2(new_n916), .ZN(new_n928));
  INV_X1    g0728(.A(new_n347), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n345), .A2(new_n699), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n648), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n345), .B(new_n699), .C1(new_n379), .C2(new_n347), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n368), .A2(new_n699), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n844), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n935), .B1(new_n685), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n928), .A2(new_n933), .A3(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n898), .A2(new_n891), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n927), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n659), .A2(new_n740), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n657), .B1(new_n733), .B2(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n941), .B(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n839), .B1(new_n931), .B2(new_n932), .ZN(new_n945));
  OAI211_X1 g0745(.A(KEYINPUT31), .B(new_n699), .C1(new_n753), .C2(new_n754), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n744), .A2(new_n757), .A3(new_n946), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n915), .A2(new_n945), .A3(new_n916), .A4(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT40), .ZN(new_n949));
  AND3_X1   g0749(.A1(new_n947), .A2(new_n877), .A3(new_n933), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n949), .B1(new_n921), .B2(new_n913), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n948), .A2(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n646), .A2(new_n700), .B1(new_n756), .B2(new_n755), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n659), .B1(new_n946), .B2(new_n953), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n952), .A2(new_n954), .ZN(new_n956));
  INV_X1    g0756(.A(G330), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n944), .A2(new_n958), .B1(new_n207), .B2(new_n763), .ZN(new_n959));
  AND2_X1   g0759(.A1(new_n944), .A2(new_n958), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n889), .B1(new_n959), .B2(new_n960), .ZN(G367));
  NAND2_X1  g0761(.A1(new_n718), .A2(new_n700), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n708), .A2(new_n711), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(KEYINPUT95), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n962), .B1(new_n964), .B2(new_n712), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n669), .A2(new_n699), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n539), .B(new_n586), .C1(new_n583), .C2(new_n700), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n969), .A2(KEYINPUT42), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n710), .A2(new_n586), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n699), .B1(new_n971), .B2(new_n539), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(new_n969), .B2(KEYINPUT42), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n581), .A2(new_n700), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT109), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n672), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n662), .B2(new_n976), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n970), .A2(new_n973), .B1(KEYINPUT43), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n716), .A2(new_n968), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n981), .B(new_n982), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n725), .B(KEYINPUT41), .Z(new_n984));
  AND3_X1   g0784(.A1(new_n964), .A2(new_n712), .A3(new_n962), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n707), .B1(new_n985), .B2(new_n965), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n985), .A2(new_n965), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n987), .A2(G330), .A3(new_n706), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n761), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(KEYINPUT110), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n719), .A2(new_n720), .A3(new_n968), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT45), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n992), .A2(new_n993), .ZN(new_n995));
  INV_X1    g0795(.A(new_n968), .ZN(new_n996));
  AOI21_X1  g0796(.A(KEYINPUT44), .B1(new_n721), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT44), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n998), .B(new_n968), .C1(new_n719), .C2(new_n720), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n994), .A2(new_n995), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n716), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT110), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n989), .A2(new_n1002), .A3(new_n761), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n997), .A2(new_n999), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n992), .B(new_n993), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1004), .A2(new_n717), .A3(new_n1005), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n991), .A2(new_n1001), .A3(new_n1003), .A4(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n984), .B1(new_n1007), .B2(new_n761), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n764), .B(KEYINPUT111), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n983), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n767), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n1012), .A2(new_n240), .B1(new_n230), .B2(new_n572), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n850), .B1(new_n781), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n280), .B1(new_n296), .B2(new_n805), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n812), .A2(new_n281), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(G143), .B2(new_n802), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n202), .B2(new_n810), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n1015), .B(new_n1018), .C1(G137), .C2(new_n789), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n803), .A2(new_n791), .B1(new_n808), .B2(G50), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1020), .A2(KEYINPUT113), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n797), .A2(G68), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1020), .A2(KEYINPUT113), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1019), .A2(new_n1021), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n796), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n1025), .A2(G107), .B1(new_n813), .B2(G97), .ZN(new_n1026));
  INV_X1    g0826(.A(G311), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1026), .B1(new_n821), .B2(new_n859), .C1(new_n1027), .C2(new_n861), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n810), .A2(new_n474), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(KEYINPUT46), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1028), .B1(KEYINPUT112), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n412), .B1(new_n808), .B2(G283), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n458), .B2(new_n805), .C1(KEYINPUT46), .C2(new_n1029), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(G317), .B2(new_n789), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1031), .B(new_n1034), .C1(KEYINPUT112), .C2(new_n1030), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1024), .A2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT114), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT47), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1014), .B1(new_n1038), .B2(new_n779), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n777), .B2(new_n978), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1011), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT115), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1041), .B(new_n1042), .ZN(G387));
  OR2_X1    g0843(.A1(new_n989), .A2(new_n761), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n726), .B1(new_n989), .B2(new_n761), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n715), .A2(new_n778), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n767), .B1(new_n237), .B2(new_n551), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n280), .A2(new_n230), .A3(new_n727), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  OR3_X1    g0850(.A1(new_n300), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1051));
  OAI21_X1  g0851(.A(KEYINPUT50), .B1(new_n300), .B2(G50), .ZN(new_n1052));
  AOI21_X1  g0852(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1051), .A2(new_n728), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n1050), .A2(new_n1054), .B1(new_n352), .B2(new_n724), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n850), .B1(new_n1055), .B2(new_n781), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n797), .A2(new_n361), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n201), .B2(new_n805), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT116), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n803), .A2(new_n357), .B1(new_n808), .B2(G68), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT117), .Z(new_n1061));
  AOI21_X1  g0861(.A(new_n404), .B1(new_n813), .B2(G97), .ZN(new_n1062));
  INV_X1    g0862(.A(G159), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1062), .B1(new_n281), .B2(new_n810), .C1(new_n861), .C2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G150), .B2(new_n789), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1059), .A2(new_n1061), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n789), .A2(G326), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n412), .B1(new_n813), .B2(G116), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n796), .A2(new_n867), .B1(new_n810), .B2(new_n821), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT118), .Z(new_n1070));
  INV_X1    g0870(.A(KEYINPUT48), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n458), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n806), .A2(G317), .B1(new_n808), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n802), .A2(G322), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1073), .B(new_n1074), .C1(new_n1027), .C2(new_n859), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1070), .B1(new_n1071), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n1071), .B2(new_n1075), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT49), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1067), .B(new_n1068), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1066), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1056), .B1(new_n1081), .B2(new_n779), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1047), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n986), .A2(new_n988), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1083), .B1(new_n1084), .B2(new_n1009), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1046), .A2(new_n1086), .ZN(G393));
  NAND2_X1  g0887(.A1(new_n1006), .A2(new_n1001), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n990), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1007), .A2(new_n1089), .A3(new_n725), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1088), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n996), .A2(new_n778), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G150), .A2(new_n802), .B1(new_n806), .B2(G159), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT51), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n789), .A2(G143), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n404), .B(new_n872), .C1(new_n357), .C2(new_n808), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n797), .A2(G77), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n803), .A2(G50), .B1(new_n811), .B2(G68), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n789), .A2(G322), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n280), .B1(G294), .B2(new_n808), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n811), .A2(G283), .B1(new_n813), .B2(G107), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(G116), .A2(new_n1025), .B1(new_n803), .B2(new_n1072), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(G317), .A2(new_n802), .B1(new_n806), .B2(G311), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT52), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n1094), .A2(new_n1099), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n1107), .A2(new_n779), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n767), .A2(new_n247), .B1(G97), .B2(new_n724), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n765), .B(new_n1108), .C1(new_n780), .C2(new_n1109), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1091), .A2(new_n1010), .B1(new_n1092), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1090), .A2(new_n1111), .ZN(G390));
  NAND3_X1  g0912(.A1(new_n917), .A2(new_n775), .A3(new_n923), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n850), .B1(new_n357), .B2(new_n853), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(KEYINPUT54), .B(G143), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n805), .A2(new_n857), .B1(new_n807), .B2(new_n1115), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n590), .B(new_n1116), .C1(new_n789), .C2(G125), .ZN(new_n1117));
  INV_X1    g0917(.A(G128), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n861), .A2(new_n1118), .B1(new_n812), .B2(new_n201), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(G137), .B2(new_n803), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n810), .A2(new_n296), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT53), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n797), .A2(G159), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1117), .A2(new_n1120), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n788), .A2(new_n821), .B1(new_n203), .B2(new_n812), .ZN(new_n1125));
  OR2_X1    g0925(.A1(new_n1125), .A2(KEYINPUT121), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(KEYINPUT121), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n590), .B1(new_n474), .B2(new_n805), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(G87), .B2(new_n811), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1126), .A2(new_n1097), .A3(new_n1127), .A4(new_n1129), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n802), .A2(G283), .B1(new_n808), .B2(G97), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n352), .B2(new_n859), .ZN(new_n1132));
  XOR2_X1   g0932(.A(new_n1132), .B(KEYINPUT120), .Z(new_n1133));
  OAI21_X1  g0933(.A(new_n1124), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1114), .B1(new_n1134), .B2(new_n779), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1113), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n926), .B1(new_n921), .B2(new_n913), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n737), .A2(new_n739), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n934), .B1(new_n1138), .B2(new_n844), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n933), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1137), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n926), .B1(new_n937), .B2(new_n933), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1141), .B1(new_n1142), .B2(new_n924), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n945), .A2(G330), .A3(new_n947), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n760), .A2(G330), .A3(new_n877), .A4(new_n933), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1141), .B(new_n1147), .C1(new_n1142), .C2(new_n924), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1136), .B1(new_n1149), .B2(new_n1009), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n760), .A2(G330), .A3(new_n877), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n1140), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n1144), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n1147), .A2(new_n1139), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n947), .A2(G330), .A3(new_n877), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n1140), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n937), .A2(new_n1155), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n957), .B1(new_n953), .B2(new_n946), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n450), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n943), .A2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(KEYINPUT119), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1163));
  AOI221_X4 g0963(.A(new_n657), .B1(new_n1160), .B2(new_n450), .C1(new_n733), .C2(new_n942), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1158), .A2(new_n1139), .A3(new_n1147), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n945), .A2(new_n1160), .B1(new_n1153), .B2(new_n1140), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n937), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1165), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT119), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1164), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1163), .A2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n725), .B1(new_n1152), .B2(new_n1171), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n1159), .A2(new_n1162), .A3(KEYINPUT119), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1169), .B1(new_n1164), .B2(new_n1168), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1175), .A2(new_n1149), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1151), .B1(new_n1172), .B2(new_n1176), .ZN(G378));
  OAI21_X1  g0977(.A(new_n1164), .B1(new_n1175), .B2(new_n1149), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n948), .A2(new_n949), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n957), .B1(new_n950), .B2(new_n951), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n303), .A2(new_n697), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n656), .A2(new_n384), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1184), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(new_n316), .B2(new_n385), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1183), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1184), .B1(new_n656), .B2(new_n384), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n316), .A2(new_n385), .A3(new_n1186), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1189), .A2(new_n1190), .A3(new_n1182), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1188), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1181), .A2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1140), .B1(new_n845), .B2(new_n935), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n939), .B1(new_n1195), .B2(new_n928), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1179), .A2(new_n1192), .A3(new_n1180), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1194), .A2(new_n927), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n1179), .A2(new_n1192), .A3(new_n1180), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1192), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n941), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1198), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(KEYINPUT57), .B1(new_n1178), .B2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1162), .B1(new_n1152), .B2(new_n1171), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1202), .A2(KEYINPUT57), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n725), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1203), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1193), .A2(new_n775), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n850), .B1(G50), .B2(new_n853), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n257), .A2(new_n412), .ZN(new_n1210));
  AOI211_X1 g1010(.A(G50), .B(new_n1210), .C1(new_n270), .C2(new_n253), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n812), .A2(new_n202), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n859), .A2(new_n319), .B1(new_n810), .B2(new_n281), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(G116), .C2(new_n802), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n789), .A2(G283), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1210), .B1(new_n352), .B2(new_n805), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n361), .B2(new_n808), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1214), .A2(new_n1022), .A3(new_n1215), .A4(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT58), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1211), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n797), .A2(G150), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n805), .A2(new_n1118), .B1(new_n807), .B2(new_n860), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(G132), .B2(new_n803), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1115), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n802), .A2(G125), .B1(new_n811), .B2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1221), .A2(new_n1223), .A3(new_n1225), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1226), .A2(KEYINPUT59), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(KEYINPUT59), .ZN(new_n1228));
  AOI211_X1 g1028(.A(G33), .B(G41), .C1(new_n813), .C2(new_n791), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(KEYINPUT122), .B(G124), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1228), .B(new_n1229), .C1(new_n788), .C2(new_n1230), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1220), .B1(new_n1219), .B2(new_n1218), .C1(new_n1227), .C2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1209), .B1(new_n1232), .B2(new_n779), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1202), .A2(new_n1010), .B1(new_n1208), .B2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1207), .A2(KEYINPUT123), .A3(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(KEYINPUT123), .B1(new_n1207), .B2(new_n1234), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1236), .A2(new_n1237), .ZN(G375));
  OAI21_X1  g1038(.A(new_n850), .B1(G68), .B2(new_n853), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1239), .B(KEYINPUT124), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n805), .A2(new_n867), .B1(new_n807), .B2(new_n352), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n280), .B(new_n1241), .C1(new_n789), .C2(G303), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1016), .B1(G294), .B2(new_n802), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n803), .A2(G116), .B1(new_n811), .B2(G97), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1242), .A2(new_n1057), .A3(new_n1243), .A4(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT125), .ZN(new_n1246));
  OR2_X1    g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n861), .A2(new_n857), .B1(new_n810), .B2(new_n1063), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1212), .B(new_n1248), .C1(new_n803), .C2(new_n1224), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n797), .A2(G50), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n789), .A2(G128), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n412), .B1(new_n805), .B2(new_n860), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(G150), .B2(new_n808), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .A4(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1247), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1240), .B1(new_n1256), .B2(new_n779), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1257), .B1(new_n933), .B2(new_n878), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(new_n1159), .B2(new_n1009), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1159), .A2(new_n1162), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1163), .A2(new_n1170), .A3(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1260), .B1(new_n1262), .B2(new_n984), .ZN(G381));
  AND2_X1   g1063(.A1(new_n852), .A2(new_n879), .ZN(new_n1264));
  AOI211_X1 g1064(.A(G396), .B(new_n1085), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  OR4_X1    g1066(.A1(G390), .A2(G378), .A3(G381), .A4(new_n1266), .ZN(new_n1267));
  OR3_X1    g1067(.A1(G375), .A2(G387), .A3(new_n1267), .ZN(G407));
  AOI21_X1  g1068(.A(new_n726), .B1(new_n1175), .B2(new_n1149), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1152), .A2(new_n1171), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1150), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1271), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1272));
  OAI211_X1 g1072(.A(G407), .B(G213), .C1(G343), .C2(new_n1272), .ZN(G409));
  INV_X1    g1073(.A(KEYINPUT126), .ZN(new_n1274));
  INV_X1    g1074(.A(G396), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1275), .B1(new_n1046), .B2(new_n1086), .ZN(new_n1276));
  OAI21_X1  g1076(.A(G390), .B1(new_n1265), .B2(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1042), .B1(new_n1276), .B2(new_n1265), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1278), .A2(new_n1090), .A3(new_n1111), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1277), .A2(new_n1279), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(new_n1280), .B(new_n1041), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT61), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n698), .A2(G213), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  OAI211_X1 g1084(.A(G378), .B(new_n1234), .C1(new_n1203), .C2(new_n1206), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1202), .ZN(new_n1286));
  NOR3_X1   g1086(.A1(new_n1204), .A2(new_n1286), .A3(new_n984), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1234), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1271), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1284), .B1(new_n1285), .B2(new_n1289), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1262), .A2(KEYINPUT60), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT60), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1292), .B1(new_n1164), .B2(new_n1168), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n725), .ZN(new_n1294));
  OAI211_X1 g1094(.A(G384), .B(new_n1260), .C1(new_n1291), .C2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1294), .B1(new_n1262), .B2(KEYINPUT60), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1264), .B1(new_n1296), .B2(new_n1259), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1284), .A2(G2897), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1295), .A2(new_n1297), .A3(new_n1299), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1282), .B1(new_n1290), .B2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT62), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1298), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1305), .B1(new_n1290), .B2(new_n1306), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1304), .A2(new_n1307), .ZN(new_n1308));
  AOI211_X1 g1108(.A(new_n1284), .B(new_n1298), .C1(new_n1285), .C2(new_n1289), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n1305), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1281), .B1(new_n1308), .B2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1290), .A2(KEYINPUT63), .A3(new_n1306), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1312), .B(new_n1282), .C1(new_n1290), .C2(new_n1303), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1281), .B1(KEYINPUT63), .B2(new_n1309), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1274), .B1(new_n1311), .B2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1304), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1290), .A2(new_n1306), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT63), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1317), .A2(new_n1320), .A3(new_n1281), .A4(new_n1312), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1318), .A2(KEYINPUT62), .ZN(new_n1322));
  NOR3_X1   g1122(.A1(new_n1322), .A2(new_n1304), .A3(new_n1307), .ZN(new_n1323));
  OAI211_X1 g1123(.A(KEYINPUT126), .B(new_n1321), .C1(new_n1323), .C2(new_n1281), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1316), .A2(new_n1324), .ZN(G405));
  NAND2_X1  g1125(.A1(new_n1207), .A2(new_n1234), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT123), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(G378), .B1(new_n1328), .B2(new_n1235), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1326), .A2(G378), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1330), .ZN(new_n1331));
  OAI211_X1 g1131(.A(KEYINPUT127), .B(new_n1306), .C1(new_n1329), .C2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1306), .A2(KEYINPUT127), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1272), .A2(new_n1333), .A3(new_n1330), .ZN(new_n1334));
  AND3_X1   g1134(.A1(new_n1332), .A2(new_n1281), .A3(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1281), .B1(new_n1332), .B2(new_n1334), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1335), .A2(new_n1336), .ZN(G402));
endmodule


