//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1 0 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT12), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G43gat), .B(G50gat), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NOR3_X1   g009(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G29gat), .ZN(new_n213));
  INV_X1    g012(.A(G36gat), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT87), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI211_X1 g014(.A(KEYINPUT15), .B(new_n208), .C1(new_n212), .C2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n208), .A2(KEYINPUT15), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT15), .ZN(new_n218));
  INV_X1    g017(.A(G43gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n219), .A2(G50gat), .ZN(new_n220));
  INV_X1    g019(.A(G50gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n221), .A2(G43gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n218), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  OR3_X1    g022(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(new_n209), .ZN(new_n225));
  INV_X1    g024(.A(new_n215), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n217), .A2(new_n223), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n216), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT17), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT88), .ZN(new_n231));
  INV_X1    g030(.A(G8gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(G15gat), .B(G22gat), .ZN(new_n233));
  INV_X1    g032(.A(G1gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT16), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n233), .A2(G1gat), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n231), .B(new_n232), .C1(new_n237), .C2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n238), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n231), .A2(new_n232), .ZN(new_n241));
  NAND2_X1  g040(.A1(KEYINPUT88), .A2(G8gat), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n240), .A2(new_n236), .A3(new_n241), .A4(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n216), .A2(new_n227), .A3(KEYINPUT17), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n230), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G229gat), .A2(G233gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n228), .A2(new_n239), .A3(new_n243), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT18), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT89), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n228), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n244), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(new_n248), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n247), .B(KEYINPUT13), .Z(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n249), .A2(KEYINPUT89), .A3(new_n250), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n253), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n246), .A2(KEYINPUT18), .A3(new_n247), .A4(new_n248), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(KEYINPUT90), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n207), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  XOR2_X1   g062(.A(new_n261), .B(KEYINPUT90), .Z(new_n264));
  NAND2_X1  g063(.A1(new_n206), .A2(new_n258), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT91), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n265), .B1(new_n266), .B2(new_n251), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n249), .A2(KEYINPUT91), .A3(new_n250), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n264), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n263), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT5), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT71), .ZN(new_n273));
  AND2_X1   g072(.A1(G113gat), .A2(G120gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(G113gat), .A2(G120gat), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(G113gat), .ZN(new_n277));
  INV_X1    g076(.A(G120gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G113gat), .A2(G120gat), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n279), .A2(KEYINPUT71), .A3(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G127gat), .B(G134gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT72), .B(KEYINPUT1), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n276), .A2(new_n281), .A3(new_n282), .A4(new_n283), .ZN(new_n284));
  XOR2_X1   g083(.A(G127gat), .B(G134gat), .Z(new_n285));
  NAND2_X1  g084(.A1(new_n279), .A2(new_n280), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n285), .B1(KEYINPUT1), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G155gat), .A2(G162gat), .ZN(new_n289));
  INV_X1    g088(.A(G155gat), .ZN(new_n290));
  INV_X1    g089(.A(G162gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G141gat), .B(G148gat), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n289), .B(new_n292), .C1(new_n293), .C2(KEYINPUT2), .ZN(new_n294));
  INV_X1    g093(.A(G141gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(G148gat), .ZN(new_n296));
  INV_X1    g095(.A(G148gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(G141gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n292), .A2(new_n289), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n289), .A2(KEYINPUT2), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n294), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n303), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n284), .A2(new_n287), .A3(new_n294), .A4(new_n302), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G225gat), .A2(G233gat), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n272), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n284), .A2(new_n287), .A3(KEYINPUT73), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT73), .B1(new_n284), .B2(new_n287), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT4), .ZN(new_n313));
  NOR4_X1   g112(.A1(new_n311), .A2(new_n312), .A3(new_n313), .A4(new_n303), .ZN(new_n314));
  AND3_X1   g113(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n300), .B1(new_n301), .B2(new_n299), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT3), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT3), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n294), .A2(new_n318), .A3(new_n302), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n317), .A2(new_n288), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n313), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(new_n321), .A3(new_n307), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n309), .B1(new_n314), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT73), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n288), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n303), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(new_n326), .A3(new_n310), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(new_n313), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n303), .A2(KEYINPUT3), .B1(new_n287), .B2(new_n284), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n308), .B1(new_n329), .B2(new_n319), .ZN(new_n330));
  OR2_X1    g129(.A1(new_n305), .A2(new_n313), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n328), .A2(new_n272), .A3(new_n330), .A4(new_n331), .ZN(new_n332));
  XOR2_X1   g131(.A(G1gat), .B(G29gat), .Z(new_n333));
  XNOR2_X1  g132(.A(new_n333), .B(KEYINPUT0), .ZN(new_n334));
  XNOR2_X1  g133(.A(G57gat), .B(G85gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n323), .A2(new_n332), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT6), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT80), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n336), .B1(new_n323), .B2(new_n332), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT80), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n337), .A2(new_n343), .A3(new_n338), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n340), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT81), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n323), .A2(new_n332), .ZN(new_n347));
  INV_X1    g146(.A(new_n336), .ZN(new_n348));
  AND4_X1   g147(.A1(new_n346), .A2(new_n347), .A3(KEYINPUT6), .A4(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n346), .B1(new_n341), .B2(KEYINPUT6), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n345), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G8gat), .B(G36gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n353), .B(KEYINPUT77), .ZN(new_n354));
  XNOR2_X1  g153(.A(G64gat), .B(G92gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n354), .B(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G197gat), .B(G204gat), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT22), .ZN(new_n358));
  INV_X1    g157(.A(G211gat), .ZN(new_n359));
  INV_X1    g158(.A(G218gat), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G211gat), .B(G218gat), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT75), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n363), .A2(new_n357), .A3(new_n361), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n362), .A2(KEYINPUT75), .A3(new_n364), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G226gat), .A2(G233gat), .ZN(new_n372));
  XOR2_X1   g171(.A(new_n372), .B(KEYINPUT76), .Z(new_n373));
  NAND2_X1  g172(.A1(G183gat), .A2(G190gat), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT70), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n376));
  NOR2_X1   g175(.A1(G169gat), .A2(G176gat), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT26), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NOR3_X1   g180(.A1(new_n376), .A2(new_n377), .A3(new_n375), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n374), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(G190gat), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT27), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n385), .A2(KEYINPUT69), .A3(G183gat), .ZN(new_n386));
  AND2_X1   g185(.A1(KEYINPUT69), .A2(G183gat), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n384), .B(new_n386), .C1(new_n387), .C2(new_n385), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT28), .ZN(new_n389));
  XNOR2_X1  g188(.A(KEYINPUT27), .B(G183gat), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n389), .A2(G190gat), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n388), .A2(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n383), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT25), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT66), .B1(new_n377), .B2(KEYINPUT23), .ZN(new_n395));
  NAND2_X1  g194(.A1(G169gat), .A2(G176gat), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT66), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT23), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n397), .B(new_n398), .C1(G169gat), .C2(G176gat), .ZN(new_n399));
  INV_X1    g198(.A(G169gat), .ZN(new_n400));
  INV_X1    g199(.A(G176gat), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n400), .A2(new_n401), .A3(KEYINPUT23), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n395), .A2(new_n396), .A3(new_n399), .A4(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT24), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n374), .A2(new_n404), .ZN(new_n405));
  OR2_X1    g204(.A1(G183gat), .A2(G190gat), .ZN(new_n406));
  NAND3_X1  g205(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n394), .B1(new_n403), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT67), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n399), .A2(new_n396), .A3(new_n402), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n400), .A2(new_n401), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n397), .B1(new_n412), .B2(new_n398), .ZN(new_n413));
  NOR3_X1   g212(.A1(new_n411), .A2(new_n413), .A3(new_n394), .ZN(new_n414));
  OR2_X1    g213(.A1(new_n405), .A2(KEYINPUT68), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n405), .A2(KEYINPUT68), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n415), .A2(new_n406), .A3(new_n407), .A4(new_n416), .ZN(new_n417));
  AOI22_X1  g216(.A1(new_n409), .A2(new_n410), .B1(new_n414), .B2(new_n417), .ZN(new_n418));
  OAI211_X1 g217(.A(KEYINPUT67), .B(new_n394), .C1(new_n403), .C2(new_n408), .ZN(new_n419));
  AOI211_X1 g218(.A(new_n373), .B(new_n393), .C1(new_n418), .C2(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n373), .A2(KEYINPUT29), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n409), .A2(new_n410), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n414), .A2(new_n417), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n422), .A2(new_n419), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n393), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n421), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n371), .B1(new_n420), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n373), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n424), .A2(new_n428), .A3(new_n425), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n393), .B1(new_n418), .B2(new_n419), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n429), .B(new_n370), .C1(new_n430), .C2(new_n421), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n356), .B1(new_n427), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n427), .A2(new_n356), .A3(new_n431), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT78), .ZN(new_n434));
  AOI22_X1  g233(.A1(KEYINPUT30), .A2(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n427), .A2(new_n431), .ZN(new_n436));
  INV_X1    g235(.A(new_n356), .ZN(new_n437));
  AND4_X1   g236(.A1(new_n434), .A2(new_n436), .A3(KEYINPUT30), .A4(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n432), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT79), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT30), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT79), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n432), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n352), .A2(new_n439), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n424), .A2(new_n425), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n311), .A2(new_n312), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n430), .A2(new_n448), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(G227gat), .A2(G233gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n453), .B(KEYINPUT64), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT34), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  XOR2_X1   g254(.A(new_n454), .B(KEYINPUT65), .Z(new_n456));
  NOR2_X1   g255(.A1(new_n456), .A2(KEYINPUT34), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n450), .A2(new_n451), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(G15gat), .B(G43gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(KEYINPUT74), .ZN(new_n461));
  INV_X1    g260(.A(G71gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n461), .B(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(G99gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n463), .B(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n456), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n466), .B1(new_n450), .B2(new_n451), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n465), .B1(new_n467), .B2(KEYINPUT33), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT32), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  AOI221_X4 g270(.A(new_n469), .B1(new_n465), .B2(KEYINPUT33), .C1(new_n452), .C2(new_n456), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n459), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n452), .A2(new_n456), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT32), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT33), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(new_n477), .A3(new_n465), .ZN(new_n478));
  INV_X1    g277(.A(new_n459), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n468), .A2(new_n470), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT83), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n365), .A2(new_n367), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT29), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n326), .B1(new_n485), .B2(new_n318), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n368), .A2(new_n369), .B1(new_n319), .B2(new_n484), .ZN(new_n487));
  INV_X1    g286(.A(G228gat), .ZN(new_n488));
  INV_X1    g287(.A(G233gat), .ZN(new_n489));
  OAI22_X1  g288(.A1(new_n486), .A2(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n487), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n488), .A2(new_n489), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n368), .A2(new_n484), .A3(new_n369), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n326), .B1(new_n494), .B2(new_n318), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n490), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(G22gat), .ZN(new_n497));
  INV_X1    g296(.A(G22gat), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n490), .B(new_n498), .C1(new_n493), .C2(new_n495), .ZN(new_n499));
  XNOR2_X1  g298(.A(KEYINPUT31), .B(G50gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(KEYINPUT82), .ZN(new_n501));
  XNOR2_X1  g300(.A(G78gat), .B(G106gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  AND4_X1   g302(.A1(new_n482), .A2(new_n497), .A3(new_n499), .A4(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n499), .A2(KEYINPUT83), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n505), .A2(new_n503), .B1(new_n497), .B2(new_n499), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n473), .A2(new_n481), .A3(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT35), .B1(new_n446), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT86), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g310(.A(KEYINPUT86), .B(KEYINPUT35), .C1(new_n446), .C2(new_n508), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n439), .A2(new_n445), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n473), .A2(new_n481), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n342), .A2(new_n338), .A3(new_n337), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n351), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n507), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n518), .A2(KEYINPUT35), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n515), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n511), .A2(new_n512), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n328), .A2(new_n320), .A3(new_n331), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(new_n308), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n304), .A2(new_n305), .A3(new_n307), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n523), .A2(KEYINPUT39), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT39), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n522), .A2(new_n526), .A3(new_n308), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(new_n336), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT40), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n341), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n525), .A2(KEYINPUT40), .A3(new_n336), .A4(new_n527), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n513), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT38), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n427), .A2(KEYINPUT37), .A3(new_n431), .ZN(new_n535));
  AOI21_X1  g334(.A(KEYINPUT85), .B1(new_n535), .B2(new_n356), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT37), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n536), .B1(new_n537), .B2(new_n436), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n535), .A2(KEYINPUT85), .A3(new_n356), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n534), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n441), .A2(new_n444), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT38), .B1(new_n436), .B2(new_n537), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n542), .A2(new_n356), .A3(new_n535), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n541), .A2(new_n543), .A3(new_n351), .A4(new_n516), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n533), .B(new_n507), .C1(new_n540), .C2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT36), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n514), .B(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n507), .A2(KEYINPUT84), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT84), .ZN(new_n549));
  NOR3_X1   g348(.A1(new_n504), .A2(new_n506), .A3(new_n549), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(new_n446), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n545), .A2(new_n547), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n271), .B1(new_n521), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G99gat), .B(G106gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(G99gat), .A2(G106gat), .ZN(new_n556));
  INV_X1    g355(.A(G85gat), .ZN(new_n557));
  INV_X1    g356(.A(G92gat), .ZN(new_n558));
  AOI22_X1  g357(.A1(KEYINPUT8), .A2(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT7), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT97), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT97), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT7), .ZN(new_n563));
  AND2_X1   g362(.A1(G85gat), .A2(G92gat), .ZN(new_n564));
  AND3_X1   g363(.A1(new_n561), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n564), .B1(new_n561), .B2(new_n563), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n555), .B(new_n559), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT98), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n561), .A2(new_n563), .ZN(new_n570));
  INV_X1    g369(.A(new_n564), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n561), .A2(new_n563), .A3(new_n564), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n574), .A2(KEYINPUT98), .A3(new_n555), .A4(new_n559), .ZN(new_n575));
  INV_X1    g374(.A(new_n555), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n559), .B1(new_n565), .B2(new_n566), .ZN(new_n577));
  AOI22_X1  g376(.A1(new_n569), .A2(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(new_n228), .ZN(new_n579));
  NAND3_X1  g378(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n230), .A2(new_n245), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n579), .B(new_n580), .C1(new_n581), .C2(new_n578), .ZN(new_n582));
  XNOR2_X1  g381(.A(G190gat), .B(G218gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(KEYINPUT99), .ZN(new_n585));
  XOR2_X1   g384(.A(G134gat), .B(G162gat), .Z(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT96), .ZN(new_n587));
  AOI21_X1  g386(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n582), .B(new_n583), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n590), .A2(new_n591), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G120gat), .B(G148gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(G176gat), .B(G204gat), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n595), .B(new_n596), .Z(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT100), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n577), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n574), .A2(KEYINPUT100), .A3(new_n559), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n600), .A2(new_n601), .A3(new_n576), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n569), .A2(new_n575), .ZN(new_n603));
  OAI21_X1  g402(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n604), .B1(G57gat), .B2(G64gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(G71gat), .B(G78gat), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT92), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(G57gat), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT9), .ZN(new_n611));
  NAND2_X1  g410(.A1(G71gat), .A2(G78gat), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n610), .A2(G64gat), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT93), .ZN(new_n614));
  INV_X1    g413(.A(G64gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n609), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n613), .A2(new_n614), .A3(new_n616), .A4(new_n606), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n606), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n612), .A2(new_n611), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n619), .B1(new_n609), .B2(new_n615), .ZN(new_n620));
  OAI21_X1  g419(.A(KEYINPUT93), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n607), .B1(new_n617), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n602), .A2(new_n603), .A3(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n623), .B1(new_n578), .B2(new_n622), .ZN(new_n624));
  NAND2_X1  g423(.A1(G230gat), .A2(G233gat), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(KEYINPUT101), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT101), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n624), .A2(new_n629), .A3(new_n626), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT10), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n623), .B(new_n632), .C1(new_n578), .C2(new_n622), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n578), .A2(KEYINPUT10), .A3(new_n622), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n626), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n598), .B1(new_n631), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n633), .A2(new_n634), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n625), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n638), .A2(new_n597), .A3(new_n628), .A4(new_n630), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT94), .B(KEYINPUT21), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n622), .A2(new_n641), .ZN(new_n642));
  AND2_X1   g441(.A1(G231gat), .A2(G233gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(G127gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  AOI22_X1  g445(.A1(new_n622), .A2(KEYINPUT21), .B1(new_n239), .B2(new_n243), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT95), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(G155gat), .ZN(new_n651));
  XOR2_X1   g450(.A(G183gat), .B(G211gat), .Z(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n648), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n648), .A2(new_n654), .ZN(new_n656));
  AOI211_X1 g455(.A(new_n594), .B(new_n640), .C1(new_n655), .C2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n352), .B(KEYINPUT102), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n554), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g459(.A1(new_n554), .A2(new_n657), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n232), .B1(new_n662), .B2(new_n513), .ZN(new_n663));
  INV_X1    g462(.A(new_n513), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT16), .B(G8gat), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n661), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT42), .B1(new_n663), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n667), .B1(KEYINPUT42), .B2(new_n666), .ZN(G1325gat));
  NOR3_X1   g467(.A1(new_n661), .A2(G15gat), .A3(new_n514), .ZN(new_n669));
  INV_X1    g468(.A(new_n547), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n662), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n669), .B1(G15gat), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT103), .ZN(G1326gat));
  INV_X1    g472(.A(new_n551), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n661), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT43), .B(G22gat), .Z(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1327gat));
  NAND2_X1  g476(.A1(new_n521), .A2(new_n553), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n594), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n594), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n682), .B1(new_n521), .B2(new_n553), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(KEYINPUT44), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n655), .A2(new_n656), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n640), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n689), .A2(new_n271), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n685), .A2(new_n658), .A3(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n213), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n693), .B1(new_n692), .B2(new_n691), .ZN(new_n694));
  AND4_X1   g493(.A1(new_n554), .A2(new_n594), .A3(new_n687), .A4(new_n688), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n695), .A2(new_n213), .A3(new_n658), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT45), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n694), .A2(new_n697), .ZN(G1328gat));
  NAND3_X1  g497(.A1(new_n695), .A2(new_n214), .A3(new_n513), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n699), .B(KEYINPUT46), .Z(new_n700));
  AND2_X1   g499(.A1(new_n685), .A2(new_n690), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n701), .A2(new_n513), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n700), .B1(new_n702), .B2(new_n214), .ZN(G1329gat));
  NAND3_X1  g502(.A1(new_n685), .A2(new_n670), .A3(new_n690), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(G43gat), .ZN(new_n705));
  INV_X1    g504(.A(new_n514), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n695), .A2(new_n219), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT47), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n705), .A2(KEYINPUT47), .A3(new_n707), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(G1330gat));
  AOI21_X1  g511(.A(new_n221), .B1(new_n701), .B2(new_n518), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n695), .A2(new_n221), .A3(new_n551), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT48), .ZN(new_n715));
  OR2_X1    g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n685), .A2(new_n551), .A3(new_n690), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n714), .B1(new_n717), .B2(G50gat), .ZN(new_n718));
  OAI22_X1  g517(.A1(new_n713), .A2(new_n716), .B1(new_n718), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g518(.A1(new_n686), .A2(new_n271), .A3(new_n682), .A4(new_n640), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n720), .B1(new_n521), .B2(new_n553), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n658), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT105), .B(G57gat), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1332gat));
  AOI21_X1  g523(.A(new_n664), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n726), .B(KEYINPUT106), .Z(new_n727));
  NOR2_X1   g526(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1333gat));
  AOI21_X1  g528(.A(new_n462), .B1(new_n721), .B2(new_n670), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n514), .A2(G71gat), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n730), .B1(new_n721), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g532(.A1(new_n721), .A2(new_n551), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g534(.A1(new_n686), .A2(new_n270), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n678), .A2(new_n594), .A3(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT51), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n683), .A2(KEYINPUT51), .A3(new_n736), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n741), .A2(new_n557), .A3(new_n640), .A4(new_n658), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n686), .A2(new_n270), .A3(new_n688), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n685), .A2(new_n743), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n744), .A2(new_n658), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n742), .B1(new_n745), .B2(new_n557), .ZN(G1336gat));
  NOR2_X1   g545(.A1(new_n664), .A2(G92gat), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n741), .A2(new_n640), .A3(new_n747), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n681), .A2(new_n513), .A3(new_n684), .A4(new_n743), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G92gat), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n748), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT108), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n748), .A2(new_n750), .A3(KEYINPUT108), .A4(new_n751), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT107), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n750), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n749), .A2(KEYINPUT107), .A3(G92gat), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n758), .A2(new_n759), .A3(new_n748), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT52), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n756), .A2(new_n761), .ZN(G1337gat));
  NAND4_X1  g561(.A1(new_n741), .A2(new_n464), .A3(new_n706), .A4(new_n640), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n744), .A2(new_n670), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n763), .B1(new_n764), .B2(new_n464), .ZN(G1338gat));
  NAND4_X1  g564(.A1(new_n681), .A2(new_n551), .A3(new_n684), .A4(new_n743), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(G106gat), .ZN(new_n767));
  INV_X1    g566(.A(new_n741), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n688), .A2(G106gat), .A3(new_n507), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(KEYINPUT109), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n767), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT53), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n681), .A2(new_n518), .A3(new_n684), .A4(new_n743), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT53), .B1(new_n773), .B2(G106gat), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n775), .B1(new_n741), .B2(new_n769), .ZN(new_n776));
  INV_X1    g575(.A(new_n769), .ZN(new_n777));
  AOI211_X1 g576(.A(KEYINPUT110), .B(new_n777), .C1(new_n739), .C2(new_n740), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n774), .B(KEYINPUT111), .C1(new_n776), .C2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  AND4_X1   g579(.A1(KEYINPUT51), .A2(new_n678), .A3(new_n594), .A4(new_n736), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT51), .B1(new_n683), .B2(new_n736), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n769), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(KEYINPUT110), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n741), .A2(new_n775), .A3(new_n769), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT111), .B1(new_n786), .B2(new_n774), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n772), .B1(new_n780), .B2(new_n787), .ZN(G1339gat));
  NAND3_X1  g587(.A1(new_n633), .A2(new_n626), .A3(new_n634), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n638), .A2(KEYINPUT54), .A3(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n597), .B1(new_n635), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n790), .A2(KEYINPUT55), .A3(new_n792), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n270), .A2(new_n795), .A3(new_n639), .A4(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n247), .B1(new_n246), .B2(new_n248), .ZN(new_n798));
  OAI22_X1  g597(.A1(new_n798), .A2(KEYINPUT112), .B1(new_n256), .B2(new_n257), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n798), .A2(KEYINPUT112), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n205), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT113), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n803), .B(new_n205), .C1(new_n799), .C2(new_n800), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n640), .A2(new_n805), .A3(new_n269), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n797), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT114), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n797), .A2(KEYINPUT114), .A3(new_n806), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n809), .A2(new_n682), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n639), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT55), .B1(new_n790), .B2(new_n792), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n805), .A2(new_n269), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n814), .A2(new_n815), .A3(new_n594), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n811), .A2(new_n816), .ZN(new_n817));
  AOI22_X1  g616(.A1(new_n817), .A2(new_n687), .B1(new_n271), .B2(new_n657), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n818), .A2(new_n551), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n819), .A2(new_n515), .A3(new_n658), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n820), .A2(new_n277), .A3(new_n271), .ZN(new_n821));
  INV_X1    g620(.A(new_n658), .ZN(new_n822));
  NOR4_X1   g621(.A1(new_n818), .A2(new_n513), .A3(new_n508), .A4(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(G113gat), .B1(new_n823), .B2(new_n270), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n821), .A2(new_n824), .ZN(G1340gat));
  NOR3_X1   g624(.A1(new_n820), .A2(new_n278), .A3(new_n688), .ZN(new_n826));
  AOI21_X1  g625(.A(G120gat), .B1(new_n823), .B2(new_n640), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n826), .A2(new_n827), .ZN(G1341gat));
  NOR3_X1   g627(.A1(new_n820), .A2(new_n645), .A3(new_n687), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n823), .A2(new_n686), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(KEYINPUT115), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n831), .A2(G127gat), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(KEYINPUT115), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n829), .B1(new_n832), .B2(new_n833), .ZN(G1342gat));
  INV_X1    g633(.A(G134gat), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n823), .A2(new_n835), .A3(new_n594), .ZN(new_n836));
  XOR2_X1   g635(.A(new_n836), .B(KEYINPUT56), .Z(new_n837));
  OAI21_X1  g636(.A(G134gat), .B1(new_n820), .B2(new_n682), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(G1343gat));
  INV_X1    g638(.A(KEYINPUT58), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n670), .A2(new_n822), .A3(new_n513), .ZN(new_n841));
  XNOR2_X1  g640(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n657), .A2(new_n271), .ZN(new_n844));
  INV_X1    g643(.A(new_n816), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n594), .B1(new_n807), .B2(new_n808), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n845), .B1(new_n846), .B2(new_n810), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n844), .B1(new_n847), .B2(new_n686), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n843), .B1(new_n848), .B2(new_n518), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n850));
  OAI21_X1  g649(.A(KEYINPUT117), .B1(new_n812), .B2(new_n813), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n795), .A2(new_n852), .A3(new_n639), .A4(new_n796), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n851), .A2(new_n270), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n594), .B1(new_n854), .B2(new_n806), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n687), .B1(new_n855), .B2(new_n845), .ZN(new_n856));
  AOI211_X1 g655(.A(new_n850), .B(new_n674), .C1(new_n856), .C2(new_n844), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n270), .B(new_n841), .C1(new_n849), .C2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(G141gat), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n670), .A2(new_n822), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n848), .A2(new_n518), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT119), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n513), .A2(new_n271), .A3(G141gat), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT119), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n848), .A2(new_n864), .A3(new_n518), .A4(new_n860), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n862), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT120), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n866), .A2(new_n867), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n840), .B(new_n859), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n871));
  INV_X1    g670(.A(new_n863), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n861), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n871), .B1(new_n875), .B2(KEYINPUT58), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n873), .B1(new_n858), .B2(G141gat), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n877), .A2(KEYINPUT118), .A3(new_n840), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n870), .B1(new_n876), .B2(new_n878), .ZN(G1344gat));
  OAI211_X1 g678(.A(new_n640), .B(new_n841), .C1(new_n849), .C2(new_n857), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n297), .A2(KEYINPUT59), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n880), .A2(KEYINPUT121), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT121), .B1(new_n880), .B2(new_n881), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n856), .A2(new_n844), .ZN(new_n884));
  OAI211_X1 g683(.A(KEYINPUT122), .B(new_n850), .C1(new_n884), .C2(new_n674), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n848), .A2(new_n518), .A3(new_n843), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n674), .B1(new_n856), .B2(new_n844), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n887), .B1(new_n888), .B2(KEYINPUT57), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n885), .A2(new_n886), .A3(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n841), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(new_n688), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n297), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894));
  OAI22_X1  g693(.A1(new_n882), .A2(new_n883), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n862), .A2(new_n664), .A3(new_n865), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n896), .A2(new_n297), .A3(new_n640), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(new_n897), .ZN(G1345gat));
  NAND3_X1  g697(.A1(new_n896), .A2(new_n290), .A3(new_n686), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n849), .A2(new_n857), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n900), .A2(new_n687), .A3(new_n891), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n899), .B1(new_n290), .B2(new_n901), .ZN(G1346gat));
  AOI21_X1  g701(.A(G162gat), .B1(new_n896), .B2(new_n594), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n900), .A2(new_n891), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n682), .A2(new_n291), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(G1347gat));
  NAND3_X1  g705(.A1(new_n822), .A2(new_n513), .A3(new_n706), .ZN(new_n907));
  XOR2_X1   g706(.A(new_n907), .B(KEYINPUT124), .Z(new_n908));
  NAND2_X1  g707(.A1(new_n819), .A2(new_n908), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n909), .A2(new_n400), .A3(new_n271), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n848), .A2(KEYINPUT123), .A3(new_n822), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT123), .B1(new_n848), .B2(new_n822), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n664), .A2(new_n508), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n270), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n910), .B1(new_n917), .B2(new_n400), .ZN(G1348gat));
  NAND3_X1  g717(.A1(new_n916), .A2(new_n401), .A3(new_n640), .ZN(new_n919));
  OAI21_X1  g718(.A(G176gat), .B1(new_n909), .B2(new_n688), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(G1349gat));
  INV_X1    g720(.A(KEYINPUT125), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n922), .A2(KEYINPUT60), .ZN(new_n923));
  OAI21_X1  g722(.A(G183gat), .B1(new_n909), .B2(new_n687), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n686), .A2(new_n390), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n915), .B(new_n925), .C1(new_n912), .C2(new_n913), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n923), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n922), .A2(KEYINPUT60), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n927), .B(new_n928), .ZN(G1350gat));
  NAND3_X1  g728(.A1(new_n916), .A2(new_n384), .A3(new_n594), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n819), .A2(new_n594), .A3(new_n908), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n932), .A2(KEYINPUT61), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n384), .B1(new_n932), .B2(KEYINPUT61), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n931), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n933), .B1(new_n931), .B2(new_n934), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n930), .B1(new_n935), .B2(new_n936), .ZN(G1351gat));
  NOR3_X1   g736(.A1(new_n670), .A2(new_n664), .A3(new_n658), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n890), .A2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(G197gat), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n939), .A2(new_n940), .A3(new_n271), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n547), .A2(new_n518), .A3(new_n513), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT127), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n914), .A2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(new_n270), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n941), .B1(new_n946), .B2(new_n940), .ZN(G1352gat));
  NOR2_X1   g746(.A1(new_n688), .A2(G204gat), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  OR3_X1    g748(.A1(new_n944), .A2(KEYINPUT62), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(G204gat), .B1(new_n939), .B2(new_n688), .ZN(new_n951));
  OAI21_X1  g750(.A(KEYINPUT62), .B1(new_n944), .B2(new_n949), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(G1353gat));
  NAND3_X1  g752(.A1(new_n890), .A2(new_n686), .A3(new_n938), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n954), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n955));
  AOI21_X1  g754(.A(KEYINPUT63), .B1(new_n954), .B2(G211gat), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n686), .A2(new_n359), .ZN(new_n957));
  OAI22_X1  g756(.A1(new_n955), .A2(new_n956), .B1(new_n944), .B2(new_n957), .ZN(G1354gat));
  OAI21_X1  g757(.A(G218gat), .B1(new_n939), .B2(new_n682), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n594), .A2(new_n360), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n959), .B1(new_n944), .B2(new_n960), .ZN(G1355gat));
endmodule


