//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 0 1 1 1 1 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1292, new_n1293;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XOR2_X1   g0007(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n208));
  XNOR2_X1  g0008(.A(new_n207), .B(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n209), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n205), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  OR2_X1    g0025(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT65), .ZN(new_n227));
  AOI211_X1 g0027(.A(new_n215), .B(new_n227), .C1(KEYINPUT1), .C2(new_n225), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XOR2_X1   g0037(.A(G107), .B(G116), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(G41), .ZN(new_n244));
  INV_X1    g0044(.A(G45), .ZN(new_n245));
  AOI21_X1  g0045(.A(G1), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(G33), .A2(G41), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n247), .A2(G1), .A3(G13), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n246), .A2(new_n248), .A3(G274), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(new_n248), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(new_n246), .ZN(new_n252));
  AND2_X1   g0052(.A1(new_n252), .A2(G226), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT3), .B(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n254), .A2(G222), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(G1698), .ZN(new_n257));
  INV_X1    g0057(.A(G223), .ZN(new_n258));
  OAI221_X1 g0058(.A(new_n256), .B1(new_n202), .B2(new_n254), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  AOI211_X1 g0059(.A(new_n250), .B(new_n253), .C1(new_n259), .C2(new_n251), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G190), .ZN(new_n261));
  XNOR2_X1  g0061(.A(new_n261), .B(KEYINPUT70), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G20), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G150), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT8), .B(G58), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n211), .A2(G33), .ZN(new_n266));
  OAI221_X1 g0066(.A(new_n264), .B1(new_n201), .B2(new_n211), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n210), .ZN(new_n269));
  INV_X1    g0069(.A(G50), .ZN(new_n270));
  INV_X1    g0070(.A(G1), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(G13), .A3(G20), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n267), .A2(new_n269), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n269), .ZN(new_n275));
  OR2_X1    g0075(.A1(new_n275), .A2(KEYINPUT66), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(KEYINPUT66), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n271), .A2(G20), .ZN(new_n278));
  XNOR2_X1  g0078(.A(new_n278), .B(KEYINPUT67), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n276), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n274), .B1(new_n280), .B2(new_n270), .ZN(new_n281));
  XOR2_X1   g0081(.A(new_n281), .B(KEYINPUT9), .Z(new_n282));
  NOR2_X1   g0082(.A1(new_n262), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT69), .ZN(new_n284));
  AOI21_X1  g0084(.A(KEYINPUT10), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G200), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n283), .B1(new_n286), .B2(new_n260), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  OAI221_X1 g0088(.A(new_n283), .B1(new_n284), .B2(KEYINPUT10), .C1(new_n286), .C2(new_n260), .ZN(new_n289));
  INV_X1    g0089(.A(G179), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n260), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n291), .B(new_n281), .C1(G169), .C2(new_n260), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n288), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT18), .ZN(new_n295));
  NAND2_X1  g0095(.A1(G58), .A2(G68), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n296), .B(KEYINPUT73), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n297), .B1(G58), .B2(G68), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n298), .A2(G20), .B1(G159), .B2(new_n263), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT7), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n300), .B1(new_n254), .B2(G20), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT3), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(G33), .ZN(new_n303));
  INV_X1    g0103(.A(G33), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n304), .A2(KEYINPUT3), .ZN(new_n305));
  OAI211_X1 g0105(.A(KEYINPUT7), .B(new_n211), .C1(new_n303), .C2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(KEYINPUT72), .B1(new_n307), .B2(G68), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT72), .ZN(new_n309));
  AOI211_X1 g0109(.A(new_n309), .B(new_n217), .C1(new_n301), .C2(new_n306), .ZN(new_n310));
  OAI211_X1 g0110(.A(KEYINPUT16), .B(new_n299), .C1(new_n308), .C2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT16), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT73), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n296), .B(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(G58), .A2(G68), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G159), .ZN(new_n317));
  INV_X1    g0117(.A(new_n263), .ZN(new_n318));
  OAI22_X1  g0118(.A1(new_n316), .A2(new_n211), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n217), .B1(new_n301), .B2(new_n306), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n312), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n311), .A2(new_n269), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n265), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n280), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(new_n273), .B2(new_n323), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n271), .B1(G41), .B2(G45), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n248), .A2(G232), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n249), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(G33), .A2(G87), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT74), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n330), .B(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n304), .A2(KEYINPUT3), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n302), .A2(G33), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n333), .A2(new_n334), .A3(G226), .A4(G1698), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n333), .A2(new_n334), .A3(G223), .A4(new_n255), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n332), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n329), .B1(new_n337), .B2(new_n251), .ZN(new_n338));
  INV_X1    g0138(.A(G169), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI211_X1 g0140(.A(new_n290), .B(new_n329), .C1(new_n251), .C2(new_n337), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n295), .B1(new_n326), .B2(new_n343), .ZN(new_n344));
  AOI211_X1 g0144(.A(KEYINPUT18), .B(new_n342), .C1(new_n322), .C2(new_n325), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT75), .ZN(new_n347));
  AOI211_X1 g0147(.A(G190), .B(new_n329), .C1(new_n251), .C2(new_n337), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n337), .A2(new_n251), .ZN(new_n349));
  INV_X1    g0149(.A(new_n329), .ZN(new_n350));
  AOI21_X1  g0150(.A(G200), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n347), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G190), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n349), .A2(new_n353), .A3(new_n350), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n354), .B(KEYINPUT75), .C1(G200), .C2(new_n338), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n322), .A2(new_n325), .A3(new_n352), .A4(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT17), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n352), .A2(new_n355), .ZN(new_n358));
  XOR2_X1   g0158(.A(KEYINPUT76), .B(KEYINPUT17), .Z(new_n359));
  NAND4_X1  g0159(.A1(new_n358), .A2(new_n322), .A3(new_n325), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n346), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n254), .A2(G232), .A3(G1698), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n254), .A2(G226), .A3(new_n255), .ZN(new_n365));
  NAND2_X1  g0165(.A1(G33), .A2(G97), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n251), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n250), .B1(G238), .B2(new_n252), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT13), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n370), .B1(new_n368), .B2(new_n369), .ZN(new_n373));
  OAI21_X1  g0173(.A(G169), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT14), .ZN(new_n375));
  INV_X1    g0175(.A(new_n373), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n371), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT14), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(new_n378), .A3(G169), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n375), .B(new_n379), .C1(new_n290), .C2(new_n377), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n279), .A2(G68), .A3(new_n275), .ZN(new_n381));
  XNOR2_X1  g0181(.A(new_n381), .B(KEYINPUT71), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n263), .A2(G50), .B1(G20), .B2(new_n217), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n202), .B2(new_n266), .ZN(new_n384));
  AND2_X1   g0184(.A1(new_n384), .A2(new_n269), .ZN(new_n385));
  OR2_X1    g0185(.A1(new_n385), .A2(KEYINPUT11), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n273), .A2(new_n217), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n387), .B(KEYINPUT12), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n385), .A2(KEYINPUT11), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n382), .A2(new_n386), .A3(new_n388), .A4(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n380), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n377), .A2(G200), .ZN(new_n392));
  INV_X1    g0192(.A(new_n390), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n376), .A2(G190), .A3(new_n371), .ZN(new_n394));
  AND3_X1   g0194(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n279), .A2(G77), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n397), .A2(new_n275), .B1(new_n202), .B2(new_n273), .ZN(new_n398));
  OAI22_X1  g0198(.A1(new_n265), .A2(new_n318), .B1(new_n211), .B2(new_n202), .ZN(new_n399));
  XNOR2_X1  g0199(.A(KEYINPUT15), .B(G87), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n400), .A2(new_n266), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n269), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n252), .A2(G244), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n254), .A2(G232), .A3(new_n255), .ZN(new_n405));
  OR2_X1    g0205(.A1(KEYINPUT68), .A2(G107), .ZN(new_n406));
  NAND2_X1  g0206(.A1(KEYINPUT68), .A2(G107), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI221_X1 g0208(.A(new_n405), .B1(new_n408), .B2(new_n254), .C1(new_n257), .C2(new_n218), .ZN(new_n409));
  AOI211_X1 g0209(.A(new_n250), .B(new_n404), .C1(new_n409), .C2(new_n251), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n403), .B1(new_n410), .B2(G190), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(new_n286), .B2(new_n410), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n410), .A2(new_n290), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n403), .B1(new_n410), .B2(G169), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  AND4_X1   g0216(.A1(new_n391), .A2(new_n396), .A3(new_n412), .A4(new_n416), .ZN(new_n417));
  AND3_X1   g0217(.A1(new_n294), .A2(new_n363), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(G13), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n420), .A2(G1), .ZN(new_n421));
  INV_X1    g0221(.A(G107), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(G20), .A3(new_n422), .ZN(new_n423));
  XNOR2_X1  g0223(.A(new_n423), .B(KEYINPUT25), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n271), .A2(G33), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n272), .A2(new_n425), .A3(new_n210), .A4(new_n268), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n424), .B1(G107), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT81), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n333), .A2(new_n334), .A3(new_n211), .A4(G87), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT22), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n254), .A2(KEYINPUT22), .A3(new_n211), .A4(G87), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT23), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n434), .A2(new_n422), .A3(G20), .ZN(new_n435));
  INV_X1    g0235(.A(G116), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n435), .B1(new_n436), .B2(new_n266), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n406), .A2(G20), .A3(new_n407), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT23), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n432), .A2(new_n433), .A3(new_n438), .A4(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT24), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n437), .B1(KEYINPUT23), .B2(new_n439), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT24), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n443), .A2(new_n444), .A3(new_n433), .A4(new_n432), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n429), .B1(new_n446), .B2(new_n269), .ZN(new_n447));
  INV_X1    g0247(.A(new_n269), .ZN(new_n448));
  AOI211_X1 g0248(.A(KEYINPUT81), .B(new_n448), .C1(new_n442), .C2(new_n445), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n428), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT77), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n244), .A2(KEYINPUT5), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n271), .A2(G45), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT5), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G41), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n456), .A2(KEYINPUT77), .A3(new_n271), .A4(G45), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n244), .A2(KEYINPUT5), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n454), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n459), .A2(G264), .A3(new_n248), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n333), .A2(new_n334), .A3(G257), .A4(G1698), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n333), .A2(new_n334), .A3(G250), .A4(new_n255), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G33), .A2(G294), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n251), .ZN(new_n465));
  INV_X1    g0265(.A(G274), .ZN(new_n466));
  INV_X1    g0266(.A(new_n210), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n466), .B1(new_n467), .B2(new_n247), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n454), .A2(new_n468), .A3(new_n457), .A4(new_n458), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n460), .A2(new_n465), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G169), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(new_n290), .B2(new_n470), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n450), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n470), .A2(new_n286), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(G190), .B2(new_n470), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n428), .B(new_n475), .C1(new_n447), .C2(new_n449), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT6), .ZN(new_n478));
  INV_X1    g0278(.A(G97), .ZN(new_n479));
  NOR3_X1   g0279(.A1(new_n478), .A2(new_n479), .A3(G107), .ZN(new_n480));
  XNOR2_X1  g0280(.A(G97), .B(G107), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n480), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  OAI22_X1  g0282(.A1(new_n482), .A2(new_n211), .B1(new_n202), .B2(new_n318), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n408), .B1(new_n301), .B2(new_n306), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n269), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n272), .A2(G97), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n486), .B1(new_n427), .B2(G97), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n333), .A2(new_n334), .A3(G244), .A4(new_n255), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(G250), .A2(G1698), .ZN(new_n492));
  NAND2_X1  g0292(.A1(KEYINPUT4), .A2(G244), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n492), .B1(new_n493), .B2(G1698), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n254), .A2(new_n494), .B1(G33), .B2(G283), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n251), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n459), .A2(G257), .A3(new_n248), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n497), .A2(new_n469), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n488), .B1(G200), .B2(new_n499), .ZN(new_n500));
  AND3_X1   g0300(.A1(new_n497), .A2(new_n469), .A3(new_n498), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G190), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n497), .A2(new_n290), .A3(new_n469), .A4(new_n498), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT78), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n248), .B1(new_n491), .B2(new_n495), .ZN(new_n505));
  INV_X1    g0305(.A(new_n469), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT78), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n507), .A2(new_n508), .A3(new_n290), .A4(new_n498), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n499), .A2(new_n339), .B1(new_n485), .B2(new_n487), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n500), .A2(new_n502), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G283), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n513), .B(new_n211), .C1(G33), .C2(new_n479), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n436), .A2(G20), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n514), .A2(new_n269), .A3(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT20), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n514), .A2(KEYINPUT20), .A3(new_n269), .A4(new_n515), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n272), .A2(new_n436), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(new_n427), .B2(new_n436), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n339), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n459), .A2(G270), .A3(new_n248), .ZN(new_n524));
  OAI21_X1  g0324(.A(G303), .B1(new_n303), .B2(new_n305), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n333), .A2(new_n334), .A3(G264), .A4(G1698), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n333), .A2(new_n334), .A3(G257), .A4(new_n255), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n251), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n524), .A2(new_n529), .A3(new_n469), .ZN(new_n530));
  AOI21_X1  g0330(.A(KEYINPUT21), .B1(new_n523), .B2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n530), .A2(G200), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n520), .A2(new_n522), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n524), .A2(new_n529), .A3(G190), .A4(new_n469), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n524), .A2(new_n529), .A3(G179), .A4(new_n469), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n534), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n523), .A2(new_n530), .A3(KEYINPUT21), .ZN(new_n541));
  AND4_X1   g0341(.A1(new_n532), .A2(new_n536), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n333), .A2(new_n334), .A3(new_n211), .A4(G68), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT79), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT79), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n254), .A2(new_n545), .A3(new_n211), .A4(G68), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT19), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n406), .A2(new_n219), .A3(new_n479), .A4(new_n407), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n366), .A2(new_n211), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR3_X1   g0350(.A1(new_n266), .A2(KEYINPUT19), .A3(new_n479), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n544), .B(new_n546), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n269), .ZN(new_n553));
  INV_X1    g0353(.A(new_n400), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n554), .A2(new_n272), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n427), .A2(new_n554), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n553), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n453), .A2(new_n220), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n271), .A2(new_n466), .A3(G45), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n559), .A2(new_n248), .A3(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n333), .A2(new_n334), .A3(G244), .A4(G1698), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n333), .A2(new_n334), .A3(G238), .A4(new_n255), .ZN(new_n563));
  NAND2_X1  g0363(.A1(G33), .A2(G116), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n561), .B1(new_n565), .B2(new_n251), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n290), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n558), .B(new_n567), .C1(G169), .C2(new_n566), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT80), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n426), .A2(new_n219), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n553), .A2(new_n556), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n565), .A2(new_n251), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n559), .A2(new_n248), .A3(new_n560), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G200), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n569), .B1(new_n572), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n566), .A2(G190), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n555), .B1(new_n552), .B2(new_n269), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n580), .A2(KEYINPUT80), .A3(new_n576), .A4(new_n571), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n512), .A2(new_n542), .A3(new_n568), .A4(new_n582), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n419), .A2(new_n477), .A3(new_n583), .ZN(G372));
  INV_X1    g0384(.A(new_n292), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n288), .A2(new_n289), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n396), .A2(new_n415), .B1(new_n390), .B2(new_n380), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n357), .A2(new_n360), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n346), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n585), .B1(new_n586), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n581), .A2(new_n579), .ZN(new_n591));
  AOI211_X1 g0391(.A(new_n555), .B(new_n570), .C1(new_n552), .C2(new_n269), .ZN(new_n592));
  AOI21_X1  g0392(.A(KEYINPUT80), .B1(new_n592), .B2(new_n576), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n568), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n510), .A2(new_n511), .ZN(new_n595));
  OAI21_X1  g0395(.A(KEYINPUT26), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT82), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n574), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n561), .A2(KEYINPUT82), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n573), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n339), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT83), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n600), .A2(KEYINPUT83), .A3(new_n339), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n603), .A2(new_n558), .A3(new_n567), .A4(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n600), .A2(G200), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n592), .A2(new_n579), .A3(new_n606), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n605), .A2(new_n510), .A3(new_n607), .A4(new_n511), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n596), .B1(KEYINPUT26), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n512), .A2(new_n476), .A3(new_n607), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n532), .A2(new_n540), .A3(new_n541), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n611), .B1(new_n450), .B2(new_n472), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n605), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  OR2_X1    g0413(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n590), .B1(new_n419), .B2(new_n615), .ZN(G369));
  NAND2_X1  g0416(.A1(new_n421), .A2(new_n211), .ZN(new_n617));
  XOR2_X1   g0417(.A(new_n617), .B(KEYINPUT84), .Z(new_n618));
  OR2_X1    g0418(.A1(new_n618), .A2(KEYINPUT27), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(KEYINPUT27), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(G213), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(G343), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n473), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g0424(.A(new_n624), .B(KEYINPUT85), .ZN(new_n625));
  INV_X1    g0425(.A(new_n623), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n626), .A2(new_n450), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n625), .B1(new_n477), .B2(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n628), .A2(KEYINPUT86), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(KEYINPUT86), .ZN(new_n630));
  OR2_X1    g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n541), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n537), .A2(new_n534), .ZN(new_n633));
  NOR3_X1   g0433(.A1(new_n632), .A2(new_n531), .A3(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n626), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n473), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n623), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n631), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n626), .A2(new_n539), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n542), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n643), .B1(new_n634), .B2(new_n642), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(G330), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n640), .A2(new_n647), .ZN(G399));
  INV_X1    g0448(.A(new_n206), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n649), .A2(G41), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(G1), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n548), .A2(G116), .ZN(new_n653));
  OAI22_X1  g0453(.A1(new_n652), .A2(new_n653), .B1(new_n214), .B2(new_n651), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n654), .B(KEYINPUT28), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT26), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n656), .B1(new_n594), .B2(new_n595), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT89), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n608), .B2(new_n656), .ZN(new_n659));
  INV_X1    g0459(.A(new_n604), .ZN(new_n660));
  AOI21_X1  g0460(.A(KEYINPUT83), .B1(new_n600), .B2(new_n339), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n580), .A2(new_n557), .B1(new_n290), .B2(new_n566), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n606), .A2(new_n579), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n662), .A2(new_n663), .B1(new_n664), .B2(new_n592), .ZN(new_n665));
  INV_X1    g0465(.A(new_n595), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n665), .A2(new_n666), .A3(KEYINPUT89), .A4(KEYINPUT26), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n657), .A2(new_n659), .A3(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(new_n613), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT29), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n669), .A2(new_n670), .A3(new_n626), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n614), .A2(new_n623), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n671), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n460), .A2(new_n465), .ZN(new_n674));
  OAI21_X1  g0474(.A(KEYINPUT87), .B1(new_n674), .B2(new_n575), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT87), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n566), .A2(new_n676), .A3(new_n460), .A4(new_n465), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n675), .A2(new_n538), .A3(new_n501), .A4(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT30), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n499), .A2(new_n470), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT88), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n499), .A2(KEYINPUT88), .A3(new_n470), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n530), .A2(new_n290), .A3(new_n600), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n499), .A2(new_n679), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n687), .A2(new_n538), .A3(new_n675), .A4(new_n677), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n680), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n626), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT31), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n689), .A2(KEYINPUT31), .A3(new_n626), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n583), .A2(new_n477), .A3(new_n626), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(G330), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n673), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n655), .B1(new_n699), .B2(G1), .ZN(G364));
  INV_X1    g0500(.A(new_n645), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n420), .A2(G20), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n271), .B1(new_n702), .B2(G45), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n650), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(G330), .B2(new_n644), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n210), .B1(G20), .B2(new_n339), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n290), .A2(new_n286), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT92), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n211), .B1(new_n711), .B2(G190), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n713), .A2(KEYINPUT94), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(KEYINPUT94), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(new_n479), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n211), .A2(G190), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n711), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(new_n317), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT32), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n290), .A2(G200), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n718), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n254), .B1(new_n723), .B2(new_n202), .ZN(new_n724));
  NAND3_X1  g0524(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G190), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n725), .A2(new_n353), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OAI22_X1  g0529(.A1(new_n727), .A2(new_n217), .B1(new_n729), .B2(new_n270), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n286), .A2(G179), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(new_n718), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  AOI211_X1 g0533(.A(new_n724), .B(new_n730), .C1(G107), .C2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n731), .A2(G20), .A3(G190), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n735), .A2(KEYINPUT93), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(KEYINPUT93), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n722), .A2(G20), .A3(G190), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT91), .ZN(new_n741));
  OR2_X1    g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI22_X1  g0544(.A1(new_n739), .A2(G87), .B1(G58), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n721), .A2(new_n734), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n717), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n254), .ZN(new_n748));
  INV_X1    g0548(.A(G303), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n748), .B1(new_n738), .B2(new_n749), .ZN(new_n750));
  XOR2_X1   g0550(.A(new_n750), .B(KEYINPUT95), .Z(new_n751));
  INV_X1    g0551(.A(new_n719), .ZN(new_n752));
  AOI22_X1  g0552(.A1(new_n752), .A2(G329), .B1(new_n744), .B2(G322), .ZN(new_n753));
  INV_X1    g0553(.A(G317), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n754), .A2(KEYINPUT33), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(KEYINPUT33), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n726), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n723), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G311), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n733), .A2(G283), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n728), .A2(G326), .ZN(new_n761));
  AND4_X1   g0561(.A1(new_n757), .A2(new_n759), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G294), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n753), .B(new_n762), .C1(new_n763), .C2(new_n712), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n751), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n708), .B1(new_n747), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n705), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n254), .A2(G355), .A3(new_n206), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n242), .A2(G45), .ZN(new_n769));
  XOR2_X1   g0569(.A(new_n769), .B(KEYINPUT90), .Z(new_n770));
  NOR2_X1   g0570(.A1(new_n649), .A2(new_n254), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(G45), .B2(new_n214), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n768), .B1(G116), .B2(new_n206), .C1(new_n770), .C2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G13), .A2(G33), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(G20), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n708), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n767), .B1(new_n773), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n766), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT96), .ZN(new_n780));
  INV_X1    g0580(.A(new_n776), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n780), .B1(new_n644), .B2(new_n781), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n707), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(G396));
  NAND2_X1  g0584(.A1(new_n415), .A2(new_n623), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n626), .A2(new_n403), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(new_n412), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n786), .B1(new_n416), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n672), .A2(new_n790), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n789), .B(new_n623), .C1(new_n609), .C2(new_n613), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n698), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n705), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n791), .A2(new_n698), .A3(new_n792), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n758), .A2(G159), .B1(G137), .B2(new_n728), .ZN(new_n797));
  INV_X1    g0597(.A(G150), .ZN(new_n798));
  INV_X1    g0598(.A(new_n744), .ZN(new_n799));
  INV_X1    g0599(.A(G143), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n797), .B1(new_n798), .B2(new_n727), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(KEYINPUT34), .ZN(new_n803));
  INV_X1    g0603(.A(G132), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n254), .B1(new_n217), .B2(new_n732), .C1(new_n719), .C2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(G50), .B2(new_n739), .ZN(new_n806));
  INV_X1    g0606(.A(G58), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n803), .B(new_n806), .C1(new_n807), .C2(new_n712), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n802), .A2(KEYINPUT34), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n752), .A2(G311), .B1(new_n744), .B2(G294), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n729), .A2(new_n749), .B1(new_n723), .B2(new_n436), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(G283), .B2(new_n726), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n812), .A2(KEYINPUT97), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(KEYINPUT97), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n748), .B1(new_n732), .B2(new_n219), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(new_n739), .B2(G107), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n810), .A2(new_n813), .A3(new_n814), .A4(new_n816), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n808), .A2(new_n809), .B1(new_n717), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n708), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n708), .A2(new_n774), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n767), .B1(new_n202), .B2(new_n820), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n819), .B(new_n821), .C1(new_n789), .C2(new_n775), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n796), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(G384));
  INV_X1    g0624(.A(new_n482), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n436), .B(new_n213), .C1(new_n825), .C2(KEYINPUT35), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(KEYINPUT35), .B2(new_n825), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT36), .Z(new_n828));
  NOR3_X1   g0628(.A1(new_n314), .A2(new_n202), .A3(new_n214), .ZN(new_n829));
  OR2_X1    g0629(.A1(new_n829), .A2(KEYINPUT98), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n829), .A2(KEYINPUT98), .B1(new_n270), .B2(G68), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n271), .B(G13), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n828), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n299), .B1(new_n308), .B2(new_n310), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n834), .A2(new_n312), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n311), .A2(new_n269), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n325), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n622), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n356), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n837), .A2(new_n343), .ZN(new_n840));
  OAI21_X1  g0640(.A(KEYINPUT37), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n326), .B1(new_n343), .B2(new_n622), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n356), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n841), .B1(KEYINPUT37), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT102), .ZN(new_n845));
  INV_X1    g0645(.A(new_n838), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n845), .B1(new_n362), .B2(new_n846), .ZN(new_n847));
  AOI211_X1 g0647(.A(KEYINPUT102), .B(new_n838), .C1(new_n346), .C2(new_n361), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n844), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT38), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(KEYINPUT38), .B(new_n844), .C1(new_n847), .C2(new_n848), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT99), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n391), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n380), .A2(KEYINPUT99), .A3(new_n390), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n623), .A2(new_n393), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n395), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n855), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n857), .B1(new_n380), .B2(new_n395), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n860), .A2(KEYINPUT100), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n860), .A2(KEYINPUT100), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n859), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n789), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT104), .B1(new_n694), .B2(new_n695), .ZN(new_n865));
  INV_X1    g0665(.A(new_n488), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n499), .A2(G200), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n866), .A2(new_n502), .A3(new_n867), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n634), .A2(new_n595), .A3(new_n536), .A4(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n869), .A2(new_n594), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n473), .A2(new_n476), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n870), .A2(new_n871), .A3(new_n623), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT104), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n872), .A2(new_n873), .A3(new_n692), .A4(new_n693), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n865), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n864), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n853), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT40), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n621), .B1(new_n322), .B2(new_n325), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n326), .A2(new_n343), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT18), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n326), .A2(new_n295), .A3(new_n343), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n880), .B1(new_n588), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT103), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n842), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT37), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n843), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n842), .A2(KEYINPUT103), .A3(KEYINPUT37), .A4(new_n356), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n885), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n850), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n852), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(KEYINPUT105), .ZN(new_n894));
  NOR3_X1   g0694(.A1(new_n864), .A2(new_n875), .A3(new_n878), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT105), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n852), .A2(new_n892), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n894), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n879), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n418), .A2(new_n865), .A3(new_n874), .ZN(new_n901));
  OAI21_X1  g0701(.A(G330), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n902), .B1(new_n900), .B2(new_n901), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n792), .A2(new_n785), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n863), .ZN(new_n905));
  OR2_X1    g0705(.A1(new_n905), .A2(KEYINPUT101), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(KEYINPUT101), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n906), .A2(new_n853), .A3(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT39), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n893), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n851), .A2(KEYINPUT39), .A3(new_n852), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n855), .A2(new_n856), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n912), .A2(new_n626), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n910), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n884), .A2(new_n621), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n908), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n673), .A2(new_n418), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n917), .A2(new_n590), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n916), .B(new_n918), .Z(new_n919));
  NAND2_X1  g0719(.A1(new_n903), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n903), .A2(new_n919), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT106), .ZN(new_n922));
  OAI221_X1 g0722(.A(new_n920), .B1(new_n271), .B2(new_n702), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n921), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n924), .A2(KEYINPUT106), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n833), .B1(new_n923), .B2(new_n925), .ZN(G367));
  OAI21_X1  g0726(.A(new_n512), .B1(new_n866), .B2(new_n623), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n666), .A2(new_n626), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n631), .A2(new_n635), .A3(new_n929), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n930), .A2(KEYINPUT42), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n929), .B(KEYINPUT108), .Z(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n637), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n626), .B1(new_n933), .B2(new_n595), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n934), .B1(new_n930), .B2(KEYINPUT42), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n623), .A2(new_n592), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n605), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n665), .B2(new_n936), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n938), .B(KEYINPUT107), .Z(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n931), .A2(new_n935), .B1(KEYINPUT43), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n940), .A2(KEYINPUT43), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n941), .B(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n646), .A2(new_n932), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n943), .B(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n650), .B(KEYINPUT41), .Z(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT109), .B1(new_n640), .B2(new_n929), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT109), .ZN(new_n948));
  INV_X1    g0748(.A(new_n929), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n639), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT44), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n639), .A2(new_n949), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT45), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n947), .A2(KEYINPUT44), .A3(new_n950), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n646), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n953), .A2(new_n955), .A3(new_n647), .A4(new_n956), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n631), .B(new_n635), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(new_n701), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n958), .A2(new_n699), .A3(new_n959), .A4(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n946), .B1(new_n962), .B2(new_n699), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n945), .B1(new_n963), .B2(new_n704), .ZN(new_n964));
  INV_X1    g0764(.A(new_n771), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n777), .B1(new_n206), .B2(new_n400), .C1(new_n235), .C2(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n767), .B1(new_n966), .B2(KEYINPUT110), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(KEYINPUT110), .B2(new_n966), .ZN(new_n968));
  INV_X1    g0768(.A(new_n716), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(G68), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n254), .B1(new_n732), .B2(new_n202), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n727), .A2(new_n317), .B1(new_n729), .B2(new_n800), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n971), .B(new_n972), .C1(G50), .C2(new_n758), .ZN(new_n973));
  INV_X1    g0773(.A(G137), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n719), .A2(new_n974), .B1(new_n738), .B2(new_n807), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(G150), .B2(new_n744), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n970), .A2(new_n973), .A3(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n738), .A2(new_n436), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT46), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n748), .B1(new_n732), .B2(new_n479), .ZN(new_n980));
  XNOR2_X1  g0780(.A(KEYINPUT111), .B(G311), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n763), .A2(new_n727), .B1(new_n729), .B2(new_n981), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n980), .B(new_n982), .C1(G283), .C2(new_n758), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n752), .A2(G317), .B1(new_n744), .B2(G303), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n983), .B(new_n984), .C1(new_n408), .C2(new_n712), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n977), .B1(new_n979), .B2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT47), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n968), .B1(new_n987), .B2(new_n708), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n940), .B2(new_n781), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n964), .A2(new_n989), .ZN(G387));
  AOI21_X1  g0790(.A(new_n651), .B1(new_n961), .B2(new_n699), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n699), .B2(new_n961), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n641), .A2(new_n776), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n771), .B1(new_n232), .B2(new_n245), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n653), .A2(new_n206), .A3(new_n254), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AOI211_X1 g0796(.A(G45), .B(new_n653), .C1(G68), .C2(G77), .ZN(new_n997));
  OAI21_X1  g0797(.A(KEYINPUT50), .B1(new_n265), .B2(G50), .ZN(new_n998));
  OR3_X1    g0798(.A1(new_n265), .A2(KEYINPUT50), .A3(G50), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n996), .A2(new_n1000), .B1(new_n422), .B2(new_n649), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n777), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n705), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT112), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n969), .A2(new_n554), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n254), .B1(new_n732), .B2(new_n479), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n317), .A2(new_n729), .B1(new_n727), .B2(new_n265), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n1006), .B(new_n1007), .C1(G68), .C2(new_n758), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n799), .A2(new_n270), .B1(new_n202), .B2(new_n738), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(G150), .B2(new_n752), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1005), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n752), .A2(G326), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n254), .B1(new_n733), .B2(G116), .ZN(new_n1013));
  INV_X1    g0813(.A(G283), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n712), .A2(new_n1014), .B1(new_n738), .B2(new_n763), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n758), .A2(G303), .B1(G322), .B2(new_n728), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(new_n727), .B2(new_n981), .C1(new_n799), .C2(new_n754), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT48), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1015), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n1018), .B2(new_n1017), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT49), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1012), .B(new_n1013), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1022));
  AND2_X1   g0822(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1011), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1024), .A2(KEYINPUT113), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n708), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n1024), .B2(KEYINPUT113), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1004), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n961), .A2(new_n704), .B1(new_n993), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n992), .A2(new_n1029), .ZN(G393));
  NAND2_X1  g0830(.A1(new_n958), .A2(new_n959), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n961), .A2(new_n699), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1033), .A2(new_n650), .A3(new_n962), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n958), .A2(new_n704), .A3(new_n959), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n239), .A2(new_n771), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1036), .B(new_n777), .C1(new_n479), .C2(new_n206), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n705), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT114), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n744), .A2(G311), .B1(G317), .B2(new_n728), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT52), .Z(new_n1041));
  NAND2_X1  g0841(.A1(new_n713), .A2(G116), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n748), .B1(new_n723), .B2(new_n763), .C1(new_n422), .C2(new_n732), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(G303), .B2(new_n726), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(G322), .A2(new_n752), .B1(new_n739), .B2(G283), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n744), .A2(G159), .B1(G150), .B2(new_n728), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT51), .Z(new_n1048));
  AOI22_X1  g0848(.A1(new_n758), .A2(new_n323), .B1(G50), .B2(new_n726), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1048), .B(new_n1049), .C1(new_n202), .C2(new_n716), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n748), .B1(new_n733), .B2(G87), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n738), .B2(new_n217), .C1(new_n800), .C2(new_n719), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT115), .Z(new_n1053));
  OAI21_X1  g0853(.A(new_n1046), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1039), .B1(new_n1054), .B2(new_n708), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n932), .B2(new_n781), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n1035), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1034), .A2(new_n1057), .ZN(G390));
  AOI21_X1  g0858(.A(new_n913), .B1(new_n904), .B2(new_n863), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n910), .B2(new_n911), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT116), .ZN(new_n1062));
  AND3_X1   g0862(.A1(new_n852), .A2(new_n892), .A3(new_n896), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n896), .B1(new_n852), .B2(new_n892), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n788), .A2(new_n416), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n623), .B(new_n1066), .C1(new_n668), .C2(new_n613), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n785), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n913), .B1(new_n1068), .B2(new_n863), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1062), .B1(new_n1065), .B2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n894), .A2(new_n1069), .A3(new_n1062), .A4(new_n897), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1061), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n865), .A2(G330), .A3(new_n874), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n864), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1077));
  NOR3_X1   g0877(.A1(new_n696), .A2(new_n697), .A3(new_n790), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n864), .A2(new_n1074), .B1(new_n1078), .B2(new_n863), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n904), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT117), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n865), .A2(new_n874), .A3(new_n1081), .A4(G330), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n1082), .A2(new_n789), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1074), .A2(KEYINPUT117), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n863), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n698), .A2(new_n789), .A3(new_n863), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1068), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n1085), .A2(KEYINPUT118), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT118), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n863), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1084), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1082), .A2(new_n789), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1091), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1088), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1090), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1080), .B1(new_n1089), .B2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n894), .A2(new_n897), .A3(new_n1069), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(KEYINPUT116), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n1071), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1100), .A2(new_n1061), .A3(new_n1086), .ZN(new_n1101));
  OR2_X1    g0901(.A1(new_n419), .A2(new_n1074), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n918), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1077), .A2(new_n1097), .A3(new_n1101), .A4(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1075), .B1(new_n1100), .B2(new_n1061), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1086), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1107), .B(new_n1060), .C1(new_n1099), .C2(new_n1071), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1080), .ZN(new_n1109));
  OAI21_X1  g0909(.A(KEYINPUT118), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1094), .A2(new_n1090), .A3(new_n1095), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1109), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n1106), .A2(new_n1108), .B1(new_n1112), .B2(new_n1103), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1105), .A2(new_n1113), .A3(new_n650), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n910), .A2(new_n911), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n774), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n820), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n705), .B1(new_n323), .B2(new_n1118), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n729), .A2(new_n1014), .B1(new_n732), .B2(new_n217), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n719), .A2(new_n763), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1120), .B(new_n1121), .C1(G116), .C2(new_n744), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n408), .A2(new_n727), .B1(new_n479), .B2(new_n723), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT119), .Z(new_n1124));
  OAI211_X1 g0924(.A(new_n1122), .B(new_n1124), .C1(new_n716), .C2(new_n202), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n748), .B1(new_n738), .B2(new_n219), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT120), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n738), .A2(new_n798), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT53), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(KEYINPUT54), .B(G143), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n254), .B1(new_n723), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(G128), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n727), .A2(new_n974), .B1(new_n729), .B2(new_n1132), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1131), .B(new_n1133), .C1(G50), .C2(new_n733), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n752), .A2(G125), .B1(new_n744), .B2(G132), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1129), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n716), .A2(new_n317), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n1125), .A2(new_n1127), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1119), .B1(new_n1138), .B2(new_n708), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1115), .A2(new_n704), .B1(new_n1117), .B2(new_n1139), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1114), .A2(KEYINPUT121), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(KEYINPUT121), .B1(new_n1114), .B2(new_n1140), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(G378));
  OAI21_X1  g0943(.A(new_n970), .B1(new_n436), .B2(new_n729), .ZN(new_n1144));
  XOR2_X1   g0944(.A(new_n1144), .B(KEYINPUT122), .Z(new_n1145));
  OAI22_X1  g0945(.A1(new_n719), .A2(new_n1014), .B1(new_n738), .B2(new_n202), .ZN(new_n1146));
  AOI211_X1 g0946(.A(G41), .B(new_n254), .C1(new_n758), .C2(new_n554), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n1147), .B1(new_n807), .B2(new_n732), .C1(new_n479), .C2(new_n727), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n1146), .B(new_n1148), .C1(G107), .C2(new_n744), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1145), .A2(KEYINPUT58), .A3(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n270), .B1(G33), .B2(G41), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n748), .B2(new_n244), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n304), .B(new_n244), .C1(new_n732), .C2(new_n317), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n799), .A2(new_n1132), .B1(new_n738), .B2(new_n1130), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n758), .A2(G137), .B1(G125), .B2(new_n728), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n804), .B2(new_n727), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n716), .B2(new_n798), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1158), .A2(KEYINPUT59), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1153), .B(new_n1159), .C1(G124), .C2(new_n752), .ZN(new_n1160));
  OR2_X1    g0960(.A1(new_n1158), .A2(KEYINPUT59), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1152), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1150), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(KEYINPUT58), .B1(new_n1145), .B2(new_n1149), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n708), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n767), .B1(new_n270), .B2(new_n820), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n622), .A2(new_n281), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n294), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n293), .A2(new_n281), .A3(new_n622), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1168), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1165), .B(new_n1166), .C1(new_n1175), .C2(new_n775), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n879), .A2(G330), .A3(new_n898), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1175), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1175), .A2(new_n879), .A3(G330), .A4(new_n898), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n916), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1180), .A2(new_n916), .A3(new_n1181), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1177), .B1(new_n1186), .B2(new_n704), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1103), .B1(new_n1115), .B2(new_n1097), .ZN(new_n1188));
  AND3_X1   g0988(.A1(new_n1180), .A2(new_n916), .A3(new_n1181), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n916), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1190));
  OAI21_X1  g0990(.A(KEYINPUT57), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n650), .B1(new_n1188), .B2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1060), .B1(new_n1099), .B2(new_n1071), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1101), .B1(new_n1193), .B2(new_n1075), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1104), .B1(new_n1194), .B2(new_n1112), .ZN(new_n1195));
  AOI21_X1  g0995(.A(KEYINPUT57), .B1(new_n1195), .B2(new_n1186), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1187), .B1(new_n1192), .B2(new_n1196), .ZN(G375));
  NAND2_X1  g0997(.A1(new_n1097), .A2(new_n1104), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1112), .A2(new_n1103), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n946), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n254), .B1(new_n732), .B2(new_n807), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n804), .A2(new_n729), .B1(new_n727), .B2(new_n1130), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1202), .B(new_n1203), .C1(G150), .C2(new_n758), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n719), .A2(new_n1132), .B1(new_n738), .B2(new_n317), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(G137), .B2(new_n744), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1204), .B(new_n1206), .C1(new_n716), .C2(new_n270), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n727), .A2(new_n436), .B1(new_n729), .B2(new_n763), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n748), .B1(new_n732), .B2(new_n202), .C1(new_n408), .C2(new_n723), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1208), .B(new_n1209), .C1(G283), .C2(new_n744), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1005), .A2(new_n1210), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n719), .A2(new_n749), .B1(new_n738), .B2(new_n479), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n1212), .B(KEYINPUT123), .Z(new_n1213));
  OAI21_X1  g1013(.A(new_n1207), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT124), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1026), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n1215), .B2(new_n1214), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1217), .B(new_n705), .C1(G68), .C2(new_n1118), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1091), .B2(new_n774), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n1097), .B2(new_n704), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1201), .A2(new_n1220), .ZN(G381));
  NAND3_X1  g1021(.A1(new_n992), .A2(new_n783), .A3(new_n1029), .ZN(new_n1222));
  OR2_X1    g1022(.A1(new_n1222), .A2(G384), .ZN(new_n1223));
  OR3_X1    g1023(.A1(G390), .A2(G381), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1114), .A2(new_n1140), .ZN(new_n1225));
  OR4_X1    g1025(.A1(G387), .A2(new_n1224), .A3(new_n1225), .A4(G375), .ZN(G407));
  NOR2_X1   g1026(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1176), .B1(new_n1227), .B2(new_n703), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT57), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n1188), .B2(new_n1227), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1229), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n651), .B1(new_n1231), .B2(new_n1195), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1228), .B1(new_n1230), .B2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1225), .ZN(new_n1234));
  INV_X1    g1034(.A(G213), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1235), .A2(G343), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1233), .A2(new_n1234), .A3(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(G407), .A2(G213), .A3(new_n1237), .ZN(G409));
  INV_X1    g1038(.A(KEYINPUT127), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1195), .A2(new_n1186), .A3(new_n1200), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1240), .A2(new_n1187), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1241), .A2(new_n1225), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT121), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1225), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1114), .A2(new_n1140), .A3(KEYINPUT121), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(KEYINPUT125), .B1(new_n1246), .B2(G375), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT125), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(G378), .A2(new_n1248), .A3(new_n1233), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1242), .B1(new_n1247), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1198), .A2(KEYINPUT60), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n1251), .A2(new_n1199), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n650), .B1(new_n1251), .B2(new_n1199), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1220), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1254), .B(G384), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(new_n1250), .A2(new_n1236), .A3(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1239), .B1(new_n1257), .B2(KEYINPUT62), .ZN(new_n1258));
  NOR3_X1   g1058(.A1(new_n1246), .A2(G375), .A3(KEYINPUT125), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1248), .B1(G378), .B2(new_n1233), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n1259), .A2(new_n1260), .B1(new_n1225), .B2(new_n1241), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT126), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1236), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1261), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(KEYINPUT126), .B1(new_n1250), .B2(new_n1236), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1264), .A2(new_n1265), .A3(KEYINPUT62), .A4(new_n1255), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1261), .A2(new_n1263), .A3(new_n1255), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT62), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1267), .A2(KEYINPUT127), .A3(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1258), .A2(new_n1266), .A3(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1236), .A2(G2897), .ZN(new_n1272));
  XOR2_X1   g1072(.A(new_n1255), .B(new_n1272), .Z(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT61), .B1(new_n1271), .B2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1270), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(G393), .A2(G396), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1222), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(new_n1034), .B2(new_n1057), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1034), .A2(new_n1057), .A3(new_n1277), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1279), .A2(new_n964), .A3(new_n989), .A4(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1280), .ZN(new_n1282));
  OAI21_X1  g1082(.A(G387), .B1(new_n1282), .B2(new_n1278), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1275), .A2(new_n1284), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1284), .A2(KEYINPUT61), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1264), .A2(new_n1265), .A3(KEYINPUT63), .A4(new_n1255), .ZN(new_n1287));
  OR2_X1    g1087(.A1(new_n1257), .A2(KEYINPUT63), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1273), .B1(new_n1236), .B2(new_n1250), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1286), .A2(new_n1287), .A3(new_n1288), .A4(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1285), .A2(new_n1290), .ZN(G405));
  AOI22_X1  g1091(.A1(new_n1247), .A2(new_n1249), .B1(new_n1234), .B2(G375), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1292), .B(new_n1256), .ZN(new_n1293));
  XNOR2_X1  g1093(.A(new_n1284), .B(new_n1293), .ZN(G402));
endmodule


