//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 1 1 0 1 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 1 0 0 1 1 1 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 0 1 0 1 1 0 1 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n788, new_n789, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979;
  INV_X1    g000(.A(G183gat), .ZN(new_n202));
  INV_X1    g001(.A(G190gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND3_X1  g003(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AOI21_X1  g005(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT25), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G169gat), .ZN(new_n209));
  INV_X1    g008(.A(G176gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(new_n210), .A3(KEYINPUT23), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n212), .B1(G169gat), .B2(G176gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n211), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT66), .B1(new_n208), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n215), .ZN(new_n217));
  INV_X1    g016(.A(new_n207), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n218), .A2(new_n205), .A3(new_n204), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT66), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n217), .A2(new_n219), .A3(new_n220), .A4(KEYINPUT25), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n216), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n223));
  NOR2_X1   g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224));
  AND2_X1   g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n224), .B1(new_n225), .B2(KEYINPUT24), .ZN(new_n226));
  AOI22_X1  g025(.A1(new_n215), .A2(new_n223), .B1(new_n226), .B2(new_n218), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n211), .A2(new_n213), .A3(KEYINPUT65), .A4(new_n214), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT25), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n222), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(new_n214), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT69), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT69), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n231), .A2(new_n234), .A3(new_n214), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT26), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n236), .A2(new_n209), .A3(new_n210), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n233), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n225), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT27), .ZN(new_n241));
  AOI21_X1  g040(.A(G190gat), .B1(new_n241), .B2(G183gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n202), .A2(KEYINPUT27), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n242), .A2(KEYINPUT28), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n246), .B1(new_n241), .B2(G183gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n202), .A2(KEYINPUT67), .A3(KEYINPUT27), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(new_n242), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT28), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n245), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n249), .A2(KEYINPUT68), .A3(new_n250), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n240), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G120gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(G113gat), .ZN(new_n257));
  INV_X1    g056(.A(G113gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(G120gat), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT1), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G127gat), .B(G134gat), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT70), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AND2_X1   g061(.A1(G127gat), .A2(G134gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(G127gat), .A2(G134gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n266));
  XNOR2_X1  g065(.A(G113gat), .B(G120gat), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n265), .B(new_n266), .C1(new_n267), .C2(KEYINPUT1), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(KEYINPUT71), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n258), .A2(G120gat), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n256), .A2(G113gat), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT1), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n270), .A2(new_n274), .A3(new_n275), .A4(new_n261), .ZN(new_n276));
  AND3_X1   g075(.A1(new_n269), .A2(KEYINPUT72), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT72), .B1(new_n269), .B2(new_n276), .ZN(new_n278));
  OAI22_X1  g077(.A1(new_n230), .A2(new_n255), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n215), .A2(new_n223), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n280), .A2(new_n228), .A3(new_n219), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT25), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n283), .A2(new_n216), .A3(new_n221), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n251), .A2(new_n252), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(new_n254), .A3(new_n244), .ZN(new_n286));
  INV_X1    g085(.A(new_n240), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n275), .B1(new_n272), .B2(new_n273), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n266), .B1(new_n289), .B2(new_n265), .ZN(new_n290));
  NOR3_X1   g089(.A1(new_n260), .A2(KEYINPUT70), .A3(new_n261), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n276), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n269), .A2(KEYINPUT72), .A3(new_n276), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n284), .A2(new_n288), .A3(new_n294), .A4(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G227gat), .A2(G233gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n297), .B(KEYINPUT64), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n279), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G15gat), .B(G43gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(G71gat), .B(G99gat), .ZN(new_n301));
  XOR2_X1   g100(.A(new_n300), .B(new_n301), .Z(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT33), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n299), .A2(KEYINPUT32), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT73), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n299), .A2(KEYINPUT73), .A3(KEYINPUT32), .A4(new_n303), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT33), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n299), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n302), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n310), .B1(new_n299), .B2(KEYINPUT32), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n306), .A2(new_n307), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT34), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n279), .A2(new_n296), .ZN(new_n314));
  INV_X1    g113(.A(new_n298), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  AOI211_X1 g115(.A(KEYINPUT34), .B(new_n298), .C1(new_n279), .C2(new_n296), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n318), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n320), .B1(new_n312), .B2(KEYINPUT74), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n307), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n311), .A2(new_n309), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n322), .A2(KEYINPUT74), .A3(new_n323), .ZN(new_n324));
  OAI211_X1 g123(.A(KEYINPUT36), .B(new_n319), .C1(new_n321), .C2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT75), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n322), .A2(new_n323), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT74), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n312), .A2(KEYINPUT74), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n330), .A2(new_n320), .A3(new_n331), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n332), .A2(KEYINPUT75), .A3(KEYINPUT36), .A4(new_n319), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT36), .ZN(new_n334));
  INV_X1    g133(.A(new_n319), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n312), .A2(new_n318), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n327), .A2(new_n333), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(G225gat), .A2(G233gat), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(G141gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(G148gat), .ZN(new_n342));
  INV_X1    g141(.A(G148gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(G141gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT2), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(G155gat), .ZN(new_n348));
  INV_X1    g147(.A(G162gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G155gat), .A2(G162gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n347), .A2(KEYINPUT79), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT79), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT2), .B1(new_n342), .B2(new_n344), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n355), .B1(new_n356), .B2(new_n352), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n343), .A2(G141gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT80), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT80), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n342), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n360), .A2(new_n344), .A3(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n351), .B1(new_n350), .B2(KEYINPUT2), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n358), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n366), .A2(new_n292), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n365), .A2(new_n358), .B1(new_n269), .B2(new_n276), .ZN(new_n368));
  OAI211_X1 g167(.A(KEYINPUT82), .B(new_n340), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT5), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n366), .A2(new_n292), .ZN(new_n371));
  AOI22_X1  g170(.A1(new_n354), .A2(new_n357), .B1(new_n363), .B2(new_n364), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n372), .A2(new_n276), .A3(new_n269), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n339), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n374), .A2(KEYINPUT82), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT83), .B1(new_n370), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n340), .B1(new_n367), .B2(new_n368), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT82), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT83), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n379), .A2(new_n380), .A3(KEYINPUT5), .A4(new_n369), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT81), .ZN(new_n383));
  AND3_X1   g182(.A1(new_n358), .A2(new_n383), .A3(new_n365), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n383), .B1(new_n358), .B2(new_n365), .ZN(new_n385));
  OAI22_X1  g184(.A1(new_n384), .A2(new_n385), .B1(new_n277), .B2(new_n278), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT4), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n388), .A2(new_n340), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT3), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n372), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(new_n292), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n372), .A2(new_n390), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT4), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n373), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n389), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n382), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G1gat), .B(G29gat), .ZN(new_n398));
  INV_X1    g197(.A(G85gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT0), .B(G57gat), .ZN(new_n401));
  XOR2_X1   g200(.A(new_n400), .B(new_n401), .Z(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n387), .ZN(new_n404));
  INV_X1    g203(.A(new_n393), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n372), .A2(new_n390), .B1(new_n276), .B2(new_n269), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n405), .A2(new_n406), .B1(new_n367), .B2(KEYINPUT4), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  NOR3_X1   g207(.A1(new_n408), .A2(KEYINPUT5), .A3(new_n340), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n397), .A2(new_n403), .A3(new_n410), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n376), .A2(new_n381), .B1(new_n389), .B2(new_n395), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n402), .B1(new_n412), .B2(new_n409), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT6), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n411), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  OAI211_X1 g214(.A(KEYINPUT6), .B(new_n402), .C1(new_n412), .C2(new_n409), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(G226gat), .A2(G233gat), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n230), .A2(new_n255), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n418), .B1(new_n419), .B2(KEYINPUT29), .ZN(new_n420));
  INV_X1    g219(.A(G211gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT76), .B(G218gat), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT22), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G197gat), .B(G204gat), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n421), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n425), .A2(KEYINPUT22), .A3(new_n421), .ZN(new_n427));
  OR3_X1    g226(.A1(new_n426), .A2(G218gat), .A3(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(G218gat), .B1(new_n426), .B2(new_n427), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT77), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n284), .A2(new_n288), .ZN(new_n433));
  INV_X1    g232(.A(new_n418), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI211_X1 g234(.A(KEYINPUT77), .B(new_n418), .C1(new_n284), .C2(new_n288), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n420), .B(new_n431), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT78), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n419), .A2(new_n418), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT29), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n434), .B1(new_n433), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n430), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n437), .A2(new_n438), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n438), .B1(new_n437), .B2(new_n442), .ZN(new_n444));
  XNOR2_X1  g243(.A(G8gat), .B(G36gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(G64gat), .B(G92gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NOR3_X1   g247(.A1(new_n443), .A2(new_n444), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n437), .A2(new_n442), .A3(new_n448), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT30), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n437), .A2(new_n442), .A3(KEYINPUT30), .A4(new_n448), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n417), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n428), .A2(new_n440), .A3(new_n429), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT3), .B1(new_n457), .B2(KEYINPUT85), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n458), .B1(KEYINPUT85), .B2(new_n457), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n366), .ZN(new_n460));
  NAND2_X1  g259(.A1(G228gat), .A2(G233gat), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n391), .A2(new_n440), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n430), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n460), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n457), .A2(new_n390), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n384), .A2(new_n385), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n464), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT84), .B1(new_n469), .B2(new_n461), .ZN(new_n470));
  AOI22_X1  g269(.A1(new_n466), .A2(new_n467), .B1(new_n430), .B2(new_n463), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT84), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n471), .A2(new_n472), .A3(new_n462), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n465), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  XOR2_X1   g273(.A(G78gat), .B(G106gat), .Z(new_n475));
  XNOR2_X1  g274(.A(new_n475), .B(G22gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(KEYINPUT31), .B(G50gat), .ZN(new_n477));
  XOR2_X1   g276(.A(new_n476), .B(new_n477), .Z(new_n478));
  XNOR2_X1  g277(.A(new_n474), .B(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n456), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT88), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT37), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n439), .A2(new_n441), .A3(new_n430), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT77), .B1(new_n419), .B2(new_n418), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n433), .A2(new_n432), .A3(new_n434), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n431), .B1(new_n486), .B2(new_n420), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n483), .B1(new_n487), .B2(KEYINPUT87), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT87), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n441), .B1(new_n484), .B2(new_n485), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n489), .B1(new_n490), .B2(new_n431), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n482), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n437), .A2(new_n442), .A3(new_n482), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n448), .A2(KEYINPUT38), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n481), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n483), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n420), .B1(new_n435), .B2(new_n436), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n498), .A2(KEYINPUT87), .A3(new_n430), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n491), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT37), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n501), .A2(KEYINPUT88), .A3(new_n493), .A4(new_n494), .ZN(new_n502));
  NOR3_X1   g301(.A1(new_n443), .A2(new_n444), .A3(new_n482), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n493), .A2(new_n447), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT38), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n496), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n415), .A2(new_n416), .A3(new_n450), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT86), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT40), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT39), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n372), .B(new_n383), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n294), .A2(new_n295), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT4), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OAI22_X1  g313(.A1(new_n392), .A2(new_n393), .B1(new_n387), .B2(new_n373), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n511), .B(new_n340), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n403), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n371), .A2(new_n373), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT39), .B1(new_n518), .B2(new_n340), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n519), .B1(new_n408), .B2(new_n340), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n510), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n408), .A2(new_n340), .ZN(new_n522));
  INV_X1    g321(.A(new_n519), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n524), .A2(KEYINPUT40), .A3(new_n403), .A4(new_n516), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n413), .A2(new_n521), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n509), .B1(new_n455), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n478), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n474), .B(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n437), .A2(new_n442), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT78), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n437), .A2(new_n442), .A3(new_n438), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(new_n532), .A3(new_n447), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n533), .A2(new_n453), .A3(new_n452), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n525), .A2(new_n521), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n534), .A2(KEYINPUT86), .A3(new_n535), .A4(new_n413), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n527), .A2(new_n529), .A3(new_n536), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n338), .B(new_n480), .C1(new_n508), .C2(new_n537), .ZN(new_n538));
  NOR3_X1   g337(.A1(new_n479), .A2(new_n336), .A3(new_n335), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT35), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n539), .A2(new_n540), .A3(new_n417), .A4(new_n455), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n529), .A2(new_n332), .A3(new_n319), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT35), .B1(new_n456), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n538), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G15gat), .B(G22gat), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT16), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n546), .B1(new_n547), .B2(G1gat), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n548), .B1(G1gat), .B2(new_n546), .ZN(new_n549));
  INV_X1    g348(.A(G8gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT21), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT9), .ZN(new_n553));
  INV_X1    g352(.A(G71gat), .ZN(new_n554));
  INV_X1    g353(.A(G78gat), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OR2_X1    g355(.A1(new_n556), .A2(KEYINPUT92), .ZN(new_n557));
  XNOR2_X1  g356(.A(G71gat), .B(G78gat), .ZN(new_n558));
  XOR2_X1   g357(.A(G57gat), .B(G64gat), .Z(new_n559));
  NAND2_X1  g358(.A1(new_n556), .A2(KEYINPUT92), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .A4(new_n560), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n559), .A2(KEYINPUT9), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n561), .B1(new_n558), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n551), .B1(new_n552), .B2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT93), .ZN(new_n565));
  AND2_X1   g364(.A1(G231gat), .A2(G233gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n563), .A2(new_n552), .ZN(new_n568));
  XOR2_X1   g367(.A(G127gat), .B(G155gat), .Z(new_n569));
  XOR2_X1   g368(.A(new_n568), .B(new_n569), .Z(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n567), .B(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(G183gat), .B(G211gat), .Z(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n573), .B(new_n574), .Z(new_n575));
  XOR2_X1   g374(.A(new_n572), .B(new_n575), .Z(new_n576));
  NAND2_X1  g375(.A1(G85gat), .A2(G92gat), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n577), .B(KEYINPUT7), .Z(new_n578));
  XOR2_X1   g377(.A(KEYINPUT96), .B(G92gat), .Z(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(new_n399), .ZN(new_n580));
  INV_X1    g379(.A(G99gat), .ZN(new_n581));
  INV_X1    g380(.A(G106gat), .ZN(new_n582));
  OAI21_X1  g381(.A(KEYINPUT95), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT95), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n584), .A2(G99gat), .A3(G106gat), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n583), .A2(KEYINPUT8), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n580), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT97), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n580), .A2(KEYINPUT97), .A3(new_n586), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n578), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  XOR2_X1   g390(.A(G99gat), .B(G106gat), .Z(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n594), .B(KEYINPUT98), .Z(new_n595));
  OR3_X1    g394(.A1(new_n591), .A2(KEYINPUT99), .A3(new_n593), .ZN(new_n596));
  OAI21_X1  g395(.A(KEYINPUT99), .B1(new_n591), .B2(new_n593), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n563), .B1(new_n595), .B2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT10), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n594), .B(KEYINPUT98), .ZN(new_n601));
  OAI21_X1  g400(.A(KEYINPUT102), .B1(new_n591), .B2(new_n593), .ZN(new_n602));
  NOR3_X1   g401(.A1(new_n591), .A2(KEYINPUT102), .A3(new_n593), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n603), .A2(new_n563), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n601), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n599), .A2(new_n600), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n598), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n563), .A2(new_n600), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n607), .A2(new_n601), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(G230gat), .ZN(new_n611));
  INV_X1    g410(.A(G233gat), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G120gat), .B(G148gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(G176gat), .B(G204gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  AND2_X1   g418(.A1(new_n599), .A2(new_n605), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n615), .B(new_n619), .C1(new_n614), .C2(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n614), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n613), .B1(new_n606), .B2(new_n609), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n618), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n607), .A2(new_n601), .ZN(new_n627));
  XNOR2_X1  g426(.A(G43gat), .B(G50gat), .ZN(new_n628));
  NOR2_X1   g427(.A1(G29gat), .A2(G36gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT14), .ZN(new_n630));
  INV_X1    g429(.A(G29gat), .ZN(new_n631));
  INV_X1    g430(.A(G36gat), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI211_X1 g432(.A(KEYINPUT15), .B(new_n628), .C1(new_n630), .C2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n630), .B(KEYINPUT91), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n636));
  XOR2_X1   g435(.A(KEYINPUT90), .B(G50gat), .Z(new_n637));
  OAI21_X1  g436(.A(new_n636), .B1(new_n637), .B2(G43gat), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n633), .B1(new_n628), .B2(KEYINPUT15), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n634), .B1(new_n635), .B2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT17), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n627), .A2(KEYINPUT100), .A3(new_n642), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n607), .A2(new_n641), .A3(new_n601), .ZN(new_n648));
  NAND3_X1  g447(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G190gat), .B(G218gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT101), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT94), .ZN(new_n656));
  XNOR2_X1  g455(.A(G134gat), .B(G162gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n653), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n647), .A2(new_n659), .A3(new_n650), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n654), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n658), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n647), .A2(new_n659), .A3(new_n650), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n659), .B1(new_n647), .B2(new_n650), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n576), .A2(new_n626), .A3(new_n661), .A4(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n642), .A2(new_n551), .ZN(new_n667));
  NAND2_X1  g466(.A1(G229gat), .A2(G233gat), .ZN(new_n668));
  INV_X1    g467(.A(new_n551), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n641), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n667), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT18), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n641), .B(new_n551), .Z(new_n675));
  XOR2_X1   g474(.A(new_n668), .B(KEYINPUT13), .Z(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n673), .A2(new_n674), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n679));
  XNOR2_X1  g478(.A(G113gat), .B(G141gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g480(.A(G169gat), .B(G197gat), .Z(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT12), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n678), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n673), .A2(new_n684), .A3(new_n674), .A4(new_n677), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n666), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n545), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n417), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g494(.A1(new_n691), .A2(new_n455), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT42), .B1(new_n696), .B2(new_n550), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT16), .B(G8gat), .Z(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  MUX2_X1   g498(.A(KEYINPUT42), .B(new_n697), .S(new_n699), .Z(G1325gat));
  NOR2_X1   g499(.A1(new_n335), .A2(new_n336), .ZN(new_n701));
  AOI21_X1  g500(.A(G15gat), .B1(new_n692), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT103), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  INV_X1    g504(.A(new_n338), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n692), .A2(G15gat), .A3(new_n706), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n704), .A2(new_n705), .A3(new_n707), .ZN(G1326gat));
  NOR2_X1   g507(.A1(new_n691), .A2(new_n529), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT43), .B(G22gat), .Z(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1327gat));
  NAND2_X1  g510(.A1(new_n665), .A2(new_n661), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n713), .B1(new_n538), .B2(new_n544), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n576), .A2(new_n625), .A3(new_n689), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n718), .A2(new_n631), .A3(new_n693), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT45), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n712), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n545), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n538), .A2(new_n544), .A3(KEYINPUT104), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n722), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n714), .A2(new_n721), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n716), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT105), .ZN(new_n729));
  INV_X1    g528(.A(new_n722), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n538), .A2(KEYINPUT104), .A3(new_n544), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT104), .B1(new_n538), .B2(new_n544), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n715), .A2(KEYINPUT44), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT105), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n735), .A2(new_n736), .A3(new_n716), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n417), .B1(new_n729), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n720), .B1(new_n738), .B2(new_n631), .ZN(G1328gat));
  NAND3_X1  g538(.A1(new_n718), .A2(new_n632), .A3(new_n534), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n740), .B(KEYINPUT46), .Z(new_n741));
  AOI21_X1  g540(.A(new_n455), .B1(new_n729), .B2(new_n737), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n741), .B1(new_n742), .B2(new_n632), .ZN(G1329gat));
  AOI21_X1  g542(.A(new_n338), .B1(new_n729), .B2(new_n737), .ZN(new_n744));
  INV_X1    g543(.A(G43gat), .ZN(new_n745));
  OAI21_X1  g544(.A(KEYINPUT107), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n736), .B1(new_n735), .B2(new_n716), .ZN(new_n747));
  AOI211_X1 g546(.A(KEYINPUT105), .B(new_n717), .C1(new_n733), .C2(new_n734), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n706), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT107), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n749), .A2(new_n750), .A3(G43gat), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n718), .A2(new_n745), .A3(new_n701), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n746), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(G43gat), .B1(new_n728), .B2(new_n338), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n756), .A2(KEYINPUT47), .A3(new_n752), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n757), .ZN(G1330gat));
  OAI21_X1  g557(.A(new_n637), .B1(new_n728), .B2(new_n529), .ZN(new_n759));
  INV_X1    g558(.A(new_n637), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n718), .A2(new_n479), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n759), .A2(KEYINPUT48), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n761), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n479), .B1(new_n747), .B2(new_n748), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n763), .B1(new_n764), .B2(new_n637), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n762), .B1(new_n765), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g565(.A1(new_n724), .A2(new_n725), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n572), .B(new_n575), .ZN(new_n768));
  NOR4_X1   g567(.A1(new_n626), .A2(new_n712), .A3(new_n688), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n693), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(G57gat), .ZN(G1332gat));
  OR2_X1    g572(.A1(new_n534), .A2(KEYINPUT108), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n534), .A2(KEYINPUT108), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n776), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n771), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT109), .ZN(new_n779));
  NOR2_X1   g578(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n779), .B(new_n780), .ZN(G1333gat));
  INV_X1    g580(.A(new_n701), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n554), .B1(new_n770), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n706), .A2(G71gat), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n783), .B1(new_n770), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g584(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(G1334gat));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n479), .ZN(new_n788));
  XOR2_X1   g587(.A(KEYINPUT111), .B(G78gat), .Z(new_n789));
  XNOR2_X1  g588(.A(new_n788), .B(new_n789), .ZN(G1335gat));
  NOR2_X1   g589(.A1(new_n576), .A2(new_n688), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n735), .A2(new_n625), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(G85gat), .B1(new_n792), .B2(new_n417), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n714), .A2(new_n791), .ZN(new_n794));
  OR2_X1    g593(.A1(new_n794), .A2(KEYINPUT51), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(KEYINPUT51), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n795), .A2(new_n625), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n693), .A2(new_n399), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n793), .B1(new_n797), .B2(new_n798), .ZN(G1336gat));
  INV_X1    g598(.A(new_n792), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n579), .B1(new_n800), .B2(new_n534), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n801), .A2(KEYINPUT112), .ZN(new_n802));
  OR3_X1    g601(.A1(new_n797), .A2(G92gat), .A3(new_n776), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n803), .B1(new_n801), .B2(KEYINPUT112), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT52), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n792), .A2(new_n776), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n803), .B(new_n806), .C1(new_n579), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n805), .A2(new_n808), .ZN(G1337gat));
  OAI21_X1  g608(.A(G99gat), .B1(new_n792), .B2(new_n338), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n701), .A2(new_n581), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n810), .B1(new_n797), .B2(new_n811), .ZN(G1338gat));
  OAI21_X1  g611(.A(new_n582), .B1(new_n797), .B2(new_n529), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n479), .A2(G106gat), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n792), .B2(new_n814), .ZN(new_n815));
  XOR2_X1   g614(.A(new_n815), .B(KEYINPUT53), .Z(G1339gat));
  AOI21_X1  g615(.A(new_n668), .B1(new_n667), .B2(new_n670), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n675), .A2(new_n676), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n683), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OR2_X1    g618(.A1(new_n819), .A2(KEYINPUT114), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(KEYINPUT114), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n820), .A2(new_n687), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n822), .B1(new_n621), .B2(new_n624), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n712), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n606), .A2(new_n613), .A3(new_n609), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n826), .A2(new_n623), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n610), .A2(new_n827), .A3(new_n614), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n618), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n825), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n619), .B1(new_n623), .B2(new_n827), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n615), .A2(KEYINPUT54), .ZN(new_n833));
  OAI211_X1 g632(.A(KEYINPUT55), .B(new_n832), .C1(new_n833), .C2(new_n826), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n831), .A2(new_n834), .A3(new_n688), .A4(new_n621), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n824), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n822), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n831), .A2(new_n834), .A3(new_n621), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n712), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n836), .A2(new_n839), .A3(new_n768), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT113), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n841), .B1(new_n666), .B2(new_n688), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n712), .A2(new_n768), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n843), .A2(KEYINPUT113), .A3(new_n689), .A4(new_n626), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n840), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n845), .A2(new_n539), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(new_n693), .A3(new_n776), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT115), .ZN(new_n848));
  OAI21_X1  g647(.A(G113gat), .B1(new_n848), .B2(new_n689), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n845), .A2(new_n693), .ZN(new_n850));
  INV_X1    g649(.A(new_n542), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n776), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n688), .A2(new_n258), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n849), .B1(new_n853), .B2(new_n854), .ZN(G1340gat));
  OAI21_X1  g654(.A(G120gat), .B1(new_n848), .B2(new_n626), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n625), .A2(new_n256), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n856), .B1(new_n853), .B2(new_n857), .ZN(G1341gat));
  INV_X1    g657(.A(G127gat), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n848), .A2(new_n859), .A3(new_n768), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n852), .A2(new_n576), .A3(new_n776), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n860), .B1(new_n859), .B2(new_n861), .ZN(G1342gat));
  INV_X1    g661(.A(G134gat), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n713), .A2(new_n534), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n852), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  XOR2_X1   g664(.A(new_n865), .B(KEYINPUT56), .Z(new_n866));
  OAI21_X1  g665(.A(G134gat), .B1(new_n848), .B2(new_n713), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(G1343gat));
  INV_X1    g667(.A(KEYINPUT58), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n845), .A2(new_n479), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XOR2_X1   g672(.A(KEYINPUT116), .B(KEYINPUT57), .Z(new_n874));
  NAND2_X1  g673(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n776), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n706), .A2(new_n417), .A3(new_n876), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n873), .A2(new_n688), .A3(new_n875), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(G141gat), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n706), .A2(new_n529), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n850), .A2(KEYINPUT118), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n845), .A2(new_n693), .A3(new_n880), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT118), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n876), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n689), .A2(G141gat), .ZN(new_n886));
  AND3_X1   g685(.A1(new_n885), .A2(KEYINPUT119), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(KEYINPUT119), .B1(new_n885), .B2(new_n886), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n869), .B(new_n879), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT117), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n871), .A2(new_n877), .A3(new_n886), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n879), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n890), .B1(new_n892), .B2(KEYINPUT58), .ZN(new_n893));
  AOI211_X1 g692(.A(KEYINPUT117), .B(new_n869), .C1(new_n879), .C2(new_n891), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n889), .B1(new_n893), .B2(new_n894), .ZN(G1344gat));
  NAND3_X1  g694(.A1(new_n885), .A2(new_n343), .A3(new_n625), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n873), .A2(new_n875), .A3(new_n877), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n897), .A2(new_n626), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n898), .A2(KEYINPUT59), .A3(new_n343), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n845), .A2(new_n479), .A3(new_n874), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n836), .A2(new_n839), .A3(new_n768), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n666), .A2(new_n688), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n479), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI22_X1  g703(.A1(new_n901), .A2(KEYINPUT121), .B1(new_n904), .B2(new_n872), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT121), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n845), .A2(new_n906), .A3(new_n479), .A4(new_n874), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n626), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n877), .B(KEYINPUT120), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n900), .B1(new_n910), .B2(G148gat), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n896), .B1(new_n899), .B2(new_n911), .ZN(G1345gat));
  AOI21_X1  g711(.A(G155gat), .B1(new_n885), .B2(new_n576), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n897), .A2(new_n348), .A3(new_n768), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n913), .A2(new_n914), .ZN(G1346gat));
  OAI21_X1  g714(.A(G162gat), .B1(new_n897), .B2(new_n713), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n881), .A2(new_n884), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n917), .A2(new_n349), .A3(new_n864), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1347gat));
  NOR2_X1   g718(.A1(new_n693), .A2(new_n455), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n846), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(G169gat), .B1(new_n921), .B2(new_n689), .ZN(new_n922));
  AND3_X1   g721(.A1(new_n845), .A2(new_n417), .A3(new_n876), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(new_n851), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n688), .A2(new_n209), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(G1348gat));
  NOR3_X1   g725(.A1(new_n921), .A2(new_n210), .A3(new_n626), .ZN(new_n927));
  INV_X1    g726(.A(new_n924), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n625), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n927), .B1(new_n929), .B2(new_n210), .ZN(G1349gat));
  NAND2_X1  g729(.A1(new_n241), .A2(G183gat), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n928), .A2(new_n243), .A3(new_n931), .A4(new_n576), .ZN(new_n932));
  INV_X1    g731(.A(new_n921), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(KEYINPUT122), .A3(new_n576), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(G183gat), .ZN(new_n935));
  AOI21_X1  g734(.A(KEYINPUT122), .B1(new_n933), .B2(new_n576), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n932), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(KEYINPUT60), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT60), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n939), .B(new_n932), .C1(new_n935), .C2(new_n936), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(G1350gat));
  NAND3_X1  g740(.A1(new_n928), .A2(new_n203), .A3(new_n712), .ZN(new_n942));
  OAI21_X1  g741(.A(G190gat), .B1(new_n921), .B2(new_n713), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n943), .A2(KEYINPUT61), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n943), .A2(KEYINPUT61), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(G1351gat));
  NAND2_X1  g745(.A1(new_n923), .A2(new_n880), .ZN(new_n947));
  XOR2_X1   g746(.A(KEYINPUT123), .B(G197gat), .Z(new_n948));
  OR3_X1    g747(.A1(new_n947), .A2(new_n689), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n338), .A2(new_n920), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n950), .B1(new_n905), .B2(new_n907), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n951), .A2(new_n688), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n952), .A2(KEYINPUT124), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n948), .B1(new_n952), .B2(KEYINPUT124), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n949), .B1(new_n953), .B2(new_n954), .ZN(G1352gat));
  INV_X1    g754(.A(G204gat), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n923), .A2(new_n956), .A3(new_n625), .A4(new_n880), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT62), .ZN(new_n958));
  INV_X1    g757(.A(new_n950), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n956), .B1(new_n908), .B2(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT125), .ZN(new_n961));
  OR3_X1    g760(.A1(new_n958), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n961), .B1(new_n958), .B2(new_n960), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(G1353gat));
  NAND2_X1  g763(.A1(new_n951), .A2(new_n576), .ZN(new_n965));
  AND3_X1   g764(.A1(new_n965), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n966));
  AOI21_X1  g765(.A(KEYINPUT63), .B1(new_n965), .B2(G211gat), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n576), .A2(new_n421), .ZN(new_n968));
  OAI22_X1  g767(.A1(new_n966), .A2(new_n967), .B1(new_n947), .B2(new_n968), .ZN(G1354gat));
  INV_X1    g768(.A(G218gat), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n970), .B1(new_n947), .B2(new_n713), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n713), .A2(new_n422), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n972), .B1(new_n951), .B2(new_n973), .ZN(new_n974));
  AOI211_X1 g773(.A(KEYINPUT126), .B(new_n950), .C1(new_n905), .C2(new_n907), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n971), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(KEYINPUT127), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT127), .ZN(new_n978));
  OAI211_X1 g777(.A(new_n978), .B(new_n971), .C1(new_n974), .C2(new_n975), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n977), .A2(new_n979), .ZN(G1355gat));
endmodule


