//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n539, new_n541, new_n542, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n601, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1172,
    new_n1173, new_n1174, new_n1175;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT66), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  NAND2_X1  g031(.A1(G113), .A2(G2104), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT67), .ZN(new_n458));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  AND3_X1   g037(.A1(new_n460), .A2(new_n462), .A3(G125), .ZN(new_n463));
  OAI21_X1  g038(.A(G2105), .B1(new_n458), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND4_X1  g040(.A1(new_n460), .A2(new_n462), .A3(G137), .A4(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(G101), .A3(G2104), .ZN(new_n468));
  AND3_X1   g043(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n467), .B1(new_n466), .B2(new_n468), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(G160));
  NAND2_X1  g047(.A1(new_n460), .A2(new_n462), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(new_n465), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n473), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  OR2_X1    g056(.A1(G102), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G114), .C2(new_n465), .ZN(new_n483));
  NAND4_X1  g058(.A1(new_n460), .A2(new_n462), .A3(G126), .A4(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n460), .A2(new_n462), .A3(G138), .A4(new_n465), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT4), .ZN(new_n487));
  XNOR2_X1  g062(.A(KEYINPUT3), .B(G2104), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n488), .A2(new_n489), .A3(G138), .A4(new_n465), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n485), .B1(new_n487), .B2(new_n490), .ZN(G164));
  INV_X1    g066(.A(G543), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT5), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT5), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G543), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n493), .A2(new_n495), .A3(G62), .ZN(new_n496));
  NAND2_X1  g071(.A1(G75), .A2(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G651), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n493), .A2(new_n495), .ZN(new_n500));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT6), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G651), .ZN(new_n504));
  AND2_X1   g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n500), .A2(new_n505), .A3(G88), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n502), .A2(new_n504), .A3(G50), .A4(G543), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n499), .A2(KEYINPUT69), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT69), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n493), .A2(new_n495), .A3(new_n502), .A4(new_n504), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n507), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n501), .B1(new_n496), .B2(new_n497), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n508), .A2(new_n514), .ZN(G166));
  AND2_X1   g090(.A1(new_n505), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G51), .ZN(new_n517));
  INV_X1    g092(.A(new_n510), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G89), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n500), .A2(G63), .A3(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n517), .A2(new_n519), .A3(new_n520), .A4(new_n522), .ZN(G286));
  INV_X1    g098(.A(G286), .ZN(G168));
  AOI22_X1  g099(.A1(new_n500), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n501), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n505), .A2(G543), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT70), .B(G52), .ZN(new_n528));
  INV_X1    g103(.A(G90), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n527), .A2(new_n528), .B1(new_n529), .B2(new_n510), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n526), .A2(new_n530), .ZN(G171));
  AOI22_X1  g106(.A1(new_n500), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n501), .ZN(new_n533));
  INV_X1    g108(.A(G43), .ZN(new_n534));
  INV_X1    g109(.A(G81), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n527), .A2(new_n534), .B1(new_n535), .B2(new_n510), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G860), .ZN(G153));
  AND3_X1   g113(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G36), .ZN(G176));
  NAND2_X1  g115(.A1(G1), .A2(G3), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT8), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n539), .A2(new_n542), .ZN(G188));
  NAND3_X1  g118(.A1(new_n516), .A2(KEYINPUT9), .A3(G53), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT9), .ZN(new_n545));
  INV_X1    g120(.A(G53), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n527), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n518), .A2(G91), .ZN(new_n549));
  NAND2_X1  g124(.A1(G78), .A2(G543), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT71), .ZN(new_n551));
  OR2_X1    g126(.A1(KEYINPUT72), .A2(G65), .ZN(new_n552));
  NAND2_X1  g127(.A1(KEYINPUT72), .A2(G65), .ZN(new_n553));
  AND2_X1   g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n551), .B1(new_n500), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n549), .B1(new_n555), .B2(new_n501), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n548), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(G299));
  OR2_X1    g133(.A1(new_n526), .A2(new_n530), .ZN(G301));
  INV_X1    g134(.A(G166), .ZN(G303));
  OAI21_X1  g135(.A(G651), .B1(new_n500), .B2(G74), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n500), .A2(new_n505), .A3(G87), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n505), .A2(G49), .A3(G543), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(G288));
  INV_X1    g139(.A(G48), .ZN(new_n565));
  INV_X1    g140(.A(G86), .ZN(new_n566));
  OAI22_X1  g141(.A1(new_n527), .A2(new_n565), .B1(new_n566), .B2(new_n510), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n500), .A2(G61), .ZN(new_n568));
  NAND2_X1  g143(.A1(G73), .A2(G543), .ZN(new_n569));
  XOR2_X1   g144(.A(new_n569), .B(KEYINPUT73), .Z(new_n570));
  AOI21_X1  g145(.A(new_n501), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G305));
  AOI22_X1  g148(.A1(new_n500), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n574), .A2(new_n501), .ZN(new_n575));
  INV_X1    g150(.A(G47), .ZN(new_n576));
  XOR2_X1   g151(.A(KEYINPUT74), .B(G85), .Z(new_n577));
  OAI22_X1  g152(.A1(new_n527), .A2(new_n576), .B1(new_n510), .B2(new_n577), .ZN(new_n578));
  OR2_X1    g153(.A1(new_n575), .A2(new_n578), .ZN(G290));
  NAND2_X1  g154(.A1(G301), .A2(G868), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n500), .A2(G66), .ZN(new_n581));
  NAND2_X1  g156(.A1(G79), .A2(G543), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT77), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(KEYINPUT78), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(KEYINPUT78), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n585), .A2(G651), .A3(new_n586), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n527), .A2(KEYINPUT76), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n527), .A2(KEYINPUT76), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n588), .A2(G54), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n518), .A2(G92), .ZN(new_n591));
  XOR2_X1   g166(.A(KEYINPUT75), .B(KEYINPUT10), .Z(new_n592));
  XNOR2_X1  g167(.A(new_n591), .B(new_n592), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n587), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n580), .B1(new_n595), .B2(G868), .ZN(G284));
  OAI21_X1  g171(.A(new_n580), .B1(new_n595), .B2(G868), .ZN(G321));
  NAND2_X1  g172(.A1(G286), .A2(G868), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n598), .B1(new_n557), .B2(G868), .ZN(G297));
  OAI21_X1  g174(.A(new_n598), .B1(new_n557), .B2(G868), .ZN(G280));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n595), .B1(new_n601), .B2(G860), .ZN(G148));
  NAND4_X1  g177(.A1(new_n587), .A2(new_n601), .A3(new_n590), .A4(new_n593), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G868), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(G868), .B2(new_n537), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g181(.A1(new_n465), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT12), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(KEYINPUT13), .Z(new_n609));
  NOR2_X1   g184(.A1(KEYINPUT79), .A2(G2100), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n474), .A2(G123), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n476), .A2(G135), .ZN(new_n613));
  OR2_X1    g188(.A1(G99), .A2(G2105), .ZN(new_n614));
  OAI211_X1 g189(.A(new_n614), .B(G2104), .C1(G111), .C2(new_n465), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n612), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(G2096), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n617), .A2(new_n618), .B1(KEYINPUT79), .B2(G2100), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n611), .B(new_n619), .C1(new_n618), .C2(new_n617), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT80), .Z(G156));
  XNOR2_X1  g196(.A(G2427), .B(G2438), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2430), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT15), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(G2435), .Z(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(KEYINPUT14), .ZN(new_n626));
  XOR2_X1   g201(.A(G1341), .B(G1348), .Z(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n626), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2451), .B(G2454), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT16), .B(G2443), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n626), .B(new_n627), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(new_n632), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT81), .B(G2446), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n634), .A2(new_n636), .A3(new_n638), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(G14), .A3(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(G401));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  XNOR2_X1  g219(.A(G2072), .B(G2078), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2067), .B(G2678), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT18), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n645), .B(KEYINPUT17), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(new_n644), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n645), .A2(new_n646), .ZN(new_n652));
  AOI211_X1 g227(.A(new_n644), .B(new_n652), .C1(new_n649), .C2(new_n646), .ZN(new_n653));
  AND2_X1   g228(.A1(new_n653), .A2(KEYINPUT82), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(KEYINPUT82), .ZN(new_n655));
  OAI221_X1 g230(.A(new_n648), .B1(new_n646), .B2(new_n651), .C1(new_n654), .C2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2100), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT83), .B(G2096), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(G227));
  XNOR2_X1  g234(.A(G1956), .B(G2474), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n660), .A2(KEYINPUT84), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(KEYINPUT84), .ZN(new_n662));
  XOR2_X1   g237(.A(G1961), .B(G1966), .Z(new_n663));
  AND3_X1   g238(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G1971), .B(G1976), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT20), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n663), .B1(new_n661), .B2(new_n662), .ZN(new_n669));
  AOI22_X1  g244(.A1(new_n667), .A2(new_n668), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  OR3_X1    g245(.A1(new_n664), .A2(new_n669), .A3(new_n666), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n670), .B(new_n671), .C1(new_n668), .C2(new_n667), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G1981), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1991), .B(G1996), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT86), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT21), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT22), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n673), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT85), .B(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(G229));
  AOI22_X1  g256(.A1(new_n488), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  AOI22_X1  g258(.A1(new_n683), .A2(G2105), .B1(new_n476), .B2(G139), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT25), .Z(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G29), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G29), .B2(G33), .ZN(new_n690));
  INV_X1    g265(.A(G2072), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(G29), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G26), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n474), .A2(G128), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n476), .A2(G140), .ZN(new_n696));
  OR2_X1    g271(.A1(G104), .A2(G2105), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n697), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n695), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n694), .B1(new_n700), .B2(new_n693), .ZN(new_n701));
  MUX2_X1   g276(.A(new_n694), .B(new_n701), .S(KEYINPUT28), .Z(new_n702));
  INV_X1    g277(.A(G2067), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n705), .A2(KEYINPUT23), .A3(G20), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT23), .ZN(new_n707));
  INV_X1    g282(.A(G20), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(G16), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n706), .B(new_n709), .C1(new_n557), .C2(new_n705), .ZN(new_n710));
  INV_X1    g285(.A(G1956), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT30), .B(G28), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n712), .A2(new_n713), .B1(new_n693), .B2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT31), .ZN(new_n716));
  OAI22_X1  g291(.A1(new_n616), .A2(new_n693), .B1(new_n716), .B2(G11), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n716), .B2(G11), .ZN(new_n718));
  AND4_X1   g293(.A1(new_n692), .A2(new_n704), .A3(new_n715), .A4(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(G286), .A2(new_n705), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(KEYINPUT94), .ZN(new_n721));
  OAI21_X1  g296(.A(KEYINPUT94), .B1(G16), .B2(G21), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n721), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G1966), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(G5), .A2(G16), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G171), .B2(G16), .ZN(new_n728));
  OAI221_X1 g303(.A(new_n726), .B1(G1961), .B2(new_n728), .C1(new_n691), .C2(new_n690), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n693), .A2(G35), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G162), .B2(new_n693), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT29), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G2090), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n693), .A2(G27), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G164), .B2(new_n693), .ZN(new_n735));
  INV_X1    g310(.A(G2078), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n705), .A2(G19), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n537), .B2(new_n705), .ZN(new_n739));
  AOI22_X1  g314(.A1(G1341), .A2(new_n739), .B1(new_n728), .B2(G1961), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n733), .A2(new_n737), .A3(new_n740), .ZN(new_n741));
  OAI22_X1  g316(.A1(new_n732), .A2(G2090), .B1(new_n724), .B2(new_n725), .ZN(new_n742));
  NOR3_X1   g317(.A1(new_n729), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n739), .A2(G1341), .ZN(new_n744));
  OAI21_X1  g319(.A(KEYINPUT93), .B1(G29), .B2(G32), .ZN(new_n745));
  AOI22_X1  g320(.A1(G129), .A2(new_n474), .B1(new_n476), .B2(G141), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n465), .A2(G105), .A3(G2104), .ZN(new_n747));
  NAND3_X1  g322(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT26), .Z(new_n749));
  NAND3_X1  g324(.A1(new_n746), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n750), .A2(KEYINPUT92), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(KEYINPUT92), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n745), .B1(new_n753), .B2(G29), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT27), .B(G1996), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n753), .A2(G29), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n755), .B(new_n757), .C1(KEYINPUT93), .C2(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n758), .A2(KEYINPUT93), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n756), .B1(new_n760), .B2(new_n754), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n719), .A2(new_n743), .A3(new_n744), .A4(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT34), .ZN(new_n764));
  NAND2_X1  g339(.A1(G166), .A2(G16), .ZN(new_n765));
  INV_X1    g340(.A(G1971), .ZN(new_n766));
  NOR2_X1   g341(.A1(G16), .A2(G22), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n765), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n705), .B1(new_n508), .B2(new_n514), .ZN(new_n770));
  OAI21_X1  g345(.A(G1971), .B1(new_n770), .B2(new_n767), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G1976), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT33), .ZN(new_n774));
  NAND2_X1  g349(.A1(G288), .A2(G16), .ZN(new_n775));
  INV_X1    g350(.A(G23), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n776), .A2(G16), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n774), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  AOI211_X1 g354(.A(KEYINPUT33), .B(new_n777), .C1(G288), .C2(G16), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n773), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n775), .A2(new_n778), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n782), .A2(KEYINPUT33), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n775), .A2(new_n774), .A3(new_n778), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n783), .A2(G1976), .A3(new_n784), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n772), .A2(new_n781), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n572), .A2(G16), .ZN(new_n787));
  OR2_X1    g362(.A1(G6), .A2(G16), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT32), .B(G1981), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n789), .B(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n764), .B1(new_n786), .B2(new_n792), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n785), .A2(new_n781), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n789), .B(new_n790), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n794), .A2(new_n795), .A3(KEYINPUT34), .A4(new_n772), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(G25), .A2(G29), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n474), .A2(G119), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n476), .A2(G131), .ZN(new_n800));
  OAI21_X1  g375(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n465), .A2(G107), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n799), .B(new_n800), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT87), .Z(new_n804));
  AOI21_X1  g379(.A(new_n798), .B1(new_n804), .B2(G29), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT35), .B(G1991), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT88), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n805), .B(new_n807), .ZN(new_n808));
  MUX2_X1   g383(.A(G24), .B(G290), .S(G16), .Z(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(G1986), .Z(new_n810));
  NAND3_X1  g385(.A1(new_n797), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT89), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n797), .A2(KEYINPUT89), .A3(new_n808), .A4(new_n810), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n813), .A2(KEYINPUT36), .A3(new_n814), .ZN(new_n815));
  AND3_X1   g390(.A1(new_n797), .A2(new_n808), .A3(new_n810), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT36), .ZN(new_n817));
  AOI21_X1  g392(.A(KEYINPUT90), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n763), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n813), .A2(KEYINPUT90), .A3(KEYINPUT36), .A4(new_n814), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n705), .A2(G4), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n595), .B2(new_n705), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT91), .B(G1348), .Z(new_n823));
  XOR2_X1   g398(.A(new_n822), .B(new_n823), .Z(new_n824));
  INV_X1    g399(.A(KEYINPUT24), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n825), .A2(G34), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(G34), .ZN(new_n827));
  AOI21_X1  g402(.A(G29), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(new_n471), .B2(G29), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(G2084), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n819), .A2(new_n820), .A3(new_n824), .A4(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(G311));
  NAND2_X1  g407(.A1(new_n831), .A2(KEYINPUT95), .ZN(new_n833));
  INV_X1    g408(.A(new_n830), .ZN(new_n834));
  AOI211_X1 g409(.A(new_n834), .B(new_n763), .C1(new_n815), .C2(new_n818), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT95), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n835), .A2(new_n836), .A3(new_n820), .A4(new_n824), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n833), .A2(new_n837), .ZN(G150));
  INV_X1    g413(.A(G55), .ZN(new_n839));
  INV_X1    g414(.A(G93), .ZN(new_n840));
  OAI22_X1  g415(.A1(new_n527), .A2(new_n839), .B1(new_n840), .B2(new_n510), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n500), .A2(G67), .ZN(new_n842));
  NAND2_X1  g417(.A1(G80), .A2(G543), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n501), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT96), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(KEYINPUT96), .B1(new_n841), .B2(new_n844), .ZN(new_n848));
  AND3_X1   g423(.A1(new_n847), .A2(new_n537), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n537), .B1(new_n847), .B2(new_n848), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT38), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n594), .A2(new_n601), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n853), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT39), .ZN(new_n857));
  OAI21_X1  g432(.A(KEYINPUT97), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(G860), .B1(new_n856), .B2(new_n857), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT97), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n854), .A2(new_n860), .A3(new_n855), .A4(KEYINPUT39), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n858), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT98), .ZN(new_n863));
  OAI21_X1  g438(.A(G860), .B1(new_n841), .B2(new_n844), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT37), .Z(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(G145));
  XNOR2_X1  g441(.A(new_n471), .B(new_n480), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n616), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n476), .A2(G142), .ZN(new_n869));
  OAI21_X1  g444(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n870), .A2(KEYINPUT100), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(KEYINPUT100), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n871), .B(new_n872), .C1(G118), .C2(new_n465), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n474), .A2(G130), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n869), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n875), .B(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n608), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n804), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n753), .A2(new_n688), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n751), .A2(new_n752), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n687), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n881), .A2(new_n699), .A3(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n487), .A2(new_n490), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(KEYINPUT99), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n483), .A2(new_n484), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT99), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n487), .A2(new_n490), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n887), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n699), .B1(new_n881), .B2(new_n883), .ZN(new_n892));
  NOR3_X1   g467(.A1(new_n885), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n487), .A2(new_n490), .A3(new_n889), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n889), .B1(new_n487), .B2(new_n490), .ZN(new_n895));
  NOR3_X1   g470(.A1(new_n894), .A2(new_n895), .A3(new_n485), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n881), .A2(new_n883), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(new_n700), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n896), .B1(new_n898), .B2(new_n884), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n880), .B1(new_n893), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n891), .B1(new_n885), .B2(new_n892), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n898), .A2(new_n896), .A3(new_n884), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n879), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n900), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n903), .A2(new_n904), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n868), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(G37), .ZN(new_n908));
  INV_X1    g483(.A(new_n868), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n900), .A2(new_n909), .A3(new_n903), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n907), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT40), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT40), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n907), .A2(new_n913), .A3(new_n908), .A4(new_n910), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(G395));
  NAND2_X1  g490(.A1(new_n595), .A2(new_n557), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n594), .A2(G299), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT41), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n595), .B(new_n601), .C1(new_n849), .C2(new_n850), .ZN(new_n921));
  INV_X1    g496(.A(new_n850), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n847), .A2(new_n537), .A3(new_n848), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n603), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n916), .A2(KEYINPUT41), .A3(new_n917), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n920), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT104), .B1(new_n925), .B2(new_n918), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n916), .A2(new_n917), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT104), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n929), .A2(new_n930), .A3(new_n924), .A4(new_n921), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n927), .A2(new_n928), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT42), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT42), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n927), .A2(new_n928), .A3(new_n931), .A4(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(KEYINPUT105), .ZN(new_n937));
  XNOR2_X1  g512(.A(G290), .B(G288), .ZN(new_n938));
  XNOR2_X1  g513(.A(G166), .B(new_n572), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n938), .B(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n933), .A2(new_n942), .A3(new_n935), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n937), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n941), .B1(new_n937), .B2(new_n943), .ZN(new_n945));
  OAI21_X1  g520(.A(G868), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OR2_X1    g521(.A1(new_n845), .A2(G868), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(G295));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n947), .ZN(G331));
  XNOR2_X1  g524(.A(G301), .B(G286), .ZN(new_n950));
  OR3_X1    g525(.A1(new_n950), .A2(new_n849), .A3(new_n850), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n950), .B1(new_n849), .B2(new_n850), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n920), .A2(new_n926), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n951), .A2(new_n918), .A3(new_n952), .ZN(new_n954));
  OR3_X1    g529(.A1(new_n953), .A2(new_n954), .A3(new_n940), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n940), .B1(new_n953), .B2(new_n954), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(new_n956), .A3(new_n908), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT43), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n955), .A2(new_n956), .A3(new_n959), .A4(new_n908), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT106), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT44), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT44), .ZN(new_n964));
  AOI211_X1 g539(.A(KEYINPUT106), .B(new_n964), .C1(new_n958), .C2(new_n960), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n963), .A2(new_n965), .ZN(G397));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(new_n896), .B2(G1384), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n464), .B(G40), .C1(new_n469), .C2(new_n470), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G1996), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n753), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n699), .B(new_n703), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n882), .A2(G1996), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n806), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n975), .B1(new_n804), .B2(new_n976), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n804), .A2(new_n976), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(G290), .A2(G1986), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(G290), .A2(G1986), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n970), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT120), .ZN(new_n984));
  AOI21_X1  g559(.A(G1384), .B1(new_n886), .B2(new_n888), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n969), .B1(KEYINPUT45), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(G1966), .B1(new_n968), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n988));
  INV_X1    g563(.A(G1384), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n891), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n886), .A2(new_n888), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n989), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n969), .B1(new_n992), .B2(KEYINPUT50), .ZN(new_n993));
  XNOR2_X1  g568(.A(KEYINPUT115), .B(G2084), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n990), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n984), .B1(new_n987), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n986), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT45), .B1(new_n891), .B2(new_n989), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n725), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n990), .A2(new_n993), .A3(new_n994), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n999), .A2(KEYINPUT120), .A3(new_n1000), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n996), .A2(new_n1001), .A3(G8), .A4(G286), .ZN(new_n1002));
  OAI21_X1  g577(.A(G8), .B1(new_n987), .B2(new_n995), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n1004));
  NAND2_X1  g579(.A1(G286), .A2(G8), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT122), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT122), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1003), .A2(new_n1008), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n996), .A2(G8), .A3(new_n1001), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n1005), .B(KEYINPUT121), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1004), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1002), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n891), .A2(KEYINPUT45), .A3(new_n989), .ZN(new_n1015));
  INV_X1    g590(.A(new_n969), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT107), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1017), .B(new_n967), .C1(G164), .C2(G1384), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT107), .B1(new_n985), .B2(KEYINPUT45), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1015), .A2(new_n1016), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT108), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n1018), .A2(new_n1016), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT108), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1022), .A2(new_n1023), .A3(new_n1015), .A4(new_n1019), .ZN(new_n1024));
  AOI21_X1  g599(.A(G1971), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n985), .A2(new_n988), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n896), .A2(G1384), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1016), .B(new_n1026), .C1(new_n1027), .C2(new_n988), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1028), .A2(G2090), .ZN(new_n1029));
  OAI21_X1  g604(.A(G8), .B1(new_n1025), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n1032));
  INV_X1    g607(.A(G8), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1032), .B1(G166), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1030), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1016), .A2(new_n891), .A3(new_n989), .ZN(new_n1038));
  INV_X1    g613(.A(G288), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(G1976), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1038), .A2(G8), .A3(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1039), .A2(G1976), .ZN(new_n1042));
  OR3_X1    g617(.A1(new_n1041), .A2(KEYINPUT52), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G1981), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT49), .B1(new_n572), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT49), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1046), .B(G1981), .C1(new_n567), .C2(new_n571), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n572), .A2(new_n1044), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1048), .A2(KEYINPUT111), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(KEYINPUT111), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1051), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1052));
  AND2_X1   g627(.A1(new_n1038), .A2(G8), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1050), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT110), .ZN(new_n1055));
  AND3_X1   g630(.A1(new_n1041), .A2(new_n1055), .A3(KEYINPUT52), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1055), .B1(new_n1041), .B2(KEYINPUT52), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1043), .B(new_n1054), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g634(.A(new_n1035), .B(KEYINPUT109), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n990), .A2(new_n993), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1061), .A2(G2090), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1060), .B(G8), .C1(new_n1025), .C2(new_n1062), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1037), .A2(new_n1059), .A3(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1021), .A2(new_n736), .A3(new_n1024), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n1066));
  INV_X1    g641(.A(G1961), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n1065), .A2(new_n1066), .B1(new_n1067), .B2(new_n1061), .ZN(new_n1068));
  XNOR2_X1  g643(.A(G301), .B(KEYINPUT54), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n736), .A2(KEYINPUT53), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT123), .ZN(new_n1072));
  XNOR2_X1  g647(.A(new_n969), .B(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n968), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1071), .B1(new_n1074), .B2(KEYINPUT124), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1074), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT124), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1076), .A2(new_n1077), .B1(KEYINPUT45), .B2(new_n1027), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n1075), .A2(KEYINPUT125), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT125), .B1(new_n1078), .B2(new_n1075), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1068), .B(new_n1070), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n968), .A2(new_n986), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1068), .B1(new_n1071), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n1069), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1014), .A2(new_n1064), .A3(new_n1081), .A4(new_n1084), .ZN(new_n1085));
  XOR2_X1   g660(.A(KEYINPUT117), .B(KEYINPUT58), .Z(new_n1086));
  XNOR2_X1  g661(.A(new_n1086), .B(G1341), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1038), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1088), .B1(new_n1020), .B2(G1996), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n537), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n1091));
  OR2_X1    g666(.A1(new_n1091), .A2(KEYINPUT118), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(KEYINPUT118), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1090), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1094), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1020), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT56), .B(G2072), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n1096), .A2(new_n1097), .B1(new_n1028), .B2(new_n711), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n557), .B(KEYINPUT57), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT61), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1102), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT61), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1104), .A2(new_n1105), .A3(new_n1100), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1095), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n823), .B1(new_n990), .B2(new_n993), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1038), .A2(G2067), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT116), .ZN(new_n1111));
  OR3_X1    g686(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1111), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT60), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1108), .B(new_n594), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1115), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n595), .B1(new_n1117), .B2(KEYINPUT119), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1116), .A2(new_n1118), .B1(KEYINPUT119), .B2(new_n1117), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1107), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1101), .A2(new_n594), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1102), .B1(new_n1122), .B2(new_n1114), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1085), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1014), .A2(KEYINPUT62), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1037), .A2(new_n1059), .A3(new_n1063), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1083), .A2(G171), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT62), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1129), .B(new_n1002), .C1(new_n1010), .C2(new_n1013), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1125), .A2(new_n1128), .A3(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1003), .A2(G286), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n766), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1062), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1033), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1059), .B(new_n1132), .C1(new_n1136), .C2(new_n1035), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT63), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1033), .B1(new_n999), .B2(new_n1000), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT63), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1139), .A2(new_n1140), .A3(G168), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1141), .B1(new_n1030), .B2(new_n1036), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1063), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1059), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  XOR2_X1   g719(.A(new_n1049), .B(KEYINPUT112), .Z(new_n1145));
  NAND2_X1  g720(.A1(new_n1039), .A2(new_n773), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(KEYINPUT113), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1145), .B1(new_n1054), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT114), .ZN(new_n1149));
  OR2_X1    g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1150), .A2(new_n1053), .A3(new_n1151), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1138), .A2(new_n1144), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1131), .A2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n983), .B1(new_n1124), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n970), .ZN(new_n1156));
  OR3_X1    g731(.A1(new_n979), .A2(KEYINPUT126), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n970), .A2(new_n982), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n1158), .B(KEYINPUT48), .ZN(new_n1159));
  OAI21_X1  g734(.A(KEYINPUT126), .B1(new_n979), .B2(new_n1156), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1157), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1156), .B1(new_n753), .B2(new_n973), .ZN(new_n1162));
  AND3_X1   g737(.A1(new_n970), .A2(KEYINPUT46), .A3(new_n971), .ZN(new_n1163));
  AOI21_X1  g738(.A(KEYINPUT46), .B1(new_n970), .B2(new_n971), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1165), .B(KEYINPUT47), .ZN(new_n1166));
  AOI22_X1  g741(.A1(new_n975), .A2(new_n978), .B1(new_n703), .B2(new_n700), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1167), .A2(new_n1156), .ZN(new_n1168));
  NOR3_X1   g743(.A1(new_n1161), .A2(new_n1166), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1155), .A2(new_n1169), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g745(.A(G319), .ZN(new_n1172));
  OR3_X1    g746(.A1(G227), .A2(KEYINPUT127), .A3(new_n1172), .ZN(new_n1173));
  AND3_X1   g747(.A1(new_n642), .A2(new_n1173), .A3(new_n680), .ZN(new_n1174));
  OAI21_X1  g748(.A(KEYINPUT127), .B1(G227), .B2(new_n1172), .ZN(new_n1175));
  NAND4_X1  g749(.A1(new_n911), .A2(new_n1174), .A3(new_n961), .A4(new_n1175), .ZN(G225));
  INV_X1    g750(.A(G225), .ZN(G308));
endmodule


