//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 0 1 1 0 0 1 0 1 1 0 0 1 0 0 1 0 1 0 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n529, new_n530, new_n531, new_n532, new_n533, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n547, new_n549, new_n550, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n561, new_n562,
    new_n564, new_n565, new_n566, new_n568, new_n569, new_n570, new_n571,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n583, new_n584, new_n585, new_n588, new_n589, new_n591,
    new_n592, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1114, new_n1115, new_n1116, new_n1117;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT64), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI211_X1 g038(.A(new_n461), .B(G125), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n461), .B1(new_n471), .B2(G125), .ZN(new_n472));
  OAI21_X1  g047(.A(G2105), .B1(new_n466), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(G137), .ZN(new_n474));
  NAND2_X1  g049(.A1(G101), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  AND2_X1   g055(.A1(new_n471), .A2(KEYINPUT66), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n471), .A2(KEYINPUT66), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(new_n477), .ZN(new_n484));
  MUX2_X1   g059(.A(G100), .B(G112), .S(G2105), .Z(new_n485));
  AOI22_X1  g060(.A1(new_n484), .A2(G124), .B1(G2104), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n483), .A2(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  NAND2_X1  g065(.A1(KEYINPUT4), .A2(G138), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n491), .B1(new_n469), .B2(new_n470), .ZN(new_n492));
  AND2_X1   g067(.A1(G102), .A2(G2104), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n477), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G126), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(new_n469), .B2(new_n470), .ZN(new_n496));
  AND2_X1   g071(.A1(G114), .A2(G2104), .ZN(new_n497));
  OAI21_X1  g072(.A(G2105), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g073(.A(G138), .B(new_n477), .C1(new_n462), .C2(new_n463), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n494), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  XNOR2_X1  g078(.A(KEYINPUT6), .B(G651), .ZN(new_n504));
  AND2_X1   g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT67), .ZN(new_n506));
  AND3_X1   g081(.A1(new_n505), .A2(new_n506), .A3(G50), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n506), .B1(new_n505), .B2(G50), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT68), .B1(new_n510), .B2(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT68), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(new_n513), .A3(G543), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n511), .A2(new_n514), .B1(KEYINPUT5), .B2(new_n510), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(new_n504), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n517), .A2(new_n520), .ZN(G166));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XOR2_X1   g097(.A(new_n522), .B(KEYINPUT7), .Z(new_n523));
  AND3_X1   g098(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n524));
  AOI211_X1 g099(.A(new_n523), .B(new_n524), .C1(G51), .C2(new_n505), .ZN(new_n525));
  INV_X1    g100(.A(G89), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n526), .B2(new_n516), .ZN(G286));
  INV_X1    g102(.A(G286), .ZN(G168));
  AOI22_X1  g103(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n519), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n505), .A2(G52), .ZN(new_n531));
  XOR2_X1   g106(.A(KEYINPUT69), .B(G90), .Z(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n516), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n530), .A2(new_n533), .ZN(G171));
  AOI22_X1  g109(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT70), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n535), .A2(new_n536), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n537), .A2(G651), .A3(new_n538), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n515), .A2(new_n504), .ZN(new_n540));
  XNOR2_X1  g115(.A(KEYINPUT71), .B(G81), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n540), .A2(new_n541), .B1(G43), .B2(new_n505), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT72), .ZN(G153));
  AND3_X1   g121(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G36), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n547), .A2(new_n550), .ZN(G188));
  AOI22_X1  g126(.A1(new_n515), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G91), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n552), .A2(new_n519), .B1(new_n553), .B2(new_n516), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n505), .A2(G53), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(G299));
  INV_X1    g133(.A(G171), .ZN(G301));
  INV_X1    g134(.A(G166), .ZN(G303));
  AOI22_X1  g135(.A1(new_n540), .A2(G87), .B1(G49), .B2(new_n505), .ZN(new_n561));
  OAI21_X1  g136(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(G288));
  NAND2_X1  g138(.A1(new_n505), .A2(G48), .ZN(new_n564));
  INV_X1    g139(.A(G86), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n515), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n566));
  OAI221_X1 g141(.A(new_n564), .B1(new_n516), .B2(new_n565), .C1(new_n566), .C2(new_n519), .ZN(G305));
  AOI22_X1  g142(.A1(new_n540), .A2(G85), .B1(G47), .B2(new_n505), .ZN(new_n568));
  XOR2_X1   g143(.A(new_n568), .B(KEYINPUT73), .Z(new_n569));
  AOI22_X1  g144(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n570));
  OR2_X1    g145(.A1(new_n570), .A2(new_n519), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(G290));
  NAND2_X1  g147(.A1(new_n540), .A2(G92), .ZN(new_n573));
  XOR2_X1   g148(.A(new_n573), .B(KEYINPUT10), .Z(new_n574));
  NAND2_X1  g149(.A1(new_n515), .A2(G66), .ZN(new_n575));
  INV_X1    g150(.A(G79), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n576), .B2(new_n510), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n577), .A2(G651), .B1(G54), .B2(new_n505), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n579), .A2(G868), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n580), .B1(G868), .B2(G171), .ZN(G284));
  AOI21_X1  g156(.A(new_n580), .B1(G868), .B2(G171), .ZN(G321));
  NAND2_X1  g157(.A1(G286), .A2(G868), .ZN(new_n583));
  XOR2_X1   g158(.A(new_n583), .B(KEYINPUT74), .Z(new_n584));
  INV_X1    g159(.A(G299), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(G868), .B2(new_n585), .ZN(G297));
  OAI21_X1  g161(.A(new_n584), .B1(G868), .B2(new_n585), .ZN(G280));
  AND2_X1   g162(.A1(new_n574), .A2(new_n578), .ZN(new_n588));
  INV_X1    g163(.A(G559), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n589), .B2(G860), .ZN(G148));
  NOR2_X1   g165(.A1(new_n543), .A2(G868), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n579), .A2(G559), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n591), .B1(new_n592), .B2(G868), .ZN(G323));
  XNOR2_X1  g168(.A(G323), .B(KEYINPUT11), .ZN(G282));
  MUX2_X1   g169(.A(G99), .B(G111), .S(G2105), .Z(new_n595));
  AOI22_X1  g170(.A1(new_n484), .A2(G123), .B1(G2104), .B2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(G135), .ZN(new_n597));
  INV_X1    g172(.A(new_n487), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(G2096), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n599), .B(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n477), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT12), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT13), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(G2100), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(G156));
  INV_X1    g181(.A(KEYINPUT14), .ZN(new_n607));
  XOR2_X1   g182(.A(KEYINPUT15), .B(G2435), .Z(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(G2438), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(G2427), .ZN(new_n610));
  INV_X1    g185(.A(G2430), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n607), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(new_n611), .B2(new_n610), .ZN(new_n613));
  XNOR2_X1  g188(.A(G2451), .B(G2454), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT16), .ZN(new_n615));
  XOR2_X1   g190(.A(G2443), .B(G2446), .Z(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(G1341), .B(G1348), .Z(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT75), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n617), .B(new_n619), .ZN(new_n620));
  OR2_X1    g195(.A1(new_n613), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n613), .A2(new_n620), .ZN(new_n622));
  AND3_X1   g197(.A1(new_n621), .A2(G14), .A3(new_n622), .ZN(G401));
  XOR2_X1   g198(.A(G2084), .B(G2090), .Z(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2067), .B(G2678), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(G2072), .B(G2078), .Z(new_n628));
  NOR3_X1   g203(.A1(new_n625), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT77), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT76), .B(KEYINPUT18), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT17), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n628), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n626), .B1(new_n634), .B2(new_n624), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n624), .ZN(new_n636));
  INV_X1    g211(.A(new_n628), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n633), .B1(new_n625), .B2(new_n627), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n635), .B(new_n636), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n632), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(new_n600), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2100), .ZN(G227));
  XNOR2_X1  g217(.A(G1961), .B(G1966), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT78), .ZN(new_n644));
  XOR2_X1   g219(.A(G1956), .B(G2474), .Z(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1971), .B(G1976), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT19), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(KEYINPUT79), .B(KEYINPUT20), .Z(new_n650));
  AND2_X1   g225(.A1(new_n646), .A2(new_n648), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n644), .A2(new_n645), .ZN(new_n652));
  AOI22_X1  g227(.A1(new_n649), .A2(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI221_X1 g228(.A(new_n653), .B1(new_n648), .B2(new_n652), .C1(new_n649), .C2(new_n650), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1991), .B(G1996), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1981), .B(G1986), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n656), .B(new_n659), .ZN(G229));
  MUX2_X1   g235(.A(G24), .B(G290), .S(G16), .Z(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT83), .B(G1986), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(KEYINPUT80), .B(G29), .Z(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n665), .A2(G25), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n484), .A2(G119), .ZN(new_n667));
  MUX2_X1   g242(.A(G95), .B(G107), .S(G2105), .Z(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(G2104), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(G131), .B2(new_n487), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n666), .B1(new_n671), .B2(new_n665), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT82), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT35), .B(G1991), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT81), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n673), .B(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(G16), .A2(G23), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT84), .ZN(new_n678));
  XNOR2_X1  g253(.A(G288), .B(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n677), .B1(new_n679), .B2(G16), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT33), .B(G1976), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n680), .B(new_n681), .Z(new_n682));
  NOR2_X1   g257(.A1(G6), .A2(G16), .ZN(new_n683));
  INV_X1    g258(.A(G305), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n683), .B1(new_n684), .B2(G16), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT32), .B(G1981), .Z(new_n686));
  XOR2_X1   g261(.A(new_n685), .B(new_n686), .Z(new_n687));
  NOR2_X1   g262(.A1(G16), .A2(G22), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(G166), .B2(G16), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1971), .ZN(new_n690));
  NOR3_X1   g265(.A1(new_n682), .A2(new_n687), .A3(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT34), .ZN(new_n692));
  AOI211_X1 g267(.A(new_n663), .B(new_n676), .C1(new_n691), .C2(new_n692), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT36), .ZN(new_n695));
  AOI22_X1  g270(.A1(new_n693), .A2(new_n694), .B1(KEYINPUT85), .B2(new_n695), .ZN(new_n696));
  OR3_X1    g271(.A1(new_n696), .A2(KEYINPUT85), .A3(new_n695), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(KEYINPUT85), .B2(new_n695), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n484), .A2(G129), .ZN(new_n699));
  NAND3_X1  g274(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT26), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  AND2_X1   g278(.A1(G105), .A2(G2104), .ZN(new_n704));
  AOI22_X1  g279(.A1(new_n702), .A2(new_n703), .B1(new_n477), .B2(new_n704), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n699), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n487), .A2(G141), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G29), .ZN(new_n709));
  NOR2_X1   g284(.A1(G29), .A2(G32), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n709), .B1(KEYINPUT92), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(KEYINPUT92), .B2(new_n709), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT27), .B(G1996), .Z(new_n713));
  XOR2_X1   g288(.A(new_n712), .B(new_n713), .Z(new_n714));
  INV_X1    g289(.A(G16), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G21), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G168), .B2(new_n715), .ZN(new_n717));
  INV_X1    g292(.A(G1966), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT31), .B(G11), .Z(new_n720));
  INV_X1    g295(.A(G28), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n721), .A2(KEYINPUT30), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT93), .Z(new_n723));
  AOI21_X1  g298(.A(G29), .B1(new_n721), .B2(KEYINPUT30), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n720), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n719), .B(new_n725), .C1(new_n599), .C2(new_n664), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n715), .A2(G5), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G171), .B2(new_n715), .ZN(new_n728));
  INV_X1    g303(.A(G2084), .ZN(new_n729));
  NOR2_X1   g304(.A1(KEYINPUT24), .A2(G34), .ZN(new_n730));
  AND2_X1   g305(.A1(KEYINPUT24), .A2(G34), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n664), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n479), .B2(new_n733), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n728), .A2(G1961), .B1(new_n729), .B2(new_n734), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n734), .A2(new_n729), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n735), .B(new_n736), .C1(G1961), .C2(new_n728), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n665), .A2(G27), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G164), .B2(new_n665), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT94), .B(G2078), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT91), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n743), .A2(new_n477), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n487), .A2(G139), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n477), .A2(G103), .A3(G2104), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT90), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT89), .B(KEYINPUT25), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  OAI211_X1 g324(.A(new_n745), .B(new_n749), .C1(new_n742), .C2(new_n744), .ZN(new_n750));
  MUX2_X1   g325(.A(G33), .B(new_n750), .S(G29), .Z(new_n751));
  AOI21_X1  g326(.A(new_n741), .B1(new_n751), .B2(G2072), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G2072), .B2(new_n751), .ZN(new_n753));
  NOR4_X1   g328(.A1(new_n714), .A2(new_n726), .A3(new_n737), .A4(new_n753), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n754), .A2(KEYINPUT95), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n754), .A2(KEYINPUT95), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n665), .A2(G35), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G162), .B2(new_n665), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT29), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G2090), .ZN(new_n760));
  NOR2_X1   g335(.A1(G16), .A2(G19), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n544), .B2(G16), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G1341), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n715), .A2(G20), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT23), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n585), .B2(new_n715), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(G1956), .Z(new_n768));
  NAND2_X1  g343(.A1(new_n664), .A2(G26), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT28), .Z(new_n770));
  NAND2_X1  g345(.A1(new_n484), .A2(G128), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT86), .Z(new_n772));
  MUX2_X1   g347(.A(G104), .B(G116), .S(G2105), .Z(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G2104), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT87), .Z(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n487), .B2(G140), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n770), .B1(new_n777), .B2(G29), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT88), .B(G2067), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(G4), .A2(G16), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n588), .B2(G16), .ZN(new_n782));
  INV_X1    g357(.A(G1348), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n764), .A2(new_n768), .A3(new_n780), .A4(new_n784), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n755), .A2(new_n756), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n697), .A2(new_n698), .A3(new_n786), .ZN(G150));
  INV_X1    g362(.A(G150), .ZN(G311));
  AOI22_X1  g363(.A1(new_n540), .A2(G93), .B1(G55), .B2(new_n505), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n519), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(G860), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT37), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n543), .B(new_n791), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT38), .Z(new_n795));
  NOR2_X1   g370(.A1(new_n579), .A2(new_n589), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n798), .A2(KEYINPUT39), .ZN(new_n799));
  INV_X1    g374(.A(G860), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n798), .B2(KEYINPUT39), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n793), .B1(new_n799), .B2(new_n801), .ZN(G145));
  XNOR2_X1  g377(.A(new_n671), .B(KEYINPUT97), .ZN(new_n803));
  MUX2_X1   g378(.A(G106), .B(G118), .S(G2105), .Z(new_n804));
  AOI22_X1  g379(.A1(new_n484), .A2(G130), .B1(G2104), .B2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(G142), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n805), .B1(new_n806), .B2(new_n598), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(new_n603), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n803), .B(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT96), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n502), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n494), .A2(new_n498), .A3(KEYINPUT96), .A4(new_n501), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n777), .B(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n809), .B(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n708), .B(new_n750), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n489), .B(G160), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(new_n599), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n817), .A2(new_n819), .ZN(new_n821));
  XOR2_X1   g396(.A(KEYINPUT98), .B(G37), .Z(new_n822));
  NAND3_X1  g397(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g399(.A1(new_n791), .A2(G868), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n588), .A2(G299), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(KEYINPUT99), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n579), .A2(new_n585), .ZN(new_n828));
  OR3_X1    g403(.A1(new_n579), .A2(KEYINPUT99), .A3(new_n585), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n794), .B(new_n592), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n826), .A2(new_n828), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT41), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n830), .B2(new_n835), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(new_n832), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n833), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT42), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(G290), .B(new_n679), .ZN(new_n842));
  XNOR2_X1  g417(.A(G166), .B(new_n684), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n841), .B(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n825), .B1(new_n845), .B2(G868), .ZN(G331));
  XNOR2_X1  g421(.A(G331), .B(KEYINPUT100), .ZN(G295));
  INV_X1    g422(.A(KEYINPUT44), .ZN(new_n848));
  XNOR2_X1  g423(.A(G286), .B(G301), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n794), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n837), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n831), .B2(new_n850), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n852), .A2(new_n844), .ZN(new_n853));
  INV_X1    g428(.A(G37), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n855), .B1(new_n844), .B2(new_n852), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT43), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n850), .A2(KEYINPUT41), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(new_n834), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n860), .B(new_n844), .C1(new_n830), .C2(new_n859), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n853), .A2(new_n822), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(KEYINPUT43), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n848), .B1(new_n858), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n856), .A2(KEYINPUT43), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n862), .A2(new_n857), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n864), .B1(new_n848), .B2(new_n867), .ZN(G397));
  INV_X1    g443(.A(G1384), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n502), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(KEYINPUT50), .ZN(new_n871));
  XOR2_X1   g446(.A(KEYINPUT103), .B(KEYINPUT50), .Z(new_n872));
  NAND3_X1  g447(.A1(new_n502), .A2(new_n869), .A3(new_n872), .ZN(new_n873));
  AND3_X1   g448(.A1(new_n473), .A2(G40), .A3(new_n478), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n871), .A2(new_n729), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT111), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n473), .A2(G40), .A3(new_n478), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n878), .B1(KEYINPUT50), .B2(new_n870), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n879), .A2(KEYINPUT111), .A3(new_n729), .A4(new_n873), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT45), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n870), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n869), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(new_n874), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(new_n718), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n877), .A2(new_n880), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT119), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n877), .A2(new_n880), .A3(new_n885), .A4(KEYINPUT119), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI211_X1 g465(.A(KEYINPUT51), .B(G8), .C1(new_n890), .C2(G286), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n886), .A2(G8), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT51), .ZN(new_n893));
  NAND2_X1  g468(.A1(G286), .A2(G8), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n894), .B1(new_n888), .B2(new_n889), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT120), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT120), .ZN(new_n900));
  AOI211_X1 g475(.A(new_n900), .B(new_n897), .C1(new_n891), .C2(new_n895), .ZN(new_n901));
  NOR3_X1   g476(.A1(new_n899), .A2(new_n901), .A3(KEYINPUT62), .ZN(new_n902));
  INV_X1    g477(.A(new_n870), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n874), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(G8), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(G1976), .ZN(new_n907));
  AOI21_X1  g482(.A(KEYINPUT52), .B1(G288), .B2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(G288), .B(KEYINPUT84), .ZN(new_n909));
  OAI211_X1 g484(.A(new_n906), .B(new_n908), .C1(new_n909), .C2(new_n907), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n905), .B1(new_n679), .B2(G1976), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT52), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT106), .B1(G305), .B2(G1981), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n564), .B1(new_n565), .B2(new_n516), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  OR2_X1    g491(.A1(new_n566), .A2(new_n519), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n918));
  INV_X1    g493(.A(G1981), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n916), .A2(new_n917), .A3(new_n918), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n915), .A2(KEYINPUT107), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT107), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n564), .B(new_n922), .C1(new_n565), .C2(new_n516), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n921), .A2(new_n917), .A3(new_n923), .ZN(new_n924));
  AOI22_X1  g499(.A1(new_n914), .A2(new_n920), .B1(new_n924), .B2(G1981), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n906), .B1(new_n925), .B2(KEYINPUT49), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n914), .A2(new_n920), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n924), .A2(G1981), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n927), .A2(KEYINPUT49), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT108), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n927), .A2(new_n928), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT49), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n925), .A2(KEYINPUT49), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n933), .A2(new_n934), .A3(new_n935), .A4(new_n906), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n913), .B1(new_n930), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n903), .A2(new_n872), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n874), .B1(KEYINPUT50), .B2(new_n870), .ZN(new_n939));
  NOR3_X1   g514(.A1(new_n938), .A2(new_n939), .A3(G2090), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n878), .B1(new_n881), .B2(new_n870), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n811), .A2(KEYINPUT45), .A3(new_n869), .A4(new_n812), .ZN(new_n942));
  AOI21_X1  g517(.A(G1971), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(G8), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(G8), .B1(new_n517), .B2(new_n520), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT55), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n945), .B(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n944), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n941), .A2(new_n942), .ZN(new_n950));
  INV_X1    g525(.A(G1971), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G2090), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n879), .A2(new_n953), .A3(new_n873), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n952), .A2(KEYINPUT104), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT104), .ZN(new_n956));
  AND4_X1   g531(.A1(new_n953), .A2(new_n871), .A3(new_n873), .A4(new_n874), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n956), .B1(new_n943), .B2(new_n957), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n955), .A2(new_n958), .A3(G8), .A4(new_n947), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n959), .A2(KEYINPUT105), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n959), .A2(KEYINPUT105), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n937), .B(new_n949), .C1(new_n960), .C2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT123), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n879), .A2(new_n873), .ZN(new_n965));
  OR2_X1    g540(.A1(new_n965), .A2(G1961), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT53), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n967), .A2(G2078), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n941), .A2(new_n883), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  XOR2_X1   g545(.A(KEYINPUT121), .B(KEYINPUT53), .Z(new_n971));
  OAI21_X1  g546(.A(new_n971), .B1(new_n950), .B2(G2078), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(G171), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT122), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT122), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n976), .B(G171), .C1(new_n970), .C2(new_n973), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n959), .B(KEYINPUT105), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n979), .A2(KEYINPUT123), .A3(new_n949), .A4(new_n937), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n964), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT124), .B1(new_n902), .B2(new_n981), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n964), .A2(new_n978), .A3(new_n980), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n896), .A2(new_n898), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n900), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT62), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n896), .A2(KEYINPUT120), .A3(new_n898), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT124), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n983), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n899), .A2(new_n901), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT125), .B1(new_n991), .B2(new_n986), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT125), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n993), .B(KEYINPUT62), .C1(new_n899), .C2(new_n901), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n982), .A2(new_n990), .A3(new_n992), .A4(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT63), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n892), .A2(G286), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n955), .A2(new_n958), .A3(G8), .ZN(new_n999));
  AOI211_X1 g574(.A(new_n996), .B(new_n998), .C1(new_n948), .C2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n1000), .A2(new_n979), .A3(new_n937), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n996), .B1(new_n962), .B2(new_n998), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n930), .A2(new_n936), .ZN(new_n1004));
  NOR2_X1   g579(.A1(G288), .A2(G1976), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n1004), .A2(new_n1005), .B1(new_n914), .B2(new_n920), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n1006), .A2(KEYINPUT110), .ZN(new_n1007));
  XOR2_X1   g582(.A(new_n905), .B(KEYINPUT109), .Z(new_n1008));
  AOI21_X1  g583(.A(new_n1008), .B1(new_n1006), .B2(KEYINPUT110), .ZN(new_n1009));
  INV_X1    g584(.A(new_n979), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n1007), .A2(new_n1009), .B1(new_n1010), .B2(new_n937), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1003), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n555), .A2(KEYINPUT113), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT57), .ZN(new_n1014));
  NAND3_X1  g589(.A1(G299), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n557), .B(new_n555), .C1(KEYINPUT113), .C2(KEYINPUT57), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(KEYINPUT112), .B(G1956), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1018), .B1(new_n938), .B2(new_n939), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT56), .B(G2072), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n941), .A2(new_n942), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1017), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n874), .A2(new_n903), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT114), .B1(new_n878), .B2(new_n870), .ZN(new_n1025));
  AOI21_X1  g600(.A(G2067), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n879), .A2(new_n873), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n783), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n579), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1017), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1022), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(KEYINPUT117), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1017), .A2(new_n1019), .A3(new_n1034), .A4(new_n1021), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT61), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT118), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1036), .A2(KEYINPUT118), .A3(KEYINPUT61), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  XOR2_X1   g616(.A(KEYINPUT115), .B(KEYINPUT61), .Z(new_n1042));
  AND3_X1   g617(.A1(new_n1017), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1042), .B1(new_n1043), .B2(new_n1022), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT116), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1029), .ZN(new_n1046));
  NOR4_X1   g621(.A1(new_n1046), .A2(new_n1026), .A3(KEYINPUT60), .A4(new_n579), .ZN(new_n1047));
  XOR2_X1   g622(.A(KEYINPUT58), .B(G1341), .Z(new_n1048));
  NAND3_X1  g623(.A1(new_n1024), .A2(new_n1025), .A3(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1049), .B1(G1996), .B2(new_n950), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(new_n544), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT59), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT59), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1050), .A2(new_n1053), .A3(new_n544), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1047), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n1046), .A2(new_n1026), .A3(new_n588), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT60), .B1(new_n1056), .B2(new_n1030), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1058), .B(new_n1042), .C1(new_n1043), .C2(new_n1022), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1045), .A2(new_n1055), .A3(new_n1057), .A4(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1032), .B1(new_n1041), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT45), .B1(new_n813), .B2(new_n869), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n942), .A2(new_n874), .A3(new_n968), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n966), .B(new_n972), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1064));
  OR2_X1    g639(.A1(new_n1064), .A2(G171), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n975), .A2(new_n1065), .A3(new_n977), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n966), .A2(G301), .A3(new_n972), .A4(new_n969), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1067), .B1(new_n1064), .B2(G171), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1066), .A2(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1061), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1071), .A2(new_n991), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n964), .A2(new_n980), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1012), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n995), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1062), .A2(new_n874), .ZN(new_n1076));
  OR2_X1    g651(.A1(G290), .A2(G1986), .ZN(new_n1077));
  XOR2_X1   g652(.A(new_n1077), .B(KEYINPUT101), .Z(new_n1078));
  NAND2_X1  g653(.A1(G290), .A2(G1986), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1076), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  OR2_X1    g655(.A1(new_n1076), .A2(G1996), .ZN(new_n1081));
  INV_X1    g656(.A(new_n708), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  XNOR2_X1  g658(.A(new_n777), .B(G2067), .ZN(new_n1084));
  XNOR2_X1  g659(.A(new_n1076), .B(KEYINPUT102), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1083), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n671), .B(new_n674), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1085), .A2(G1996), .A3(new_n1082), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1086), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n1080), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1075), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT126), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1078), .A2(new_n1076), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n1095), .B(KEYINPUT48), .ZN(new_n1096));
  OR2_X1    g671(.A1(new_n1096), .A2(new_n1090), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n671), .A2(new_n674), .ZN(new_n1099));
  OAI22_X1  g674(.A1(new_n1098), .A2(new_n1099), .B1(G2067), .B2(new_n777), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n1085), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n1081), .B(KEYINPUT46), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1085), .A2(new_n1082), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1105), .B(KEYINPUT47), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1097), .A2(new_n1101), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1093), .A2(new_n1094), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1091), .B1(new_n995), .B2(new_n1074), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT126), .B1(new_n1110), .B2(new_n1107), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g687(.A1(new_n865), .A2(new_n866), .ZN(new_n1114));
  NOR3_X1   g688(.A1(G227), .A2(new_n459), .A3(G401), .ZN(new_n1115));
  XNOR2_X1  g689(.A(new_n1115), .B(KEYINPUT127), .ZN(new_n1116));
  NOR2_X1   g690(.A1(new_n1116), .A2(G229), .ZN(new_n1117));
  AND3_X1   g691(.A1(new_n1114), .A2(new_n823), .A3(new_n1117), .ZN(G308));
  NAND3_X1  g692(.A1(new_n1114), .A2(new_n823), .A3(new_n1117), .ZN(G225));
endmodule


