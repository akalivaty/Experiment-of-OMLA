//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 0 1 0 1 0 1 0 1 0 1 0 1 0 0 1 1 1 1 0 0 0 0 1 1 1 0 1 0 0 1 1 1 1 0 0 1 1 1 1 1 1 0 0 1 1 1 1 0 1 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n866, new_n867, new_n869, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n999, new_n1000;
  INV_X1    g000(.A(KEYINPUT29), .ZN(new_n202));
  NOR2_X1   g001(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G190gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT24), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT24), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n210), .A2(G183gat), .A3(G190gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n207), .A2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G169gat), .ZN(new_n216));
  INV_X1    g015(.A(G176gat), .ZN(new_n217));
  OAI22_X1  g016(.A1(new_n216), .A2(new_n217), .B1(KEYINPUT65), .B2(KEYINPUT23), .ZN(new_n218));
  NAND2_X1  g017(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n215), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT25), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT23), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n223), .A2(G176gat), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n222), .B1(new_n224), .B2(new_n216), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n213), .A2(new_n221), .A3(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n229), .A2(new_n223), .B1(G169gat), .B2(G176gat), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n214), .B1(new_n230), .B2(new_n219), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT64), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT64), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G169gat), .ZN(new_n234));
  AND3_X1   g033(.A1(new_n224), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n228), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(KEYINPUT64), .B(G169gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(new_n224), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n221), .A2(KEYINPUT66), .A3(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n212), .B1(G183gat), .B2(G190gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n236), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n227), .B1(new_n241), .B2(new_n222), .ZN(new_n242));
  INV_X1    g041(.A(G183gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(KEYINPUT27), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT27), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(G183gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n244), .A2(new_n246), .A3(new_n205), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT28), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT26), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n249), .A2(new_n216), .A3(new_n217), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n250), .B(new_n251), .C1(new_n216), .C2(new_n217), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n248), .A2(new_n208), .A3(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(G183gat), .ZN(new_n257));
  AND2_X1   g056(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n257), .B(KEYINPUT27), .C1(new_n258), .C2(new_n203), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n245), .B1(new_n256), .B2(new_n243), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n255), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n253), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n202), .B1(new_n242), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G226gat), .A2(G233gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT75), .ZN(new_n266));
  AND2_X1   g065(.A1(G211gat), .A2(G218gat), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n267), .A2(KEYINPUT22), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(G197gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT74), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT74), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(G197gat), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n271), .A2(new_n273), .A3(G204gat), .ZN(new_n274));
  AOI21_X1  g073(.A(G204gat), .B1(new_n271), .B2(new_n273), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n269), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g075(.A1(G211gat), .A2(G218gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n267), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(G204gat), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n272), .A2(G197gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n270), .A2(KEYINPUT74), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n271), .A2(new_n273), .A3(G204gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n278), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(new_n286), .A3(new_n269), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n279), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT75), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n263), .A2(new_n289), .A3(new_n264), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n241), .A2(new_n222), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(new_n226), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT69), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n293), .B1(new_n253), .B2(new_n261), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n259), .A2(new_n260), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(new_n254), .ZN(new_n296));
  AOI22_X1  g095(.A1(new_n247), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n296), .A2(KEYINPUT69), .A3(new_n252), .A4(new_n297), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n292), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n264), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n266), .A2(new_n288), .A3(new_n290), .A4(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT76), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n265), .A2(KEYINPUT75), .B1(new_n301), .B2(new_n300), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n306), .A2(KEYINPUT76), .A3(new_n288), .A4(new_n290), .ZN(new_n307));
  AOI211_X1 g106(.A(KEYINPUT29), .B(new_n301), .C1(new_n292), .C2(new_n299), .ZN(new_n308));
  NOR3_X1   g107(.A1(new_n242), .A2(new_n264), .A3(new_n262), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n288), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  XOR2_X1   g111(.A(G8gat), .B(G36gat), .Z(new_n313));
  XNOR2_X1  g112(.A(new_n313), .B(KEYINPUT77), .ZN(new_n314));
  XNOR2_X1  g113(.A(G64gat), .B(G92gat), .ZN(new_n315));
  XOR2_X1   g114(.A(new_n314), .B(new_n315), .Z(new_n316));
  NAND4_X1  g115(.A1(new_n305), .A2(new_n307), .A3(new_n312), .A4(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT30), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n305), .A2(new_n307), .A3(new_n312), .ZN(new_n320));
  XOR2_X1   g119(.A(new_n316), .B(KEYINPUT78), .Z(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G155gat), .B(G162gat), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(G141gat), .ZN(new_n325));
  INV_X1    g124(.A(G148gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(G141gat), .A2(G148gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n324), .B1(KEYINPUT2), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT79), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n327), .A2(KEYINPUT79), .A3(new_n328), .ZN(new_n333));
  INV_X1    g132(.A(G155gat), .ZN(new_n334));
  INV_X1    g133(.A(G162gat), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT2), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT80), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n332), .A2(new_n333), .A3(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n323), .B1(new_n336), .B2(new_n337), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n330), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT3), .ZN(new_n342));
  INV_X1    g141(.A(G113gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n343), .A2(G120gat), .ZN(new_n344));
  INV_X1    g143(.A(G120gat), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n345), .A2(G113gat), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n344), .B1(KEYINPUT70), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT70), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n348), .B1(new_n345), .B2(G113gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  XOR2_X1   g149(.A(G127gat), .B(G134gat), .Z(new_n351));
  NOR2_X1   g150(.A1(new_n351), .A2(KEYINPUT1), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT1), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n354), .B1(new_n344), .B2(new_n346), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(new_n351), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT81), .B(KEYINPUT3), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n330), .B(new_n358), .C1(new_n339), .C2(new_n340), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n342), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT4), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n361), .B1(new_n357), .B2(new_n341), .ZN(new_n362));
  INV_X1    g161(.A(new_n341), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n350), .A2(new_n352), .B1(new_n355), .B2(new_n351), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n363), .A2(KEYINPUT4), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n360), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G225gat), .A2(G233gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT5), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n364), .B(new_n330), .C1(new_n340), .C2(new_n339), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n357), .A2(new_n341), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n367), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI22_X1  g171(.A1(new_n366), .A2(new_n368), .B1(new_n369), .B2(new_n372), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n365), .A2(new_n362), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n374), .A2(KEYINPUT5), .A3(new_n367), .A4(new_n360), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G1gat), .B(G29gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(KEYINPUT0), .ZN(new_n378));
  XNOR2_X1  g177(.A(G57gat), .B(G85gat), .ZN(new_n379));
  XOR2_X1   g178(.A(new_n378), .B(new_n379), .Z(new_n380));
  NAND2_X1  g179(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n380), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n373), .A2(new_n375), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT6), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n381), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n373), .A2(new_n375), .A3(KEYINPUT6), .A4(new_n382), .ZN(new_n386));
  AND2_X1   g185(.A1(new_n386), .A2(KEYINPUT82), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n386), .A2(KEYINPUT82), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n385), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n303), .A2(new_n304), .B1(new_n311), .B2(new_n310), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n390), .A2(KEYINPUT30), .A3(new_n307), .A4(new_n316), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n319), .A2(new_n322), .A3(new_n389), .A4(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(G22gat), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n288), .B1(new_n202), .B2(new_n359), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(G228gat), .ZN(new_n396));
  INV_X1    g195(.A(G233gat), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT29), .B1(new_n279), .B2(new_n287), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n341), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n395), .A2(new_n342), .A3(new_n398), .A4(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n286), .B1(new_n285), .B2(new_n269), .ZN(new_n402));
  AOI211_X1 g201(.A(new_n278), .B(new_n268), .C1(new_n283), .C2(new_n284), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n202), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT84), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT84), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n288), .A2(new_n406), .A3(new_n202), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(new_n358), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n394), .B1(new_n408), .B2(new_n341), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n393), .B(new_n401), .C1(new_n409), .C2(new_n398), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT85), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n407), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n358), .B1(new_n399), .B2(new_n406), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n341), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n398), .B1(new_n415), .B2(new_n395), .ZN(new_n416));
  INV_X1    g215(.A(new_n401), .ZN(new_n417));
  OAI21_X1  g216(.A(G22gat), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G78gat), .B(G106gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT31), .B(G50gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n358), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n422), .B1(new_n404), .B2(KEYINPUT84), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n363), .B1(new_n423), .B2(new_n407), .ZN(new_n424));
  OAI22_X1  g223(.A1(new_n424), .A2(new_n394), .B1(new_n396), .B2(new_n397), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n425), .A2(KEYINPUT85), .A3(new_n393), .A4(new_n401), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n412), .A2(new_n418), .A3(new_n421), .A4(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n421), .B(KEYINPUT83), .ZN(new_n428));
  INV_X1    g227(.A(new_n410), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n393), .B1(new_n425), .B2(new_n401), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n292), .A2(new_n357), .A3(new_n299), .ZN(new_n433));
  NAND2_X1  g232(.A1(G227gat), .A2(G233gat), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n294), .A2(new_n298), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n364), .B1(new_n242), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n433), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT32), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT33), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  XOR2_X1   g240(.A(G15gat), .B(G43gat), .Z(new_n442));
  XNOR2_X1  g241(.A(G71gat), .B(G99gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n442), .B(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n439), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n444), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n438), .B(KEYINPUT32), .C1(new_n440), .C2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n357), .B1(new_n292), .B2(new_n299), .ZN(new_n449));
  NOR3_X1   g248(.A1(new_n242), .A2(new_n436), .A3(new_n364), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n434), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT72), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT34), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n453), .B1(new_n434), .B2(KEYINPUT71), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n433), .A2(new_n437), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT72), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(new_n456), .A3(new_n434), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n452), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n454), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n456), .B1(new_n455), .B2(new_n434), .ZN(new_n460));
  AOI211_X1 g259(.A(KEYINPUT72), .B(new_n435), .C1(new_n433), .C2(new_n437), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n448), .A2(new_n458), .A3(new_n462), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n445), .A2(new_n447), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n458), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n432), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT35), .B1(new_n392), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT73), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n464), .A2(new_n465), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n448), .B1(new_n458), .B2(new_n462), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT35), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n463), .A2(KEYINPUT73), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n472), .A2(new_n473), .A3(new_n432), .A4(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n468), .B1(new_n475), .B2(new_n392), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n392), .A2(new_n432), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n288), .B1(new_n308), .B2(new_n309), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n288), .B1(new_n306), .B2(new_n290), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n478), .B1(new_n479), .B2(KEYINPUT87), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n266), .A2(new_n290), .A3(new_n302), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT87), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n481), .A2(new_n482), .A3(new_n288), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT37), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT37), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n305), .A2(new_n307), .A3(new_n485), .A4(new_n312), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT38), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n321), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n484), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n316), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n485), .B1(new_n390), .B2(new_n307), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT38), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AND2_X1   g293(.A1(new_n373), .A2(new_n375), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT82), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n495), .A2(new_n496), .A3(KEYINPUT6), .A4(new_n382), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n386), .A2(KEYINPUT82), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT6), .B1(new_n376), .B2(new_n380), .ZN(new_n499));
  AOI22_X1  g298(.A1(new_n497), .A2(new_n498), .B1(new_n499), .B2(new_n383), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n317), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n490), .A2(new_n494), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n319), .A2(new_n391), .A3(new_n322), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n366), .A2(new_n368), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n505), .A2(KEYINPUT39), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n506), .A2(new_n382), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n370), .A2(new_n371), .A3(new_n367), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT39), .ZN(new_n509));
  OR2_X1    g308(.A1(new_n509), .A2(KEYINPUT86), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(KEYINPUT86), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n510), .A2(new_n505), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n507), .A2(KEYINPUT40), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(new_n383), .ZN(new_n514));
  AOI21_X1  g313(.A(KEYINPUT40), .B1(new_n507), .B2(new_n512), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n504), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n503), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n477), .B1(new_n518), .B2(new_n432), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT36), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n472), .A2(new_n520), .A3(new_n474), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n520), .B1(new_n466), .B2(new_n463), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n476), .B1(new_n519), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(G229gat), .A2(G233gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(G15gat), .B(G22gat), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT16), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n527), .B1(new_n528), .B2(G1gat), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n529), .B1(G1gat), .B2(new_n527), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n530), .A2(G8gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(G8gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G43gat), .B(G50gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(KEYINPUT15), .ZN(new_n535));
  INV_X1    g334(.A(G29gat), .ZN(new_n536));
  INV_X1    g335(.A(G36gat), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n536), .A2(new_n537), .A3(KEYINPUT14), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT14), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n539), .B1(G29gat), .B2(G36gat), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n538), .B(new_n540), .C1(new_n536), .C2(new_n537), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n535), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(KEYINPUT15), .A3(new_n534), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n533), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n546));
  AOI21_X1  g345(.A(KEYINPUT89), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT89), .ZN(new_n548));
  AOI211_X1 g347(.A(new_n548), .B(KEYINPUT17), .C1(new_n542), .C2(new_n543), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n533), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n542), .A2(KEYINPUT17), .A3(new_n543), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n526), .B(new_n545), .C1(new_n550), .C2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n533), .B(new_n544), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n526), .B(KEYINPUT13), .Z(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n551), .B(new_n552), .C1(new_n547), .C2(new_n549), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n560), .A2(KEYINPUT18), .A3(new_n526), .A4(new_n545), .ZN(new_n561));
  XNOR2_X1  g360(.A(G113gat), .B(G141gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G169gat), .B(G197gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n566), .B(KEYINPUT12), .Z(new_n567));
  NAND4_X1  g366(.A1(new_n556), .A2(new_n559), .A3(new_n561), .A4(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT91), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n561), .A2(new_n559), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n571), .A2(KEYINPUT91), .A3(new_n556), .A4(new_n567), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n556), .ZN(new_n574));
  INV_X1    g373(.A(new_n567), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n525), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G57gat), .B(G64gat), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(G71gat), .B(G78gat), .Z(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT21), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G231gat), .A2(G233gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(G127gat), .B(G155gat), .Z(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT20), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n587), .B(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G183gat), .B(G211gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n551), .B1(new_n584), .B2(new_n583), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT93), .ZN(new_n594));
  XOR2_X1   g393(.A(KEYINPUT92), .B(KEYINPUT19), .Z(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n592), .A2(new_n596), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(G85gat), .ZN(new_n601));
  INV_X1    g400(.A(G92gat), .ZN(new_n602));
  OAI21_X1  g401(.A(KEYINPUT94), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT94), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n604), .A2(G85gat), .A3(G92gat), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n603), .A2(KEYINPUT7), .A3(new_n605), .ZN(new_n606));
  OR2_X1    g405(.A1(G99gat), .A2(G106gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(G99gat), .A2(G106gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT7), .ZN(new_n610));
  OAI211_X1 g409(.A(KEYINPUT94), .B(new_n610), .C1(new_n601), .C2(new_n602), .ZN(new_n611));
  AOI22_X1  g410(.A1(KEYINPUT8), .A2(new_n608), .B1(new_n601), .B2(new_n602), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n606), .A2(new_n609), .A3(new_n611), .A4(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n606), .A2(new_n611), .A3(new_n612), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n614), .A2(new_n608), .A3(new_n607), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n544), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT95), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n615), .A2(new_n613), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n552), .B(new_n621), .C1(new_n547), .C2(new_n549), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(G190gat), .B(G218gat), .Z(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G134gat), .B(G162gat), .ZN(new_n626));
  AOI21_X1  g425(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n624), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n620), .A2(new_n629), .A3(new_n622), .ZN(new_n630));
  AND3_X1   g429(.A1(new_n625), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n628), .B1(new_n625), .B2(new_n630), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n621), .A2(new_n583), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT10), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n621), .A2(new_n583), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  OR3_X1    g436(.A1(new_n621), .A2(new_n583), .A3(new_n635), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(G230gat), .A2(G233gat), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n640), .B1(new_n634), .B2(new_n636), .ZN(new_n643));
  XNOR2_X1  g442(.A(G120gat), .B(G148gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(G176gat), .B(G204gat), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n644), .B(new_n645), .Z(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  OR3_X1    g446(.A1(new_n642), .A2(new_n643), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n640), .B(KEYINPUT96), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n649), .B1(new_n637), .B2(new_n638), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n647), .B1(new_n650), .B2(new_n643), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n600), .A2(new_n633), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n578), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n654), .A2(new_n389), .ZN(new_n655));
  XOR2_X1   g454(.A(KEYINPUT97), .B(G1gat), .Z(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(G1324gat));
  INV_X1    g456(.A(new_n654), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT16), .B(G8gat), .Z(new_n659));
  NAND3_X1  g458(.A1(new_n658), .A2(new_n504), .A3(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT42), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n658), .A2(new_n504), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(G8gat), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n660), .A2(new_n661), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n662), .A2(new_n664), .A3(new_n665), .ZN(G1325gat));
  AOI21_X1  g465(.A(KEYINPUT73), .B1(new_n466), .B2(new_n463), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n462), .A2(new_n458), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n469), .B1(new_n668), .B2(new_n448), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n667), .A2(KEYINPUT36), .A3(new_n669), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n670), .A2(new_n522), .A3(KEYINPUT98), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT98), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n672), .B1(new_n521), .B2(new_n523), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n674), .A2(KEYINPUT99), .ZN(new_n675));
  OAI21_X1  g474(.A(KEYINPUT98), .B1(new_n670), .B2(new_n522), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n521), .A2(new_n672), .A3(new_n523), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT99), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(G15gat), .B1(new_n654), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n472), .A2(new_n474), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n684), .A2(G15gat), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n683), .B1(new_n654), .B2(new_n685), .ZN(G1326gat));
  NOR2_X1   g485(.A1(new_n654), .A2(new_n432), .ZN(new_n687));
  XOR2_X1   g486(.A(KEYINPUT43), .B(G22gat), .Z(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1327gat));
  INV_X1    g488(.A(new_n633), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n690), .A2(new_n599), .A3(new_n652), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n578), .A2(new_n536), .A3(new_n500), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT45), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n525), .A2(new_n633), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT44), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT101), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n476), .A2(new_n696), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n468), .B(KEYINPUT101), .C1(new_n475), .C2(new_n392), .ZN(new_n698));
  OAI211_X1 g497(.A(new_n697), .B(new_n698), .C1(new_n674), .C2(new_n519), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n699), .A2(new_n700), .A3(new_n633), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n695), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n652), .B(KEYINPUT100), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n573), .A2(new_n576), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n703), .A2(new_n704), .A3(new_n599), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(G29gat), .B1(new_n706), .B2(new_n389), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n693), .A2(new_n707), .ZN(G1328gat));
  NAND4_X1  g507(.A1(new_n578), .A2(new_n537), .A3(new_n504), .A4(new_n691), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(KEYINPUT46), .Z(new_n710));
  AND2_X1   g509(.A1(new_n702), .A2(new_n705), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n504), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT102), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(G36gat), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n712), .A2(new_n713), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n710), .B1(new_n715), .B2(new_n716), .ZN(G1329gat));
  INV_X1    g516(.A(G43gat), .ZN(new_n718));
  INV_X1    g517(.A(new_n684), .ZN(new_n719));
  AND4_X1   g518(.A1(new_n718), .A2(new_n578), .A3(new_n719), .A4(new_n691), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT47), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT103), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n723), .B1(new_n706), .B2(new_n678), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(G43gat), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n706), .A2(new_n723), .A3(new_n678), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n722), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n718), .B1(new_n711), .B2(new_n681), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n721), .B1(new_n728), .B2(new_n720), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(G1330gat));
  OAI21_X1  g529(.A(G50gat), .B1(new_n706), .B2(new_n432), .ZN(new_n731));
  INV_X1    g530(.A(G50gat), .ZN(new_n732));
  INV_X1    g531(.A(new_n432), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n578), .A2(new_n732), .A3(new_n733), .A4(new_n691), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT48), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1331gat));
  NOR2_X1   g536(.A1(new_n600), .A2(new_n633), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n738), .A2(new_n704), .A3(new_n703), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT104), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n699), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n741), .A2(new_n389), .ZN(new_n742));
  XNOR2_X1  g541(.A(KEYINPUT105), .B(G57gat), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(G1332gat));
  AND2_X1   g543(.A1(new_n740), .A2(new_n699), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT49), .ZN(new_n746));
  INV_X1    g545(.A(G64gat), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n504), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  XOR2_X1   g547(.A(new_n748), .B(KEYINPUT106), .Z(new_n749));
  NAND2_X1  g548(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n746), .A2(new_n747), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1333gat));
  AND3_X1   g551(.A1(new_n745), .A2(G71gat), .A3(new_n681), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT107), .B1(new_n745), .B2(new_n719), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n754), .A2(G71gat), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n745), .A2(KEYINPUT107), .A3(new_n719), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n753), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  XOR2_X1   g556(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(G1334gat));
  NAND2_X1  g558(.A1(new_n745), .A2(new_n733), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g560(.A1(new_n600), .A2(new_n704), .ZN(new_n762));
  INV_X1    g561(.A(new_n652), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n702), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(G85gat), .B1(new_n765), .B2(new_n389), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n762), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n699), .A2(new_n633), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(KEYINPUT109), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT109), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n699), .A2(new_n771), .A3(new_n633), .A4(new_n768), .ZN(new_n772));
  INV_X1    g571(.A(new_n762), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n699), .A2(new_n633), .A3(new_n773), .ZN(new_n774));
  AOI22_X1  g573(.A1(new_n770), .A2(new_n772), .B1(new_n767), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n500), .A2(new_n652), .A3(new_n601), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT110), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n766), .B1(new_n775), .B2(new_n777), .ZN(G1336gat));
  NAND3_X1  g577(.A1(new_n703), .A2(new_n602), .A3(new_n504), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n774), .A2(new_n767), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n769), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n633), .A2(new_n700), .ZN(new_n783));
  INV_X1    g582(.A(new_n698), .ZN(new_n784));
  INV_X1    g583(.A(new_n477), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n482), .B1(new_n481), .B2(new_n288), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n479), .A2(KEYINPUT87), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n786), .A2(new_n787), .A3(new_n478), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n488), .B1(new_n788), .B2(KEYINPUT37), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n501), .B1(new_n789), .B2(new_n486), .ZN(new_n790));
  AOI22_X1  g589(.A1(new_n790), .A2(new_n494), .B1(new_n504), .B2(new_n516), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n785), .B1(new_n791), .B2(new_n733), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n784), .B1(new_n792), .B2(new_n678), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n783), .B1(new_n793), .B2(new_n697), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n700), .B1(new_n525), .B2(new_n633), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n504), .B(new_n764), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  AOI22_X1  g595(.A1(new_n780), .A2(new_n782), .B1(new_n796), .B2(G92gat), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798));
  OAI21_X1  g597(.A(KEYINPUT111), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT111), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n796), .A2(G92gat), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n779), .B1(new_n781), .B2(new_n769), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n800), .B(KEYINPUT52), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n796), .A2(G92gat), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n798), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n770), .A2(new_n772), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n779), .B1(new_n808), .B2(new_n781), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n805), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT52), .B1(new_n796), .B2(G92gat), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n811), .B(KEYINPUT112), .C1(new_n775), .C2(new_n779), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n804), .A2(new_n813), .ZN(G1337gat));
  OAI21_X1  g613(.A(G99gat), .B1(new_n765), .B2(new_n682), .ZN(new_n815));
  OR3_X1    g614(.A1(new_n684), .A2(G99gat), .A3(new_n763), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n815), .B1(new_n775), .B2(new_n816), .ZN(G1338gat));
  NAND3_X1  g616(.A1(new_n702), .A2(new_n733), .A3(new_n764), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(G106gat), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT113), .ZN(new_n820));
  INV_X1    g619(.A(new_n703), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n821), .A2(G106gat), .A3(new_n432), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n823), .B1(new_n781), .B2(new_n769), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n819), .B1(new_n820), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n824), .A2(new_n820), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT53), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n819), .B(new_n828), .C1(new_n775), .C2(new_n823), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(G1339gat));
  INV_X1    g629(.A(new_n649), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n641), .B(KEYINPUT54), .C1(new_n639), .C2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT55), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n646), .B1(new_n650), .B2(new_n834), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n832), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n833), .B1(new_n832), .B2(new_n835), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n648), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OR3_X1    g637(.A1(new_n838), .A2(new_n631), .A3(new_n632), .ZN(new_n839));
  INV_X1    g638(.A(new_n566), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n526), .B1(new_n560), .B2(new_n545), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n557), .A2(new_n558), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(KEYINPUT114), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n573), .A2(new_n844), .ZN(new_n845));
  OR2_X1    g644(.A1(new_n839), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n573), .A2(new_n844), .A3(new_n652), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n847), .B1(new_n704), .B2(new_n838), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n690), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n599), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n738), .A2(new_n704), .A3(new_n763), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n853), .A2(new_n389), .A3(new_n504), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n684), .A2(new_n733), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n856), .A2(new_n343), .A3(new_n704), .ZN(new_n857));
  INV_X1    g656(.A(new_n467), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n577), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n857), .B1(new_n343), .B2(new_n861), .ZN(G1340gat));
  NOR3_X1   g661(.A1(new_n856), .A2(new_n345), .A3(new_n821), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n860), .A2(new_n652), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n863), .B1(new_n345), .B2(new_n864), .ZN(G1341gat));
  OAI21_X1  g664(.A(G127gat), .B1(new_n856), .B2(new_n600), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n600), .A2(G127gat), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n866), .B1(new_n859), .B2(new_n867), .ZN(G1342gat));
  OR3_X1    g667(.A1(new_n859), .A2(G134gat), .A3(new_n690), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n869), .A2(KEYINPUT56), .ZN(new_n870));
  OAI21_X1  g669(.A(G134gat), .B1(new_n856), .B2(new_n690), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(KEYINPUT56), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(G1343gat));
  NOR4_X1   g672(.A1(new_n853), .A2(new_n389), .A3(new_n432), .A4(new_n504), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n682), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n325), .B1(new_n875), .B2(new_n704), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n877), .B1(new_n853), .B2(new_n432), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT115), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n839), .A2(new_n845), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n838), .A2(KEYINPUT117), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT117), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n882), .B(new_n648), .C1(new_n836), .C2(new_n837), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n881), .A2(new_n577), .A3(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT116), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n847), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n573), .A2(new_n844), .A3(KEYINPUT116), .A4(new_n652), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n884), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n880), .B1(new_n888), .B2(new_n690), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n851), .B1(new_n889), .B2(new_n599), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n432), .A2(new_n877), .ZN(new_n891));
  AOI22_X1  g690(.A1(new_n878), .A2(new_n879), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI211_X1 g691(.A(KEYINPUT115), .B(new_n877), .C1(new_n853), .C2(new_n432), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n504), .A2(new_n389), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n678), .A2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n704), .A2(new_n325), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n876), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT58), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n876), .B(KEYINPUT58), .C1(new_n898), .C2(new_n900), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(G1344gat));
  INV_X1    g704(.A(new_n875), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(new_n326), .A3(new_n652), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n896), .B1(new_n892), .B2(new_n893), .ZN(new_n908));
  AOI211_X1 g707(.A(KEYINPUT59), .B(new_n326), .C1(new_n908), .C2(new_n652), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT59), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT118), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n600), .B1(new_n889), .B2(new_n911), .ZN(new_n912));
  AOI211_X1 g711(.A(KEYINPUT118), .B(new_n880), .C1(new_n888), .C2(new_n690), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n851), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n432), .A2(KEYINPUT57), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT57), .B1(new_n853), .B2(new_n432), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n916), .A2(new_n652), .A3(new_n897), .A4(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n910), .B1(new_n918), .B2(G148gat), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n907), .B1(new_n909), .B2(new_n919), .ZN(G1345gat));
  OAI21_X1  g719(.A(G155gat), .B1(new_n898), .B2(new_n600), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n906), .A2(new_n334), .A3(new_n599), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(G1346gat));
  OAI21_X1  g722(.A(new_n335), .B1(new_n875), .B2(new_n690), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n690), .A2(new_n335), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n924), .B1(new_n898), .B2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT119), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n924), .B(KEYINPUT119), .C1(new_n898), .C2(new_n926), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1347gat));
  OR2_X1    g730(.A1(new_n850), .A2(new_n852), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n504), .A2(new_n389), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n932), .A2(new_n858), .A3(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n936), .A2(new_n237), .A3(new_n577), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT120), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n932), .A2(new_n938), .A3(new_n855), .A4(new_n934), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n855), .B(new_n934), .C1(new_n850), .C2(new_n852), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT120), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n939), .A2(new_n577), .A3(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT121), .ZN(new_n943));
  AND3_X1   g742(.A1(new_n942), .A2(new_n943), .A3(G169gat), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n943), .B1(new_n942), .B2(G169gat), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n937), .B1(new_n944), .B2(new_n945), .ZN(G1348gat));
  NAND3_X1  g745(.A1(new_n936), .A2(new_n217), .A3(new_n652), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n939), .A2(new_n703), .A3(new_n941), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n947), .B1(new_n948), .B2(new_n217), .ZN(G1349gat));
  NAND3_X1  g748(.A1(new_n599), .A2(new_n244), .A3(new_n246), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n935), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n939), .A2(new_n599), .A3(new_n941), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n258), .A2(new_n203), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n951), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT123), .ZN(new_n956));
  AND4_X1   g755(.A1(KEYINPUT122), .A2(new_n955), .A3(new_n956), .A4(KEYINPUT60), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n955), .A2(KEYINPUT122), .ZN(new_n958));
  AOI21_X1  g757(.A(KEYINPUT60), .B1(new_n955), .B2(new_n956), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(G1350gat));
  NAND3_X1  g759(.A1(new_n936), .A2(new_n205), .A3(new_n633), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n939), .A2(new_n633), .A3(new_n941), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT61), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n962), .A2(new_n963), .A3(G190gat), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n963), .B1(new_n962), .B2(G190gat), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n961), .B1(new_n964), .B2(new_n965), .ZN(G1351gat));
  NOR2_X1   g765(.A1(new_n681), .A2(new_n933), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n916), .A2(new_n917), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(G197gat), .B1(new_n968), .B2(new_n704), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n853), .A2(new_n432), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  INV_X1    g770(.A(new_n971), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n972), .A2(new_n270), .A3(new_n577), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n969), .A2(new_n973), .ZN(G1352gat));
  XNOR2_X1  g773(.A(KEYINPUT124), .B(G204gat), .ZN(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n976), .B1(new_n968), .B2(new_n821), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n972), .A2(new_n652), .A3(new_n975), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n978), .A2(KEYINPUT62), .ZN(new_n979));
  NOR3_X1   g778(.A1(new_n971), .A2(new_n763), .A3(new_n976), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT62), .ZN(new_n981));
  AND3_X1   g780(.A1(new_n980), .A2(KEYINPUT125), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g781(.A(KEYINPUT125), .B1(new_n980), .B2(new_n981), .ZN(new_n983));
  OAI211_X1 g782(.A(new_n977), .B(new_n979), .C1(new_n982), .C2(new_n983), .ZN(G1353gat));
  NAND4_X1  g783(.A1(new_n916), .A2(new_n967), .A3(new_n599), .A4(new_n917), .ZN(new_n985));
  NOR2_X1   g784(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n985), .A2(G211gat), .A3(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(G211gat), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n972), .A2(new_n988), .A3(new_n599), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  XOR2_X1   g789(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n991));
  INV_X1    g790(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n992), .B1(new_n985), .B2(G211gat), .ZN(new_n993));
  OAI21_X1  g792(.A(KEYINPUT127), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  INV_X1    g793(.A(new_n993), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT127), .ZN(new_n996));
  NAND4_X1  g795(.A1(new_n995), .A2(new_n996), .A3(new_n989), .A4(new_n987), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n994), .A2(new_n997), .ZN(G1354gat));
  OAI21_X1  g797(.A(G218gat), .B1(new_n968), .B2(new_n690), .ZN(new_n999));
  OR2_X1    g798(.A1(new_n690), .A2(G218gat), .ZN(new_n1000));
  OAI21_X1  g799(.A(new_n999), .B1(new_n971), .B2(new_n1000), .ZN(G1355gat));
endmodule


