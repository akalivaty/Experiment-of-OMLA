//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n803, new_n804, new_n805, new_n807,
    new_n808, new_n809, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n866, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n202));
  OR3_X1    g001(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n203));
  OAI21_X1  g002(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT24), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n212));
  NOR3_X1   g011(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT25), .B1(new_n207), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT25), .ZN(new_n215));
  AOI22_X1  g014(.A1(new_n203), .A2(new_n204), .B1(G169gat), .B2(G176gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n212), .B(KEYINPUT64), .ZN(new_n217));
  OR2_X1    g016(.A1(new_n210), .A2(new_n211), .ZN(new_n218));
  OAI211_X1 g017(.A(new_n215), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(new_n206), .ZN(new_n222));
  NOR3_X1   g021(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n208), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n224), .A2(KEYINPUT65), .ZN(new_n225));
  XOR2_X1   g024(.A(KEYINPUT27), .B(G183gat), .Z(new_n226));
  OR3_X1    g025(.A1(new_n226), .A2(KEYINPUT28), .A3(G190gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n224), .A2(KEYINPUT65), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT28), .B1(new_n226), .B2(G190gat), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n225), .A2(new_n227), .A3(new_n228), .A4(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n220), .A2(new_n230), .ZN(new_n231));
  AND3_X1   g030(.A1(new_n231), .A2(G226gat), .A3(G233gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT69), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT29), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n231), .A2(new_n234), .B1(G226gat), .B2(G233gat), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n231), .A2(G226gat), .A3(G233gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT69), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT67), .B(G197gat), .ZN(new_n240));
  INV_X1    g039(.A(G204gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT22), .ZN(new_n243));
  INV_X1    g042(.A(G211gat), .ZN(new_n244));
  INV_X1    g043(.A(G218gat), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n242), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G211gat), .B(G218gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n242), .A2(new_n250), .A3(new_n246), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n233), .A2(new_n236), .A3(new_n239), .A4(new_n254), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n253), .B(new_n252), .C1(new_n235), .C2(new_n232), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  XOR2_X1   g056(.A(G64gat), .B(G92gat), .Z(new_n258));
  XNOR2_X1  g057(.A(G8gat), .B(G36gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n261));
  XOR2_X1   g060(.A(new_n260), .B(new_n261), .Z(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT30), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n202), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n262), .B1(new_n255), .B2(new_n256), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n267), .A2(KEYINPUT72), .A3(KEYINPUT30), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n264), .A2(new_n265), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n255), .A2(new_n256), .A3(new_n262), .ZN(new_n271));
  AND3_X1   g070(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n273));
  XNOR2_X1  g072(.A(G1gat), .B(G29gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G57gat), .B(G85gat), .ZN(new_n276));
  XOR2_X1   g075(.A(new_n275), .B(new_n276), .Z(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT75), .ZN(new_n279));
  XOR2_X1   g078(.A(G127gat), .B(G134gat), .Z(new_n280));
  INV_X1    g079(.A(KEYINPUT66), .ZN(new_n281));
  XOR2_X1   g080(.A(G113gat), .B(G120gat), .Z(new_n282));
  AOI21_X1  g081(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT1), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n284), .B(new_n282), .C1(new_n280), .C2(new_n281), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G155gat), .A2(G162gat), .ZN(new_n289));
  OR2_X1    g088(.A1(G155gat), .A2(G162gat), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n289), .B1(new_n290), .B2(KEYINPUT2), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT73), .ZN(new_n292));
  INV_X1    g091(.A(G141gat), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n292), .B1(new_n293), .B2(G148gat), .ZN(new_n294));
  INV_X1    g093(.A(G148gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n295), .A2(KEYINPUT73), .A3(G141gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n295), .A2(G141gat), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n291), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G141gat), .B(G148gat), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n289), .B(new_n290), .C1(new_n300), .C2(KEYINPUT2), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n288), .B(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(G225gat), .A2(G233gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT5), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n279), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n304), .ZN(new_n308));
  INV_X1    g107(.A(new_n288), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n309), .A2(new_n302), .ZN(new_n310));
  INV_X1    g109(.A(new_n302), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n288), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n308), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n313), .A2(KEYINPUT75), .A3(KEYINPUT5), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n302), .B(KEYINPUT74), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n315), .A2(KEYINPUT4), .A3(new_n288), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT4), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n317), .B1(new_n309), .B2(new_n302), .ZN(new_n318));
  AND3_X1   g117(.A1(new_n316), .A2(new_n304), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT3), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n311), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n302), .A2(KEYINPUT3), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n309), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n307), .A2(new_n314), .B1(new_n319), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n315), .A2(new_n317), .A3(new_n288), .ZN(new_n325));
  OR2_X1    g124(.A1(new_n325), .A2(KEYINPUT77), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n325), .B(KEYINPUT77), .C1(new_n317), .C2(new_n310), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n308), .A2(KEYINPUT5), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n326), .A2(new_n327), .A3(new_n323), .A4(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n278), .B1(new_n324), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n319), .A2(new_n323), .ZN(new_n332));
  INV_X1    g131(.A(new_n314), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT75), .B1(new_n313), .B2(KEYINPUT5), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n335), .A2(new_n277), .A3(new_n329), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT6), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n331), .A2(new_n336), .A3(KEYINPUT78), .A4(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT78), .ZN(new_n339));
  OAI221_X1 g138(.A(new_n278), .B1(new_n339), .B2(KEYINPUT6), .C1(new_n324), .C2(new_n330), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n272), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(G22gat), .B(G50gat), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(G228gat), .ZN(new_n346));
  INV_X1    g145(.A(G233gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n252), .A2(KEYINPUT79), .A3(new_n234), .A4(new_n253), .ZN(new_n349));
  AND2_X1   g148(.A1(new_n349), .A2(new_n320), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n252), .A2(new_n234), .A3(new_n253), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n311), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n321), .A2(new_n234), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(new_n254), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n348), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT31), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n315), .B1(new_n351), .B2(new_n320), .ZN(new_n360));
  INV_X1    g159(.A(new_n348), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n356), .A2(new_n361), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n358), .B(new_n359), .C1(new_n360), .C2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n353), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n320), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n302), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n361), .B1(new_n366), .B2(new_n356), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n362), .A2(new_n360), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT31), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  XOR2_X1   g168(.A(G78gat), .B(G106gat), .Z(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n363), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n371), .B1(new_n363), .B2(new_n369), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n345), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n363), .A2(new_n369), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n370), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n377), .A2(new_n344), .A3(new_n372), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n375), .A2(new_n378), .A3(KEYINPUT80), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT80), .B1(new_n375), .B2(new_n378), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n343), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n303), .A2(new_n304), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT39), .ZN(new_n384));
  XOR2_X1   g183(.A(new_n384), .B(KEYINPUT81), .Z(new_n385));
  NAND3_X1  g184(.A1(new_n326), .A2(new_n327), .A3(new_n323), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(new_n308), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  OR2_X1    g187(.A1(new_n387), .A2(KEYINPUT39), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n388), .A2(new_n277), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT40), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n388), .A2(KEYINPUT40), .A3(new_n277), .A4(new_n389), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n382), .A2(new_n392), .A3(new_n331), .A4(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT37), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n263), .B1(new_n257), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n396), .B1(new_n395), .B2(new_n257), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n267), .B1(new_n397), .B2(KEYINPUT38), .ZN(new_n398));
  OAI211_X1 g197(.A(KEYINPUT6), .B(new_n278), .C1(new_n324), .C2(new_n330), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n331), .A2(new_n336), .A3(new_n337), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT38), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n236), .A2(new_n237), .A3(new_n254), .ZN(new_n402));
  AND3_X1   g201(.A1(new_n233), .A2(new_n236), .A3(new_n239), .ZN(new_n403));
  OAI211_X1 g202(.A(KEYINPUT37), .B(new_n402), .C1(new_n403), .C2(new_n254), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n396), .A2(new_n401), .A3(new_n404), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n398), .A2(new_n399), .A3(new_n400), .A4(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n375), .A2(new_n378), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n394), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n381), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G15gat), .B(G43gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(G71gat), .ZN(new_n411));
  INV_X1    g210(.A(G99gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n231), .A2(new_n288), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n309), .A2(new_n220), .A3(new_n230), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(G227gat), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n416), .A2(new_n417), .A3(new_n347), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n413), .B1(new_n418), .B2(KEYINPUT33), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT32), .ZN(new_n420));
  NOR3_X1   g219(.A1(new_n418), .A2(new_n420), .A3(KEYINPUT34), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT34), .ZN(new_n422));
  AND2_X1   g221(.A1(new_n414), .A2(new_n415), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n417), .A2(new_n347), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n422), .B1(new_n425), .B2(KEYINPUT32), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n423), .A2(new_n424), .ZN(new_n427));
  NOR3_X1   g226(.A1(new_n421), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n427), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT34), .B1(new_n418), .B2(new_n420), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n425), .A2(KEYINPUT32), .A3(new_n422), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n419), .B1(new_n428), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n427), .B1(new_n421), .B2(new_n426), .ZN(new_n434));
  INV_X1    g233(.A(new_n419), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n430), .A2(new_n431), .A3(new_n429), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n433), .A2(KEYINPUT36), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT36), .ZN(new_n439));
  NOR3_X1   g238(.A1(new_n428), .A2(new_n432), .A3(new_n419), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n435), .B1(new_n434), .B2(new_n436), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n409), .B1(new_n438), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT35), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n343), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n407), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n440), .A2(new_n441), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n400), .A2(new_n399), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n407), .A2(new_n272), .A3(new_n451), .A4(new_n447), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n444), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  OR2_X1    g253(.A1(new_n443), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(G57gat), .B(G64gat), .ZN(new_n456));
  OR2_X1    g255(.A1(new_n456), .A2(KEYINPUT87), .ZN(new_n457));
  AND2_X1   g256(.A1(G71gat), .A2(G78gat), .ZN(new_n458));
  OR2_X1    g257(.A1(new_n458), .A2(KEYINPUT9), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n456), .A2(KEYINPUT87), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n457), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(G71gat), .B(G78gat), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n459), .A2(new_n462), .ZN(new_n465));
  INV_X1    g264(.A(G64gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(G57gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(KEYINPUT88), .B(G57gat), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n467), .B1(new_n468), .B2(new_n466), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n464), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT21), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(G15gat), .B(G22gat), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT16), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n474), .B1(new_n475), .B2(G1gat), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n476), .B1(G1gat), .B2(new_n474), .ZN(new_n477));
  INV_X1    g276(.A(G8gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n477), .B(new_n478), .ZN(new_n479));
  OR2_X1    g278(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n471), .A2(new_n472), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n473), .A2(new_n479), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  XOR2_X1   g282(.A(KEYINPUT90), .B(KEYINPUT19), .Z(new_n484));
  XNOR2_X1  g283(.A(new_n483), .B(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G127gat), .B(G155gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n485), .B(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(G183gat), .B(G211gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(KEYINPUT91), .ZN(new_n489));
  NAND2_X1  g288(.A1(G231gat), .A2(G233gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n489), .B(new_n490), .ZN(new_n491));
  XOR2_X1   g290(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n492));
  XOR2_X1   g291(.A(new_n491), .B(new_n492), .Z(new_n493));
  XNOR2_X1  g292(.A(new_n487), .B(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT15), .ZN(new_n495));
  INV_X1    g294(.A(G50gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(G43gat), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT83), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n497), .B(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(G43gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(G50gat), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT84), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n495), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n501), .A2(new_n497), .A3(KEYINPUT15), .ZN(new_n505));
  NOR2_X1   g304(.A1(G29gat), .A2(G36gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(KEYINPUT14), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(G29gat), .A2(G36gat), .ZN(new_n509));
  XOR2_X1   g308(.A(new_n509), .B(KEYINPUT85), .Z(new_n510));
  NAND4_X1  g309(.A1(new_n504), .A2(new_n505), .A3(new_n508), .A4(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n505), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n508), .A2(KEYINPUT82), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT82), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n509), .B1(new_n507), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n512), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n517), .B(KEYINPUT17), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT94), .ZN(new_n519));
  XOR2_X1   g318(.A(G99gat), .B(G106gat), .Z(new_n520));
  NAND2_X1  g319(.A1(G99gat), .A2(G106gat), .ZN(new_n521));
  INV_X1    g320(.A(G85gat), .ZN(new_n522));
  INV_X1    g321(.A(G92gat), .ZN(new_n523));
  AOI22_X1  g322(.A1(KEYINPUT8), .A2(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT92), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n528));
  AND2_X1   g327(.A1(G85gat), .A2(G92gat), .ZN(new_n529));
  AND3_X1   g328(.A1(new_n528), .A2(new_n529), .A3(KEYINPUT93), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT93), .B1(new_n528), .B2(new_n529), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n527), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT93), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT7), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n534), .A2(KEYINPUT92), .ZN(new_n535));
  NAND2_X1  g334(.A1(G85gat), .A2(G92gat), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n533), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n527), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n528), .A2(new_n529), .A3(KEYINPUT93), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AOI211_X1 g339(.A(new_n520), .B(new_n525), .C1(new_n532), .C2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n520), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n532), .A2(new_n540), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n542), .B1(new_n543), .B2(new_n524), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n518), .B(new_n519), .C1(new_n541), .C2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n546));
  INV_X1    g345(.A(new_n517), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n547), .B1(new_n519), .B2(KEYINPUT17), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n543), .A2(new_n542), .A3(new_n524), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n538), .B1(new_n537), .B2(new_n539), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n524), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n520), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n548), .A2(new_n549), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n545), .A2(new_n546), .A3(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G134gat), .B(G162gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(G190gat), .B(G218gat), .Z(new_n558));
  AOI21_X1  g357(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n557), .B(new_n560), .Z(new_n561));
  AND3_X1   g360(.A1(new_n455), .A2(new_n494), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G230gat), .A2(G233gat), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n471), .B1(new_n544), .B2(new_n541), .ZN(new_n565));
  AOI22_X1  g364(.A1(new_n461), .A2(new_n463), .B1(new_n469), .B2(new_n465), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n553), .A2(new_n549), .A3(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT10), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n565), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n553), .A2(new_n549), .A3(KEYINPUT10), .A4(new_n566), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n564), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n563), .B1(new_n565), .B2(new_n567), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G120gat), .B(G148gat), .ZN(new_n574));
  INV_X1    g373(.A(G176gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(new_n241), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n579), .A2(KEYINPUT95), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(KEYINPUT95), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT96), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n569), .A2(new_n570), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n583), .B1(new_n584), .B2(new_n563), .ZN(new_n585));
  AOI211_X1 g384(.A(KEYINPUT96), .B(new_n564), .C1(new_n569), .C2(new_n570), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n572), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n578), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n582), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n518), .A2(new_n479), .ZN(new_n592));
  NAND2_X1  g391(.A1(G229gat), .A2(G233gat), .ZN(new_n593));
  OR2_X1    g392(.A1(new_n547), .A2(new_n479), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT18), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT86), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n592), .A2(KEYINPUT18), .A3(new_n593), .A4(new_n594), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n517), .B(new_n479), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n593), .B(KEYINPUT13), .ZN(new_n601));
  OR2_X1    g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G113gat), .B(G141gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(G197gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT11), .ZN(new_n606));
  INV_X1    g405(.A(G169gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n608), .B(KEYINPUT12), .Z(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT86), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n595), .A2(new_n611), .A3(new_n596), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n598), .A2(new_n603), .A3(new_n610), .A4(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n597), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n602), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n609), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n591), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n562), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n620), .A2(new_n342), .ZN(new_n621));
  XOR2_X1   g420(.A(KEYINPUT97), .B(G1gat), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(G1324gat));
  INV_X1    g422(.A(new_n620), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n478), .B1(new_n624), .B2(new_n382), .ZN(new_n625));
  NOR2_X1   g424(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n475), .A2(new_n478), .ZN(new_n627));
  NOR4_X1   g426(.A1(new_n620), .A2(new_n272), .A3(new_n626), .A4(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(KEYINPUT42), .B1(new_n625), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n629), .B1(KEYINPUT42), .B2(new_n628), .ZN(G1325gat));
  NOR3_X1   g429(.A1(new_n440), .A2(new_n441), .A3(new_n439), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT36), .B1(new_n433), .B2(new_n437), .ZN(new_n632));
  OAI21_X1  g431(.A(KEYINPUT98), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT98), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n442), .A2(new_n634), .A3(new_n438), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n624), .A2(G15gat), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(G15gat), .B1(new_n624), .B2(new_n447), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(G1326gat));
  NOR2_X1   g439(.A1(new_n379), .A2(new_n380), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n620), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(KEYINPUT43), .B(G22gat), .Z(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(G1327gat));
  XNOR2_X1  g443(.A(new_n557), .B(new_n560), .ZN(new_n645));
  AND2_X1   g444(.A1(new_n455), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n493), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n487), .B(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n646), .A2(new_n619), .A3(new_n648), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n649), .A2(G29gat), .A3(new_n342), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n650), .B(KEYINPUT45), .Z(new_n651));
  INV_X1    g450(.A(KEYINPUT44), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n381), .A2(new_n636), .A3(new_n408), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT101), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n381), .A2(new_n636), .A3(KEYINPUT101), .A4(new_n408), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n454), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n652), .B1(new_n657), .B2(new_n561), .ZN(new_n658));
  OAI211_X1 g457(.A(KEYINPUT44), .B(new_n645), .C1(new_n443), .C2(new_n454), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n494), .B(KEYINPUT99), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(new_n619), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n664), .B(KEYINPUT100), .Z(new_n665));
  NAND3_X1  g464(.A1(new_n661), .A2(new_n341), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(G29gat), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n667), .ZN(G1328gat));
  OR3_X1    g467(.A1(new_n649), .A2(G36gat), .A3(new_n272), .ZN(new_n669));
  OR2_X1    g468(.A1(new_n669), .A2(KEYINPUT46), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n661), .A2(new_n382), .A3(new_n665), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n671), .A2(KEYINPUT102), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(KEYINPUT102), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n672), .A2(G36gat), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n669), .A2(KEYINPUT46), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n670), .A2(new_n674), .A3(new_n675), .ZN(G1329gat));
  OAI21_X1  g475(.A(new_n500), .B1(new_n649), .B2(new_n448), .ZN(new_n677));
  NAND2_X1  g476(.A1(KEYINPUT103), .A2(KEYINPUT47), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n661), .A2(G43gat), .A3(new_n637), .A4(new_n665), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(KEYINPUT103), .A2(KEYINPUT47), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n680), .B(new_n681), .Z(G1330gat));
  OR3_X1    g481(.A1(new_n649), .A2(G50gat), .A3(new_n641), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n661), .A2(new_n446), .A3(new_n665), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n683), .B(KEYINPUT48), .C1(new_n496), .C2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n641), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n661), .A2(new_n686), .A3(new_n665), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(G50gat), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n685), .B1(new_n689), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g489(.A1(new_n561), .A2(new_n618), .A3(new_n494), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n657), .A2(new_n590), .A3(new_n691), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n341), .B(KEYINPUT104), .Z(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT105), .Z(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(new_n468), .ZN(G1332gat));
  INV_X1    g496(.A(KEYINPUT49), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n692), .B1(new_n698), .B2(new_n466), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(new_n272), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT106), .ZN(new_n701));
  NOR2_X1   g500(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1333gat));
  NAND3_X1  g502(.A1(new_n692), .A2(G71gat), .A3(new_n637), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n692), .A2(new_n447), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n704), .B1(new_n705), .B2(G71gat), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n686), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT107), .B(G78gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1335gat));
  NAND2_X1  g509(.A1(new_n655), .A2(new_n656), .ZN(new_n711));
  INV_X1    g510(.A(new_n454), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n494), .A2(new_n617), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n713), .A2(new_n645), .A3(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT51), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n713), .A2(KEYINPUT51), .A3(new_n645), .A4(new_n714), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n719), .A2(new_n590), .ZN(new_n720));
  AOI21_X1  g519(.A(G85gat), .B1(new_n720), .B2(new_n341), .ZN(new_n721));
  INV_X1    g520(.A(new_n714), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n660), .A2(new_n590), .A3(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n342), .A2(new_n522), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n721), .B1(new_n723), .B2(new_n724), .ZN(G1336gat));
  AND2_X1   g524(.A1(new_n723), .A2(new_n382), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n591), .A2(new_n382), .A3(new_n523), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT108), .ZN(new_n728));
  OAI22_X1  g527(.A1(new_n726), .A2(new_n523), .B1(new_n719), .B2(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT52), .ZN(G1337gat));
  AOI21_X1  g529(.A(G99gat), .B1(new_n720), .B2(new_n447), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n636), .A2(new_n412), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n731), .B1(new_n723), .B2(new_n732), .ZN(G1338gat));
  INV_X1    g532(.A(KEYINPUT53), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n722), .A2(new_n590), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n658), .A2(new_n686), .A3(new_n659), .A4(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT109), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n736), .A2(new_n737), .A3(G106gat), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n737), .B1(new_n736), .B2(G106gat), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n717), .A2(new_n718), .ZN(new_n741));
  INV_X1    g540(.A(G106gat), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n741), .A2(new_n742), .A3(new_n591), .A4(new_n446), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n734), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n658), .A2(new_n446), .A3(new_n659), .A4(new_n735), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G106gat), .ZN(new_n746));
  XOR2_X1   g545(.A(KEYINPUT110), .B(KEYINPUT53), .Z(new_n747));
  NAND3_X1  g546(.A1(new_n743), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(KEYINPUT111), .B1(new_n744), .B2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n739), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n736), .A2(new_n737), .A3(G106gat), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n743), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT53), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT111), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n754), .A2(new_n755), .A3(new_n748), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n750), .A2(new_n756), .ZN(G1339gat));
  NAND2_X1  g556(.A1(new_n584), .A2(new_n563), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n569), .A2(new_n564), .A3(new_n570), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n758), .A2(KEYINPUT54), .A3(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT54), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n585), .B2(new_n586), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT112), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n762), .A2(new_n763), .A3(new_n577), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n763), .B1(new_n762), .B2(new_n577), .ZN(new_n765));
  OAI211_X1 g564(.A(KEYINPUT55), .B(new_n760), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n582), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n561), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n615), .B1(KEYINPUT86), .B2(new_n597), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n612), .A2(new_n610), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n600), .A2(new_n601), .ZN(new_n772));
  OR2_X1    g571(.A1(new_n772), .A2(KEYINPUT113), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(KEYINPUT113), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n592), .A2(new_n594), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n773), .B(new_n774), .C1(new_n775), .C2(new_n593), .ZN(new_n776));
  AOI22_X1  g575(.A1(new_n770), .A2(new_n771), .B1(new_n608), .B2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n760), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n758), .A2(KEYINPUT96), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n571), .A2(new_n583), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT54), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT112), .B1(new_n781), .B2(new_n578), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n762), .A2(new_n763), .A3(new_n577), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n778), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n769), .B(new_n777), .C1(KEYINPUT55), .C2(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n777), .B1(new_n582), .B2(new_n589), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n617), .B1(new_n784), .B2(KEYINPUT55), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n787), .B2(new_n768), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n561), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n662), .B1(new_n785), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n691), .A2(new_n591), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n792), .A2(new_n272), .A3(new_n694), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n793), .A2(new_n446), .A3(new_n448), .ZN(new_n794));
  INV_X1    g593(.A(G113gat), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n794), .A2(new_n795), .A3(new_n617), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n790), .A2(new_n791), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n797), .A2(new_n686), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n342), .A2(new_n382), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n798), .A2(new_n447), .A3(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(G113gat), .B1(new_n800), .B2(new_n618), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n796), .A2(new_n801), .ZN(G1340gat));
  INV_X1    g601(.A(G120gat), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n794), .A2(new_n803), .A3(new_n591), .ZN(new_n804));
  OAI21_X1  g603(.A(G120gat), .B1(new_n800), .B2(new_n590), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(G1341gat));
  INV_X1    g605(.A(G127gat), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n800), .A2(new_n807), .A3(new_n663), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n794), .A2(new_n494), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n808), .B1(new_n809), .B2(new_n807), .ZN(G1342gat));
  INV_X1    g609(.A(G134gat), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n794), .A2(new_n811), .A3(new_n645), .ZN(new_n812));
  XOR2_X1   g611(.A(new_n812), .B(KEYINPUT56), .Z(new_n813));
  OAI21_X1  g612(.A(G134gat), .B1(new_n800), .B2(new_n561), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(G1343gat));
  INV_X1    g614(.A(KEYINPUT58), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n793), .A2(new_n407), .A3(new_n637), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(new_n293), .A3(new_n617), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n636), .A2(new_n799), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n792), .A2(new_n446), .ZN(new_n821));
  XNOR2_X1  g620(.A(KEYINPUT114), .B(KEYINPUT57), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n820), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  AOI211_X1 g623(.A(KEYINPUT115), .B(new_n822), .C1(new_n792), .C2(new_n446), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT116), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n788), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g627(.A(KEYINPUT116), .B(new_n786), .C1(new_n787), .C2(new_n768), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n828), .A2(new_n561), .A3(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n831));
  OR2_X1    g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n832), .A2(new_n785), .A3(new_n833), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n834), .A2(new_n648), .ZN(new_n835));
  OAI211_X1 g634(.A(KEYINPUT57), .B(new_n686), .C1(new_n835), .C2(new_n791), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n819), .B1(new_n826), .B2(new_n836), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n837), .A2(new_n617), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n816), .B(new_n818), .C1(new_n838), .C2(new_n293), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n293), .B1(new_n837), .B2(new_n617), .ZN(new_n840));
  INV_X1    g639(.A(new_n818), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT58), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n839), .A2(new_n842), .ZN(G1344gat));
  NAND3_X1  g642(.A1(new_n817), .A2(new_n295), .A3(new_n591), .ZN(new_n844));
  AOI211_X1 g643(.A(KEYINPUT59), .B(new_n295), .C1(new_n837), .C2(new_n591), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n847), .B1(new_n691), .B2(new_n591), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n648), .A2(new_n645), .A3(new_n617), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n849), .A2(KEYINPUT118), .A3(new_n590), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n830), .A2(new_n785), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n851), .B1(new_n852), .B2(new_n648), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n641), .B1(new_n853), .B2(KEYINPUT119), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n494), .B1(new_n830), .B2(new_n785), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n855), .B1(new_n856), .B2(new_n851), .ZN(new_n857));
  AOI21_X1  g656(.A(KEYINPUT57), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n821), .A2(new_n823), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OR3_X1    g659(.A1(new_n860), .A2(new_n590), .A3(new_n819), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n846), .B1(new_n861), .B2(G148gat), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n844), .B1(new_n845), .B2(new_n862), .ZN(G1345gat));
  AOI21_X1  g662(.A(G155gat), .B1(new_n817), .B2(new_n494), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n662), .A2(G155gat), .ZN(new_n865));
  XOR2_X1   g664(.A(new_n865), .B(KEYINPUT120), .Z(new_n866));
  AOI21_X1  g665(.A(new_n864), .B1(new_n837), .B2(new_n866), .ZN(G1346gat));
  AOI21_X1  g666(.A(G162gat), .B1(new_n817), .B2(new_n645), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n645), .A2(G162gat), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n868), .B1(new_n837), .B2(new_n869), .ZN(G1347gat));
  NOR2_X1   g669(.A1(new_n797), .A2(new_n341), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(new_n382), .A3(new_n449), .ZN(new_n872));
  XOR2_X1   g671(.A(new_n872), .B(KEYINPUT121), .Z(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(new_n607), .A3(new_n617), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n694), .A2(new_n272), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n447), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(KEYINPUT122), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n876), .A2(KEYINPUT122), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n798), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(G169gat), .B1(new_n879), .B2(new_n618), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n874), .A2(new_n880), .ZN(G1348gat));
  NOR3_X1   g680(.A1(new_n879), .A2(new_n575), .A3(new_n590), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n873), .A2(new_n591), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n882), .B1(new_n883), .B2(new_n575), .ZN(G1349gat));
  OAI21_X1  g683(.A(G183gat), .B1(new_n879), .B2(new_n663), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n872), .A2(new_n226), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n885), .B1(new_n886), .B2(new_n648), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT60), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n888), .A2(KEYINPUT123), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n887), .B(new_n889), .ZN(G1350gat));
  INV_X1    g689(.A(G190gat), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n873), .A2(new_n891), .A3(new_n645), .ZN(new_n892));
  OAI21_X1  g691(.A(G190gat), .B1(new_n879), .B2(new_n561), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT61), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n894), .ZN(G1351gat));
  AND4_X1   g694(.A1(new_n382), .A2(new_n871), .A3(new_n446), .A4(new_n636), .ZN(new_n896));
  XOR2_X1   g695(.A(KEYINPUT124), .B(G197gat), .Z(new_n897));
  NAND3_X1  g696(.A1(new_n896), .A2(new_n617), .A3(new_n897), .ZN(new_n898));
  XOR2_X1   g697(.A(new_n898), .B(KEYINPUT125), .Z(new_n899));
  NAND2_X1  g698(.A1(new_n875), .A2(new_n636), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n860), .A2(new_n618), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n899), .B1(new_n901), .B2(new_n897), .ZN(G1352gat));
  INV_X1    g701(.A(KEYINPUT126), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n860), .A2(new_n590), .A3(new_n900), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n904), .A2(new_n241), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n896), .A2(new_n241), .A3(new_n591), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT62), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n903), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n906), .B(new_n909), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n910), .B(KEYINPUT126), .C1(new_n241), .C2(new_n904), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n908), .A2(new_n911), .ZN(G1353gat));
  NAND3_X1  g711(.A1(new_n896), .A2(new_n244), .A3(new_n494), .ZN(new_n913));
  INV_X1    g712(.A(new_n900), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n494), .B(new_n914), .C1(new_n858), .C2(new_n859), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n915), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n916));
  AOI21_X1  g715(.A(KEYINPUT63), .B1(new_n915), .B2(G211gat), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT127), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI211_X1 g719(.A(KEYINPUT127), .B(new_n913), .C1(new_n916), .C2(new_n917), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1354gat));
  AOI21_X1  g721(.A(G218gat), .B1(new_n896), .B2(new_n645), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n860), .A2(new_n900), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n561), .A2(new_n245), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(G1355gat));
endmodule


