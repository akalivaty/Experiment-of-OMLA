//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n868, new_n869, new_n870,
    new_n872, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976, new_n977;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  AND2_X1   g004(.A1(G227gat), .A2(G233gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  AND2_X1   g006(.A1(KEYINPUT70), .A2(G127gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(KEYINPUT70), .A2(G127gat), .ZN(new_n209));
  OAI21_X1  g008(.A(G134gat), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G134gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G127gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT69), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n211), .A2(KEYINPUT69), .A3(G127gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n210), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  XOR2_X1   g015(.A(G113gat), .B(G120gat), .Z(new_n217));
  INV_X1    g016(.A(KEYINPUT1), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n211), .A2(G127gat), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n217), .A2(new_n218), .A3(new_n212), .A4(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(KEYINPUT23), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT23), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n228), .A2(KEYINPUT65), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n225), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT25), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n232), .B1(new_n224), .B2(KEYINPUT23), .ZN(new_n233));
  AND3_X1   g032(.A1(new_n230), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n235));
  OAI22_X1  g034(.A1(new_n235), .A2(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(KEYINPUT67), .A2(G183gat), .A3(G190gat), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT67), .B1(G183gat), .B2(G190gat), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n236), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G183gat), .A2(G190gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  OR2_X1    g042(.A1(G183gat), .A2(G190gat), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT24), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT66), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n243), .A2(new_n244), .A3(new_n246), .A4(new_n237), .ZN(new_n247));
  AND2_X1   g046(.A1(new_n240), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G176gat), .ZN(new_n249));
  AND2_X1   g048(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n250));
  NOR2_X1   g049(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n251));
  OAI211_X1 g050(.A(KEYINPUT23), .B(new_n249), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n241), .A2(new_n245), .ZN(new_n253));
  NAND3_X1  g052(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n244), .A3(new_n254), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n230), .A2(new_n252), .A3(new_n255), .A4(new_n231), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n234), .A2(new_n248), .B1(new_n256), .B2(new_n232), .ZN(new_n257));
  INV_X1    g056(.A(G190gat), .ZN(new_n258));
  AND2_X1   g057(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT28), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT28), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n263), .B(new_n258), .C1(new_n259), .C2(new_n260), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT26), .ZN(new_n266));
  INV_X1    g065(.A(G169gat), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n266), .A2(new_n267), .A3(new_n249), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n268), .A2(new_n231), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(new_n241), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT68), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n270), .A2(new_n273), .A3(new_n241), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n265), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n223), .B1(new_n257), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n256), .A2(new_n232), .ZN(new_n277));
  INV_X1    g076(.A(new_n231), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n228), .A2(KEYINPUT65), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n226), .A2(KEYINPUT23), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n278), .B1(new_n281), .B2(new_n225), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n282), .A2(new_n233), .A3(new_n247), .A4(new_n240), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n277), .A2(new_n283), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n270), .A2(new_n273), .A3(new_n241), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n273), .B1(new_n270), .B2(new_n241), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n262), .B(new_n264), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n217), .A2(new_n218), .A3(new_n221), .ZN(new_n288));
  AOI22_X1  g087(.A1(new_n288), .A2(new_n212), .B1(new_n216), .B2(new_n219), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n284), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n207), .B1(new_n276), .B2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT71), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT33), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n205), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n291), .A2(KEYINPUT71), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n296));
  AOI211_X1 g095(.A(new_n296), .B(new_n207), .C1(new_n276), .C2(new_n290), .ZN(new_n297));
  OAI21_X1  g096(.A(KEYINPUT32), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n276), .A2(new_n207), .A3(new_n290), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT34), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n299), .B(KEYINPUT34), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n292), .A2(KEYINPUT32), .A3(new_n303), .ZN(new_n304));
  AND3_X1   g103(.A1(new_n294), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n292), .A2(new_n293), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n304), .A2(new_n302), .B1(new_n306), .B2(new_n204), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n308), .B(KEYINPUT36), .ZN(new_n309));
  NAND2_X1  g108(.A1(G225gat), .A2(G233gat), .ZN(new_n310));
  XOR2_X1   g109(.A(G141gat), .B(G148gat), .Z(new_n311));
  OR2_X1    g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(G155gat), .A2(G162gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(KEYINPUT2), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n311), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G141gat), .B(G148gat), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n313), .B(new_n312), .C1(new_n317), .C2(KEYINPUT2), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT3), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT3), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n316), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n320), .A2(new_n223), .A3(new_n322), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n220), .A2(new_n316), .A3(new_n318), .A4(new_n222), .ZN(new_n324));
  OAI21_X1  g123(.A(KEYINPUT77), .B1(new_n324), .B2(KEYINPUT4), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT77), .ZN(new_n326));
  INV_X1    g125(.A(new_n319), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT4), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n289), .A2(new_n326), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n316), .A2(new_n318), .A3(KEYINPUT76), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT76), .B1(new_n316), .B2(new_n318), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n328), .B1(new_n333), .B2(new_n289), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n310), .B(new_n323), .C1(new_n330), .C2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT5), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n223), .A2(new_n319), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(new_n324), .ZN(new_n338));
  INV_X1    g137(.A(new_n310), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n336), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n324), .A2(new_n328), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n323), .A2(KEYINPUT4), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n333), .A2(new_n289), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n339), .A2(KEYINPUT5), .ZN(new_n345));
  AOI22_X1  g144(.A1(new_n335), .A2(new_n340), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  XOR2_X1   g145(.A(G1gat), .B(G29gat), .Z(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G57gat), .B(G85gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT6), .B1(new_n346), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n335), .A2(new_n340), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n344), .A2(new_n345), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(new_n351), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n356), .A2(KEYINPUT6), .A3(new_n351), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  XOR2_X1   g160(.A(G211gat), .B(G218gat), .Z(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT72), .B(G211gat), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT22), .B1(new_n363), .B2(G218gat), .ZN(new_n364));
  XOR2_X1   g163(.A(G197gat), .B(G204gat), .Z(new_n365));
  OAI21_X1  g164(.A(new_n362), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(G211gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT72), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT72), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(G211gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n368), .A2(new_n370), .A3(G218gat), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT22), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n362), .ZN(new_n374));
  INV_X1    g173(.A(new_n365), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n366), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(G226gat), .A2(G233gat), .ZN(new_n378));
  XOR2_X1   g177(.A(new_n378), .B(KEYINPUT73), .Z(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n380), .B1(new_n257), .B2(new_n275), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT29), .B1(new_n284), .B2(new_n287), .ZN(new_n382));
  INV_X1    g181(.A(new_n378), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n377), .B(new_n381), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT74), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT29), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n386), .B1(new_n257), .B2(new_n275), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n284), .A2(new_n287), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n387), .A2(new_n379), .B1(new_n388), .B2(new_n383), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n384), .B(new_n385), .C1(new_n389), .C2(new_n377), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n383), .B1(new_n257), .B2(new_n275), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n392), .B1(new_n382), .B2(new_n380), .ZN(new_n393));
  INV_X1    g192(.A(new_n377), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n385), .B1(new_n395), .B2(new_n384), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT37), .B1(new_n391), .B2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G8gat), .B(G36gat), .ZN(new_n398));
  INV_X1    g197(.A(G64gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(G92gat), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT85), .B(KEYINPUT37), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n395), .A2(new_n384), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n397), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT38), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n384), .B(new_n401), .C1(new_n389), .C2(new_n377), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT38), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n394), .B(new_n381), .C1(new_n382), .C2(new_n383), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n409), .B(KEYINPUT37), .C1(new_n389), .C2(new_n394), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n404), .A2(new_n408), .A3(new_n410), .A4(new_n402), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n361), .A2(new_n406), .A3(new_n407), .A4(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT29), .B1(new_n366), .B2(new_n376), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n321), .B1(new_n413), .B2(KEYINPUT81), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT81), .ZN(new_n415));
  AOI211_X1 g214(.A(new_n415), .B(KEYINPUT29), .C1(new_n366), .C2(new_n376), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n319), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT82), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n322), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n394), .B1(KEYINPUT29), .B2(new_n420), .ZN(new_n421));
  OAI211_X1 g220(.A(KEYINPUT82), .B(new_n319), .C1(new_n414), .C2(new_n416), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n419), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(G228gat), .ZN(new_n424));
  INV_X1    g223(.A(G233gat), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n426), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n421), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n366), .A2(KEYINPUT80), .A3(new_n376), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n386), .ZN(new_n431));
  NOR3_X1   g230(.A1(new_n366), .A2(KEYINPUT80), .A3(new_n374), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n321), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n333), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n429), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n427), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G78gat), .B(G106gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(KEYINPUT31), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G22gat), .B(G50gat), .ZN(new_n441));
  INV_X1    g240(.A(new_n439), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n427), .A2(new_n442), .A3(new_n436), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n440), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n441), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n442), .B1(new_n427), .B2(new_n436), .ZN(new_n446));
  AOI211_X1 g245(.A(new_n439), .B(new_n435), .C1(new_n423), .C2(new_n426), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n344), .A2(new_n310), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT39), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n337), .A2(new_n310), .A3(new_n324), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n453), .B(KEYINPUT39), .C1(new_n344), .C2(new_n310), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n452), .A2(new_n454), .A3(KEYINPUT40), .A4(new_n352), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT84), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n455), .B(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n351), .B1(new_n450), .B2(new_n451), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n454), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT83), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT40), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT83), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n458), .A2(new_n462), .A3(new_n454), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n460), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n402), .B1(new_n391), .B2(new_n396), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT30), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n407), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n407), .A2(new_n466), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT75), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT75), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n407), .A2(new_n471), .A3(new_n466), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n465), .A2(new_n468), .A3(new_n470), .A4(new_n472), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n457), .A2(new_n357), .A3(new_n464), .A4(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n412), .A2(new_n449), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n356), .A2(KEYINPUT79), .A3(new_n351), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT79), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n477), .B1(new_n346), .B2(new_n352), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n476), .A2(new_n478), .A3(new_n353), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n359), .ZN(new_n480));
  INV_X1    g279(.A(new_n473), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n444), .A2(new_n448), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n309), .A2(new_n475), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n294), .A2(new_n302), .A3(new_n304), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n304), .A2(new_n302), .ZN(new_n487));
  INV_X1    g286(.A(new_n294), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n444), .A2(new_n448), .A3(new_n486), .A4(new_n489), .ZN(new_n490));
  OAI211_X1 g289(.A(KEYINPUT87), .B(KEYINPUT35), .C1(new_n490), .C2(new_n482), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n473), .B1(new_n359), .B2(new_n479), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n493), .A2(new_n444), .A3(new_n308), .A4(new_n448), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT87), .B1(new_n494), .B2(KEYINPUT35), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT35), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n481), .A2(new_n497), .A3(new_n360), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT86), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n499), .A2(new_n500), .A3(new_n449), .A4(new_n308), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT86), .B1(new_n490), .B2(new_n498), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n485), .B1(new_n496), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(G230gat), .A2(G233gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(G99gat), .A2(G106gat), .ZN(new_n506));
  INV_X1    g305(.A(G85gat), .ZN(new_n507));
  INV_X1    g306(.A(G92gat), .ZN(new_n508));
  AOI22_X1  g307(.A1(KEYINPUT8), .A2(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT97), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n509), .B(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(G85gat), .A2(G92gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(KEYINPUT7), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  XOR2_X1   g313(.A(G99gat), .B(G106gat), .Z(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT9), .ZN(new_n517));
  INV_X1    g316(.A(G71gat), .ZN(new_n518));
  INV_X1    g317(.A(G78gat), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT95), .ZN(new_n521));
  XOR2_X1   g320(.A(G57gat), .B(G64gat), .Z(new_n522));
  INV_X1    g321(.A(KEYINPUT95), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n523), .B(new_n517), .C1(new_n518), .C2(new_n519), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n521), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G71gat), .B(G78gat), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n521), .A2(new_n522), .A3(new_n526), .A4(new_n524), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n515), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n511), .A2(new_n531), .A3(new_n513), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n531), .A2(KEYINPUT98), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n516), .A2(new_n530), .A3(new_n532), .A4(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n533), .A2(new_n528), .A3(new_n529), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n511), .A2(new_n531), .A3(new_n513), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n531), .B1(new_n511), .B2(new_n513), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n505), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT99), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(G120gat), .B(G148gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(new_n249), .ZN(new_n543));
  INV_X1    g342(.A(G204gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n546), .B1(new_n539), .B2(new_n540), .ZN(new_n547));
  INV_X1    g346(.A(new_n505), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT10), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n534), .A2(new_n538), .A3(new_n549), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n536), .A2(new_n537), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n551), .A2(KEYINPUT10), .A3(new_n530), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n548), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  OR3_X1    g352(.A1(new_n541), .A2(new_n547), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n545), .B1(new_n553), .B2(new_n539), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n504), .A2(new_n556), .ZN(new_n557));
  OR2_X1    g356(.A1(G15gat), .A2(G22gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(G15gat), .A2(G22gat), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n558), .A2(KEYINPUT88), .A3(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT88), .ZN(new_n561));
  AND2_X1   g360(.A1(G15gat), .A2(G22gat), .ZN(new_n562));
  NOR2_X1   g361(.A1(G15gat), .A2(G22gat), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(G1gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT16), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT89), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n560), .A2(new_n564), .A3(new_n566), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT90), .B(G8gat), .ZN(new_n572));
  AND2_X1   g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n565), .A2(KEYINPUT89), .A3(new_n567), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n570), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n568), .A2(new_n571), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(G8gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n578), .B1(KEYINPUT21), .B2(new_n530), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(G183gat), .ZN(new_n580));
  XOR2_X1   g379(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n530), .A2(KEYINPUT21), .ZN(new_n583));
  XOR2_X1   g382(.A(G127gat), .B(G155gat), .Z(new_n584));
  XOR2_X1   g383(.A(new_n583), .B(new_n584), .Z(new_n585));
  XOR2_X1   g384(.A(KEYINPUT96), .B(G211gat), .Z(new_n586));
  NAND2_X1  g385(.A1(G231gat), .A2(G233gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n585), .B(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n582), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n582), .A2(new_n590), .ZN(new_n592));
  AND2_X1   g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT14), .ZN(new_n594));
  INV_X1    g393(.A(G29gat), .ZN(new_n595));
  INV_X1    g394(.A(G36gat), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n597), .A2(new_n598), .B1(G29gat), .B2(G36gat), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G43gat), .B(G50gat), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n600), .A2(KEYINPUT15), .A3(new_n601), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n601), .A2(KEYINPUT15), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(KEYINPUT15), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n603), .A2(new_n604), .A3(new_n599), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n551), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n602), .A2(new_n605), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(KEYINPUT17), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT17), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n607), .B(new_n608), .C1(new_n613), .C2(new_n551), .ZN(new_n614));
  XNOR2_X1  g413(.A(G134gat), .B(G162gat), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n614), .B(new_n615), .Z(new_n616));
  XNOR2_X1  g415(.A(G190gat), .B(G218gat), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n616), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT18), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n610), .A2(new_n577), .A3(new_n575), .A4(new_n612), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n578), .A2(new_n606), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(G229gat), .A2(G233gat), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n628), .B(KEYINPUT91), .Z(new_n629));
  OAI21_X1  g428(.A(new_n624), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n575), .A2(new_n609), .A3(new_n577), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(KEYINPUT92), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT92), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n575), .A2(new_n609), .A3(new_n577), .A4(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n632), .A2(new_n626), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n629), .B(KEYINPUT13), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n629), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n625), .A2(KEYINPUT18), .A3(new_n638), .A4(new_n626), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT11), .B(G169gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G197gat), .ZN(new_n641));
  XOR2_X1   g440(.A(G113gat), .B(G141gat), .Z(new_n642));
  XOR2_X1   g441(.A(new_n641), .B(new_n642), .Z(new_n643));
  XOR2_X1   g442(.A(new_n643), .B(KEYINPUT12), .Z(new_n644));
  NAND4_X1  g443(.A1(new_n630), .A2(new_n637), .A3(new_n639), .A4(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n644), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n637), .A2(new_n639), .A3(KEYINPUT93), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n630), .ZN(new_n648));
  AOI21_X1  g447(.A(KEYINPUT93), .B1(new_n637), .B2(new_n639), .ZN(new_n649));
  OAI211_X1 g448(.A(KEYINPUT94), .B(new_n646), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n637), .A2(new_n639), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT93), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n654), .A2(new_n630), .A3(new_n647), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT94), .B1(new_n655), .B2(new_n646), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n645), .B1(new_n651), .B2(new_n656), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n557), .A2(new_n593), .A3(new_n623), .A4(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n658), .A2(new_n480), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(new_n566), .ZN(G1324gat));
  NOR2_X1   g459(.A1(new_n658), .A2(new_n481), .ZN(new_n661));
  NAND2_X1  g460(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n662));
  OR2_X1    g461(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT42), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  INV_X1    g466(.A(G8gat), .ZN(new_n668));
  OAI211_X1 g467(.A(new_n666), .B(new_n667), .C1(new_n668), .C2(new_n661), .ZN(G1325gat));
  INV_X1    g468(.A(G15gat), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n658), .A2(new_n670), .A3(new_n309), .ZN(new_n671));
  INV_X1    g470(.A(new_n308), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n670), .B1(new_n658), .B2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT100), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n674), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n671), .B1(new_n675), .B2(new_n676), .ZN(G1326gat));
  NOR2_X1   g476(.A1(new_n658), .A2(new_n449), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT43), .B(G22gat), .Z(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1327gat));
  INV_X1    g479(.A(new_n645), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT94), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n681), .B1(new_n684), .B2(new_n650), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n593), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n557), .A2(new_n622), .A3(new_n686), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n687), .A2(G29gat), .A3(new_n480), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT45), .Z(new_n689));
  INV_X1    g488(.A(KEYINPUT102), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n691), .B1(new_n504), .B2(new_n623), .ZN(new_n692));
  OAI21_X1  g491(.A(KEYINPUT35), .B1(new_n490), .B2(new_n482), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT87), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n695), .A2(new_n491), .A3(new_n502), .A4(new_n501), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n309), .A2(new_n475), .A3(new_n484), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n623), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(KEYINPUT44), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n692), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n591), .A2(new_n592), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT101), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n702), .A2(new_n685), .A3(new_n556), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n690), .B1(new_n704), .B2(new_n480), .ZN(new_n705));
  INV_X1    g504(.A(new_n480), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n700), .A2(KEYINPUT102), .A3(new_n706), .A4(new_n703), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n705), .A2(G29gat), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n689), .A2(new_n708), .ZN(G1328gat));
  NOR2_X1   g508(.A1(new_n481), .A2(G36gat), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n557), .A2(new_n622), .A3(new_n686), .A4(new_n710), .ZN(new_n711));
  OR2_X1    g510(.A1(new_n711), .A2(KEYINPUT103), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(KEYINPUT103), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(KEYINPUT104), .B1(new_n714), .B2(KEYINPUT46), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(KEYINPUT46), .ZN(new_n716));
  OAI21_X1  g515(.A(G36gat), .B1(new_n704), .B2(new_n481), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT104), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT46), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n712), .A2(new_n718), .A3(new_n719), .A4(new_n713), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n715), .A2(new_n716), .A3(new_n717), .A4(new_n720), .ZN(G1329gat));
  OR3_X1    g520(.A1(new_n687), .A2(G43gat), .A3(new_n672), .ZN(new_n722));
  INV_X1    g521(.A(new_n309), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n692), .A2(new_n723), .A3(new_n699), .A4(new_n703), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(G43gat), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT105), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(KEYINPUT47), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT47), .ZN(new_n728));
  AOI211_X1 g527(.A(KEYINPUT105), .B(new_n728), .C1(new_n722), .C2(new_n725), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n727), .A2(new_n729), .ZN(G1330gat));
  OAI21_X1  g529(.A(G50gat), .B1(new_n704), .B2(new_n449), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT48), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT106), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n687), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(G50gat), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n557), .A2(KEYINPUT106), .A3(new_n622), .A4(new_n686), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n734), .A2(new_n735), .A3(new_n483), .A4(new_n736), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n731), .A2(new_n732), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n732), .B1(new_n731), .B2(new_n737), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(G1331gat));
  NAND3_X1  g539(.A1(new_n593), .A2(new_n623), .A3(new_n685), .ZN(new_n741));
  INV_X1    g540(.A(new_n556), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT107), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n696), .A2(new_n697), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n706), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g547(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n746), .A2(new_n473), .A3(new_n749), .ZN(new_n750));
  OR2_X1    g549(.A1(new_n750), .A2(KEYINPUT108), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(KEYINPUT108), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1333gat));
  NAND3_X1  g554(.A1(new_n746), .A2(G71gat), .A3(new_n723), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n744), .A2(new_n308), .A3(new_n745), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n756), .B1(G71gat), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(KEYINPUT109), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT109), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n756), .B(new_n760), .C1(G71gat), .C2(new_n757), .ZN(new_n761));
  AND3_X1   g560(.A1(new_n759), .A2(KEYINPUT50), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT50), .B1(new_n759), .B2(new_n761), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(G1334gat));
  NAND2_X1  g563(.A1(new_n746), .A2(new_n483), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g565(.A1(new_n685), .A2(new_n701), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT110), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n768), .A2(new_n556), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n700), .A2(new_n769), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n770), .A2(G85gat), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n745), .A2(new_n622), .A3(new_n768), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT111), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n698), .A2(KEYINPUT51), .A3(new_n768), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT51), .B1(new_n698), .B2(new_n768), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n742), .B1(new_n778), .B2(KEYINPUT111), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n777), .A2(new_n779), .A3(new_n706), .ZN(new_n780));
  AOI22_X1  g579(.A1(new_n771), .A2(new_n706), .B1(new_n507), .B2(new_n780), .ZN(G1336gat));
  NOR2_X1   g580(.A1(new_n481), .A2(G92gat), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n777), .A2(new_n779), .A3(new_n782), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n692), .A2(new_n473), .A3(new_n699), .A4(new_n769), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT52), .B1(new_n784), .B2(G92gat), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n784), .A2(G92gat), .ZN(new_n788));
  INV_X1    g587(.A(new_n776), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n556), .B(new_n782), .C1(new_n789), .C2(new_n778), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n787), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(KEYINPUT112), .B1(new_n786), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n783), .A2(new_n785), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n788), .A2(new_n790), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n793), .B(new_n794), .C1(new_n795), .C2(new_n787), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n792), .A2(new_n796), .ZN(G1337gat));
  NAND3_X1  g596(.A1(new_n770), .A2(KEYINPUT113), .A3(new_n723), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n700), .A2(new_n723), .A3(new_n769), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT113), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n798), .A2(G99gat), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n777), .A2(new_n779), .ZN(new_n803));
  OR2_X1    g602(.A1(new_n803), .A2(G99gat), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n672), .B2(new_n804), .ZN(G1338gat));
  NAND4_X1  g604(.A1(new_n692), .A2(new_n483), .A3(new_n699), .A4(new_n769), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(G106gat), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT114), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n449), .A2(G106gat), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n556), .B(new_n809), .C1(new_n789), .C2(new_n778), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT115), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n742), .B1(new_n774), .B2(new_n776), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n812), .A2(new_n813), .A3(new_n809), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n806), .A2(new_n815), .A3(G106gat), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n808), .A2(new_n811), .A3(new_n814), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT53), .ZN(new_n818));
  XNOR2_X1  g617(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n819));
  INV_X1    g618(.A(new_n809), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n807), .B(new_n819), .C1(new_n803), .C2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n818), .A2(new_n821), .ZN(G1339gat));
  NAND4_X1  g621(.A1(new_n593), .A2(new_n623), .A3(new_n685), .A4(new_n742), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT117), .ZN(new_n824));
  INV_X1    g623(.A(new_n823), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT117), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n550), .A2(new_n548), .A3(new_n552), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT54), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n829), .A2(new_n553), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  XNOR2_X1  g630(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  AOI211_X1 g632(.A(new_n548), .B(new_n833), .C1(new_n550), .C2(new_n552), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n834), .A2(KEYINPUT119), .A3(new_n546), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT119), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n553), .A2(new_n832), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n836), .B1(new_n837), .B2(new_n545), .ZN(new_n838));
  OAI211_X1 g637(.A(KEYINPUT55), .B(new_n831), .C1(new_n835), .C2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n554), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n831), .B1(new_n835), .B2(new_n838), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT55), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n841), .A2(KEYINPUT120), .A3(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT120), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT119), .B1(new_n834), .B2(new_n546), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n837), .A2(new_n836), .A3(new_n545), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n830), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n844), .B1(new_n847), .B2(KEYINPUT55), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n840), .B1(new_n843), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n635), .A2(new_n636), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n850), .B1(new_n629), .B2(new_n627), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n851), .A2(new_n643), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n645), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n849), .A2(new_n622), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n853), .A2(new_n742), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n856), .B1(new_n849), .B2(new_n657), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n855), .B1(new_n857), .B2(new_n622), .ZN(new_n858));
  INV_X1    g657(.A(new_n702), .ZN(new_n859));
  AOI22_X1  g658(.A1(new_n824), .A2(new_n827), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n860), .A2(new_n490), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n480), .A2(new_n473), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n657), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g664(.A1(new_n863), .A2(new_n556), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g666(.A1(new_n863), .A2(new_n593), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n208), .A2(new_n209), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n859), .A2(new_n869), .ZN(new_n870));
  AOI22_X1  g669(.A1(new_n868), .A2(new_n869), .B1(new_n863), .B2(new_n870), .ZN(G1342gat));
  NAND2_X1  g670(.A1(new_n863), .A2(new_n622), .ZN(new_n872));
  NOR2_X1   g671(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n873));
  AND2_X1   g672(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n875), .B1(new_n872), .B2(new_n873), .ZN(G1343gat));
  NAND2_X1  g675(.A1(new_n827), .A2(new_n824), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n858), .A2(new_n859), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n879), .A2(new_n880), .A3(new_n483), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n847), .A2(KEYINPUT55), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n840), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n856), .B1(new_n657), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n855), .B1(new_n884), .B2(new_n622), .ZN(new_n885));
  AOI22_X1  g684(.A1(new_n827), .A2(new_n824), .B1(new_n885), .B2(new_n701), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT57), .B1(new_n886), .B2(new_n449), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n309), .A2(new_n862), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n881), .A2(new_n887), .A3(new_n657), .A4(new_n889), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n860), .A2(new_n449), .A3(new_n888), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n685), .A2(G141gat), .ZN(new_n892));
  AOI22_X1  g691(.A1(new_n890), .A2(G141gat), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OR2_X1    g694(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n895), .B(new_n896), .ZN(G1344gat));
  XNOR2_X1  g696(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n825), .B1(new_n885), .B2(new_n701), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n880), .B1(new_n899), .B2(new_n449), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT124), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n879), .A2(KEYINPUT57), .A3(new_n483), .ZN(new_n903));
  OAI211_X1 g702(.A(KEYINPUT124), .B(new_n880), .C1(new_n899), .C2(new_n449), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n905), .A2(new_n556), .A3(new_n889), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n898), .B1(new_n906), .B2(G148gat), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n881), .A2(new_n887), .A3(new_n889), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n908), .A2(new_n742), .ZN(new_n909));
  INV_X1    g708(.A(G148gat), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n909), .A2(KEYINPUT59), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n891), .A2(new_n910), .A3(new_n556), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n912), .A2(KEYINPUT122), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n912), .A2(KEYINPUT122), .ZN(new_n914));
  OAI22_X1  g713(.A1(new_n907), .A2(new_n911), .B1(new_n913), .B2(new_n914), .ZN(G1345gat));
  AOI21_X1  g714(.A(G155gat), .B1(new_n891), .B2(new_n593), .ZN(new_n916));
  INV_X1    g715(.A(G155gat), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n908), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n916), .B1(new_n918), .B2(new_n702), .ZN(G1346gat));
  AOI21_X1  g718(.A(G162gat), .B1(new_n891), .B2(new_n622), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n908), .A2(new_n623), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g721(.A1(new_n706), .A2(new_n481), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n861), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n657), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n250), .A2(new_n251), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT125), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT125), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n929), .B1(new_n925), .B2(G169gat), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n928), .B1(new_n927), .B2(new_n930), .ZN(G1348gat));
  NAND2_X1  g730(.A1(new_n924), .A2(new_n556), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g732(.A1(new_n861), .A2(new_n702), .A3(new_n923), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(KEYINPUT126), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT126), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n861), .A2(new_n936), .A3(new_n702), .A4(new_n923), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n935), .A2(G183gat), .A3(new_n937), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n924), .B(new_n593), .C1(new_n260), .C2(new_n259), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT60), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT60), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n938), .A2(new_n942), .A3(new_n939), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(G1350gat));
  NAND2_X1  g743(.A1(new_n924), .A2(new_n622), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n945), .A2(new_n946), .A3(new_n258), .ZN(new_n947));
  XOR2_X1   g746(.A(KEYINPUT61), .B(G190gat), .Z(new_n948));
  AOI21_X1  g747(.A(new_n947), .B1(new_n945), .B2(new_n948), .ZN(G1351gat));
  NAND2_X1  g748(.A1(new_n309), .A2(new_n923), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n905), .A2(new_n657), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(G197gat), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n860), .A2(new_n449), .A3(new_n950), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  OR2_X1    g754(.A1(new_n685), .A2(G197gat), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n953), .B1(new_n955), .B2(new_n956), .ZN(G1352gat));
  NAND3_X1  g756(.A1(new_n905), .A2(new_n556), .A3(new_n951), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(G204gat), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT62), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n954), .A2(new_n960), .A3(new_n544), .A4(new_n556), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n879), .A2(new_n544), .A3(new_n483), .A4(new_n951), .ZN(new_n962));
  OAI21_X1  g761(.A(KEYINPUT62), .B1(new_n962), .B2(new_n742), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n959), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(KEYINPUT127), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT127), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n959), .A2(new_n964), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n966), .A2(new_n968), .ZN(G1353gat));
  OR3_X1    g768(.A1(new_n955), .A2(new_n701), .A3(new_n363), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n905), .A2(new_n593), .A3(new_n951), .ZN(new_n971));
  AND3_X1   g770(.A1(new_n971), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n972));
  AOI21_X1  g771(.A(KEYINPUT63), .B1(new_n971), .B2(G211gat), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n970), .B1(new_n972), .B2(new_n973), .ZN(G1354gat));
  NAND3_X1  g773(.A1(new_n905), .A2(new_n622), .A3(new_n951), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(G218gat), .ZN(new_n976));
  OR2_X1    g775(.A1(new_n623), .A2(G218gat), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n976), .B1(new_n955), .B2(new_n977), .ZN(G1355gat));
endmodule


