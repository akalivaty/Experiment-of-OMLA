//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 0 0 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 0 0 1 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n593, new_n594, new_n595, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n637,
    new_n638, new_n641, new_n643, new_n644, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1203, new_n1204, new_n1205, new_n1206;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT65), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n459), .A2(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G101), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT69), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n460), .A2(KEYINPUT69), .A3(G101), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n466), .A2(new_n468), .A3(G137), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT70), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT70), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n465), .A2(new_n473), .A3(new_n470), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n466), .A2(new_n468), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT66), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT66), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n478), .A2(G125), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(G113), .A2(G2104), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT67), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n469), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n484));
  OR2_X1    g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI211_X1 g060(.A(KEYINPUT68), .B(new_n469), .C1(new_n480), .C2(new_n482), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n475), .B1(new_n485), .B2(new_n487), .ZN(G160));
  NOR2_X1   g063(.A1(new_n476), .A2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G136), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n476), .A2(new_n469), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G124), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT71), .B1(G100), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NOR3_X1   g069(.A1(KEYINPUT71), .A2(G100), .A3(G2105), .ZN(new_n495));
  OAI221_X1 g070(.A(G2104), .B1(G112), .B2(new_n469), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n490), .A2(new_n492), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G162));
  OR2_X1    g073(.A1(G102), .A2(G2105), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n499), .B(G2104), .C1(G114), .C2(new_n469), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n466), .A2(new_n468), .A3(G126), .A4(G2105), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n469), .A2(G138), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT72), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT72), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n503), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n478), .A2(new_n479), .A3(new_n508), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n466), .A2(new_n468), .A3(G138), .A4(new_n469), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT4), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n502), .B1(new_n509), .B2(new_n511), .ZN(G164));
  OR2_X1    g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  AND2_X1   g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  AND2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  OAI21_X1  g099(.A(G543), .B1(new_n521), .B2(new_n522), .ZN(new_n525));
  INV_X1    g100(.A(G50), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n523), .A2(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n518), .A2(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  XNOR2_X1  g104(.A(KEYINPUT6), .B(G651), .ZN(new_n530));
  AOI21_X1  g105(.A(KEYINPUT73), .B1(new_n530), .B2(G543), .ZN(new_n531));
  OAI211_X1 g106(.A(KEYINPUT73), .B(G543), .C1(new_n521), .C2(new_n522), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  OAI21_X1  g108(.A(G51), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g109(.A(G89), .B1(new_n521), .B2(new_n522), .ZN(new_n535));
  NAND2_X1  g110(.A1(G63), .A2(G651), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(KEYINPUT7), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n538), .A2(KEYINPUT7), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n537), .A2(new_n515), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n534), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(G168));
  NAND2_X1  g118(.A1(G77), .A2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n520), .A2(new_n519), .ZN(new_n545));
  INV_X1    g120(.A(G64), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  OR2_X1    g122(.A1(KEYINPUT6), .A2(G651), .ZN(new_n548));
  NAND2_X1  g123(.A1(KEYINPUT6), .A2(G651), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n513), .A2(new_n514), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n547), .A2(G651), .B1(new_n550), .B2(G90), .ZN(new_n551));
  XOR2_X1   g126(.A(KEYINPUT74), .B(G52), .Z(new_n552));
  OAI21_X1  g127(.A(new_n552), .B1(new_n531), .B2(new_n533), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n551), .A2(new_n553), .ZN(G301));
  INV_X1    g129(.A(G301), .ZN(G171));
  AOI22_X1  g130(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G81), .ZN(new_n557));
  OAI22_X1  g132(.A1(new_n556), .A2(new_n517), .B1(new_n557), .B2(new_n523), .ZN(new_n558));
  INV_X1    g133(.A(G43), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT73), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n525), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n559), .B1(new_n561), .B2(new_n532), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(new_n564));
  XOR2_X1   g139(.A(new_n564), .B(KEYINPUT75), .Z(G153));
  AND3_X1   g140(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G36), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT76), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  XOR2_X1   g146(.A(new_n571), .B(KEYINPUT77), .Z(G188));
  INV_X1    g147(.A(G543), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n573), .B1(new_n548), .B2(new_n549), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n574), .A2(new_n575), .A3(G53), .ZN(new_n576));
  INV_X1    g151(.A(G53), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT9), .B1(new_n525), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n576), .A2(new_n578), .B1(G91), .B2(new_n550), .ZN(new_n579));
  INV_X1    g154(.A(G65), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n513), .A2(new_n581), .A3(new_n514), .ZN(new_n582));
  OAI21_X1  g157(.A(KEYINPUT78), .B1(new_n520), .B2(new_n519), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n580), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AND2_X1   g159(.A1(G78), .A2(G543), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n579), .A2(new_n586), .ZN(G299));
  NAND2_X1  g162(.A1(new_n540), .A2(new_n539), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n530), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n589), .B2(new_n545), .ZN(new_n590));
  INV_X1    g165(.A(G51), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n591), .B1(new_n561), .B2(new_n532), .ZN(new_n592));
  NOR3_X1   g167(.A1(new_n590), .A2(new_n592), .A3(KEYINPUT79), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT79), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n594), .B1(new_n534), .B2(new_n541), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n593), .A2(new_n595), .ZN(G286));
  NAND2_X1  g171(.A1(new_n550), .A2(G87), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n574), .A2(G49), .ZN(new_n598));
  OAI21_X1  g173(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(G288));
  INV_X1    g175(.A(G86), .ZN(new_n601));
  INV_X1    g176(.A(G48), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n523), .A2(new_n601), .B1(new_n525), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(G73), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G61), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n545), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G651), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n603), .B1(new_n607), .B2(KEYINPUT80), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n515), .A2(G61), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n517), .B1(new_n609), .B2(new_n604), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT80), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n608), .A2(new_n612), .ZN(G305));
  NAND2_X1  g188(.A1(new_n561), .A2(new_n532), .ZN(new_n614));
  AND2_X1   g189(.A1(new_n614), .A2(G47), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n616));
  INV_X1    g191(.A(G85), .ZN(new_n617));
  OAI22_X1  g192(.A1(new_n616), .A2(new_n517), .B1(new_n617), .B2(new_n523), .ZN(new_n618));
  OR3_X1    g193(.A1(new_n615), .A2(KEYINPUT81), .A3(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(KEYINPUT81), .B1(new_n615), .B2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(G290));
  NAND2_X1  g196(.A1(G301), .A2(G868), .ZN(new_n622));
  INV_X1    g197(.A(G66), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n623), .B1(new_n582), .B2(new_n583), .ZN(new_n624));
  AND2_X1   g199(.A1(G79), .A2(G543), .ZN(new_n625));
  OAI21_X1  g200(.A(G651), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT10), .ZN(new_n627));
  INV_X1    g202(.A(G92), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n523), .B2(new_n628), .ZN(new_n629));
  NAND4_X1  g204(.A1(new_n515), .A2(new_n530), .A3(KEYINPUT10), .A4(G92), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(G54), .B1(new_n531), .B2(new_n533), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n626), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n622), .B1(new_n634), .B2(G868), .ZN(G284));
  OAI21_X1  g210(.A(new_n622), .B1(new_n634), .B2(G868), .ZN(G321));
  NOR2_X1   g211(.A1(G299), .A2(G868), .ZN(new_n637));
  INV_X1    g212(.A(G286), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n637), .B1(new_n638), .B2(G868), .ZN(G280));
  XOR2_X1   g214(.A(G280), .B(KEYINPUT82), .Z(G297));
  INV_X1    g215(.A(G559), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n634), .B1(new_n641), .B2(G860), .ZN(G148));
  NAND2_X1  g217(.A1(new_n634), .A2(new_n641), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(G868), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(G868), .B2(new_n563), .ZN(G323));
  XNOR2_X1  g220(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g221(.A1(new_n478), .A2(new_n479), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(new_n460), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT12), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT13), .ZN(new_n650));
  INV_X1    g225(.A(G2100), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n489), .A2(G135), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n491), .A2(G123), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n469), .A2(G111), .ZN(new_n656));
  OAI21_X1  g231(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n657));
  OAI211_X1 g232(.A(new_n654), .B(new_n655), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(G2096), .Z(new_n659));
  NAND3_X1  g234(.A1(new_n652), .A2(new_n653), .A3(new_n659), .ZN(G156));
  INV_X1    g235(.A(KEYINPUT14), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2427), .B(G2438), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2430), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT15), .B(G2435), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n661), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n665), .B1(new_n664), .B2(new_n663), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2451), .B(G2454), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT16), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1341), .B(G1348), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n666), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2443), .B(G2446), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  AND3_X1   g249(.A1(new_n673), .A2(G14), .A3(new_n674), .ZN(G401));
  XNOR2_X1  g250(.A(G2072), .B(G2078), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT17), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2067), .B(G2678), .ZN(new_n678));
  XOR2_X1   g253(.A(G2084), .B(G2090), .Z(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  NOR3_X1   g255(.A1(new_n677), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT83), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n677), .A2(new_n678), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n683), .B(new_n680), .C1(new_n676), .C2(new_n678), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n679), .A2(new_n676), .A3(new_n678), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT18), .Z(new_n686));
  NAND3_X1  g261(.A1(new_n682), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G2096), .B(G2100), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(G227));
  XOR2_X1   g265(.A(G1971), .B(G1976), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT19), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1956), .B(G2474), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1961), .B(G1966), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  NOR3_X1   g271(.A1(new_n692), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n692), .A2(new_n695), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT20), .Z(new_n699));
  AOI211_X1 g274(.A(new_n697), .B(new_n699), .C1(new_n692), .C2(new_n696), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1991), .B(G1996), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1981), .B(G1986), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(G229));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G6), .ZN(new_n708));
  INV_X1    g283(.A(G305), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(new_n707), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT32), .B(G1981), .Z(new_n711));
  XOR2_X1   g286(.A(new_n710), .B(new_n711), .Z(new_n712));
  NAND2_X1  g287(.A1(new_n707), .A2(G23), .ZN(new_n713));
  INV_X1    g288(.A(G288), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(new_n707), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT85), .Z(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT33), .B(G1976), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n716), .A2(new_n717), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n707), .A2(G22), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G166), .B2(new_n707), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G1971), .ZN(new_n722));
  NOR4_X1   g297(.A1(new_n712), .A2(new_n718), .A3(new_n719), .A4(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT34), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n723), .A2(new_n724), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n491), .A2(G119), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n469), .A2(G107), .ZN(new_n728));
  OAI21_X1  g303(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G131), .B2(new_n489), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT84), .Z(new_n732));
  MUX2_X1   g307(.A(G25), .B(new_n732), .S(G29), .Z(new_n733));
  XOR2_X1   g308(.A(KEYINPUT35), .B(G1991), .Z(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  MUX2_X1   g310(.A(G24), .B(G290), .S(G16), .Z(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(G1986), .Z(new_n737));
  NAND4_X1  g312(.A1(new_n725), .A2(new_n726), .A3(new_n735), .A4(new_n737), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT36), .Z(new_n739));
  INV_X1    g314(.A(G29), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G35), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G162), .B2(new_n740), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT29), .Z(new_n743));
  INV_X1    g318(.A(G2090), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n647), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n746), .A2(new_n469), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT25), .Z(new_n749));
  NAND2_X1  g324(.A1(new_n489), .A2(G139), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G29), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G29), .B2(G33), .ZN(new_n754));
  INV_X1    g329(.A(G2072), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT24), .ZN(new_n757));
  INV_X1    g332(.A(G34), .ZN(new_n758));
  AOI21_X1  g333(.A(G29), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n757), .B2(new_n758), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G160), .B2(new_n740), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(G2084), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n707), .A2(G21), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G168), .B2(new_n707), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT91), .B(G1966), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n745), .A2(new_n756), .A3(new_n762), .A4(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n754), .A2(new_n755), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT90), .Z(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G2084), .B2(new_n761), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n740), .A2(G26), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT28), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n489), .A2(G140), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n491), .A2(G128), .ZN(new_n774));
  NOR2_X1   g349(.A1(G104), .A2(G2105), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT87), .Z(new_n776));
  OAI21_X1  g351(.A(G2104), .B1(new_n469), .B2(G116), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n773), .B(new_n774), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT88), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(G29), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n780), .A2(KEYINPUT89), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n780), .A2(KEYINPUT89), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n772), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(G2067), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n563), .A2(new_n707), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n707), .B2(G19), .ZN(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n788), .A2(G1341), .ZN(new_n789));
  NOR2_X1   g364(.A1(G27), .A2(G29), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G164), .B2(G29), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT94), .B(G2078), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n788), .A2(G1341), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n789), .A2(new_n793), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(G4), .A2(G16), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT86), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(new_n633), .B2(new_n707), .ZN(new_n799));
  INV_X1    g374(.A(G1348), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n740), .A2(G32), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n489), .A2(G141), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n491), .A2(G129), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n460), .A2(G105), .ZN(new_n805));
  NAND3_X1  g380(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT26), .Z(new_n807));
  NAND4_X1  g382(.A1(new_n803), .A2(new_n804), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n802), .B1(new_n809), .B2(new_n740), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT27), .B(G1996), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(G5), .A2(G16), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT93), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(G301), .B2(new_n707), .ZN(new_n815));
  INV_X1    g390(.A(G1961), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT30), .B(G28), .ZN(new_n818));
  OR2_X1    g393(.A1(KEYINPUT31), .A2(G11), .ZN(new_n819));
  NAND2_X1  g394(.A1(KEYINPUT31), .A2(G11), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n818), .A2(new_n740), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n658), .B2(new_n740), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT92), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n815), .A2(new_n816), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n812), .A2(new_n817), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  NOR3_X1   g400(.A1(new_n796), .A2(new_n801), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n707), .A2(G20), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT23), .Z(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(G299), .B2(G16), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(G1956), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n743), .B2(new_n744), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT95), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n785), .A2(new_n826), .A3(new_n832), .ZN(new_n833));
  NOR4_X1   g408(.A1(new_n739), .A2(new_n767), .A3(new_n770), .A4(new_n833), .ZN(G311));
  INV_X1    g409(.A(G311), .ZN(G150));
  NAND2_X1  g410(.A1(new_n634), .A2(G559), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT38), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n838));
  INV_X1    g413(.A(G93), .ZN(new_n839));
  OAI22_X1  g414(.A1(new_n838), .A2(new_n517), .B1(new_n839), .B2(new_n523), .ZN(new_n840));
  INV_X1    g415(.A(G55), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(new_n561), .B2(new_n532), .ZN(new_n842));
  OAI22_X1  g417(.A1(new_n562), .A2(new_n558), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n562), .ZN(new_n844));
  NAND2_X1  g419(.A1(G68), .A2(G543), .ZN(new_n845));
  INV_X1    g420(.A(G56), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n845), .B1(new_n545), .B2(new_n846), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n847), .A2(G651), .B1(new_n550), .B2(G81), .ZN(new_n848));
  NAND2_X1  g423(.A1(G80), .A2(G543), .ZN(new_n849));
  INV_X1    g424(.A(G67), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n849), .B1(new_n545), .B2(new_n850), .ZN(new_n851));
  AOI22_X1  g426(.A1(new_n851), .A2(G651), .B1(new_n550), .B2(G93), .ZN(new_n852));
  OAI21_X1  g427(.A(G55), .B1(new_n531), .B2(new_n533), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n844), .A2(new_n848), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n843), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n837), .B(new_n856), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n857), .A2(KEYINPUT39), .ZN(new_n858));
  INV_X1    g433(.A(G860), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(KEYINPUT39), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n840), .A2(new_n842), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n862), .A2(new_n859), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT37), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT96), .ZN(G145));
  AOI22_X1  g441(.A1(G130), .A2(new_n491), .B1(new_n489), .B2(G142), .ZN(new_n867));
  OAI21_X1  g442(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n868));
  INV_X1    g443(.A(G118), .ZN(new_n869));
  AOI22_X1  g444(.A1(new_n868), .A2(KEYINPUT98), .B1(new_n869), .B2(G2105), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n870), .B1(KEYINPUT98), .B2(new_n868), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n649), .B(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n732), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT99), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT97), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(new_n747), .B2(new_n751), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n878), .A2(new_n809), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n809), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(G164), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n509), .A2(new_n511), .ZN(new_n883));
  INV_X1    g458(.A(new_n502), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n879), .A2(new_n885), .A3(new_n880), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n779), .ZN(new_n888));
  INV_X1    g463(.A(new_n779), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n882), .A2(new_n889), .A3(new_n886), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n876), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(KEYINPUT100), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT100), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n876), .A2(new_n891), .A3(new_n894), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n893), .B(new_n895), .C1(new_n891), .C2(new_n876), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n658), .B(new_n497), .ZN(new_n897));
  XOR2_X1   g472(.A(G160), .B(new_n897), .Z(new_n898));
  AOI21_X1  g473(.A(G37), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n888), .A2(new_n890), .A3(new_n874), .ZN(new_n900));
  INV_X1    g475(.A(new_n898), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n892), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT101), .ZN(new_n903));
  XNOR2_X1  g478(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n899), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n904), .B1(new_n899), .B2(new_n903), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(G395));
  XNOR2_X1  g482(.A(new_n643), .B(new_n855), .ZN(new_n908));
  AOI22_X1  g483(.A1(G54), .A2(new_n614), .B1(new_n629), .B2(new_n630), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n909), .A2(new_n586), .A3(new_n579), .A4(new_n626), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n633), .A2(G299), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n910), .A2(new_n911), .A3(KEYINPUT41), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT41), .B1(new_n910), .B2(new_n911), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n913), .B1(new_n908), .B2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT42), .ZN(new_n918));
  XNOR2_X1  g493(.A(G303), .B(G288), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n619), .A2(G305), .A3(new_n620), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(G305), .B1(new_n619), .B2(new_n620), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n923), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n925), .A2(new_n919), .A3(new_n921), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n918), .B(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(G868), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(G868), .B2(new_n862), .ZN(G295));
  OAI21_X1  g505(.A(new_n929), .B1(G868), .B2(new_n862), .ZN(G331));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n932));
  OAI21_X1  g507(.A(G171), .B1(new_n593), .B2(new_n595), .ZN(new_n933));
  NAND2_X1  g508(.A1(G301), .A2(new_n542), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n933), .A2(new_n843), .A3(new_n854), .A4(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT79), .B1(new_n590), .B2(new_n592), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n534), .A2(new_n541), .A3(new_n594), .ZN(new_n938));
  AOI21_X1  g513(.A(G301), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AND2_X1   g514(.A1(G301), .A2(new_n542), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n855), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n935), .A2(new_n936), .A3(new_n941), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n856), .A2(KEYINPUT106), .A3(new_n933), .A4(new_n934), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n912), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT104), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n935), .A2(new_n945), .A3(new_n941), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n855), .B(KEYINPUT104), .C1(new_n939), .C2(new_n940), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n946), .A2(new_n916), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT105), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n944), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n946), .A2(new_n916), .A3(new_n947), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT105), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n950), .A2(KEYINPUT107), .A3(new_n927), .A4(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n942), .A2(new_n943), .ZN(new_n954));
  INV_X1    g529(.A(new_n912), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n946), .A2(new_n916), .A3(new_n949), .A4(new_n947), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n952), .A2(new_n956), .A3(new_n927), .A4(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G37), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n942), .A2(new_n916), .A3(new_n943), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n942), .A2(new_n916), .A3(KEYINPUT108), .A4(new_n943), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n946), .A2(new_n947), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n955), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n927), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n953), .A2(new_n960), .A3(new_n961), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT109), .ZN(new_n972));
  AOI21_X1  g547(.A(G37), .B1(new_n958), .B2(new_n959), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT109), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n973), .A2(new_n974), .A3(new_n953), .A4(new_n970), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n972), .A2(KEYINPUT43), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n950), .A2(new_n952), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n969), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n978), .A2(new_n973), .A3(new_n953), .ZN(new_n979));
  XOR2_X1   g554(.A(KEYINPUT103), .B(KEYINPUT43), .Z(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n932), .B1(new_n976), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n979), .A2(new_n981), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n973), .A2(new_n953), .A3(new_n980), .A4(new_n970), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n984), .A2(new_n932), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT110), .B1(new_n983), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT110), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n979), .A2(new_n981), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT43), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n991), .B1(new_n971), .B2(KEYINPUT109), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n990), .B1(new_n992), .B2(new_n975), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n989), .B(new_n986), .C1(new_n993), .C2(new_n932), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n988), .A2(new_n994), .ZN(G397));
  AND3_X1   g570(.A1(new_n465), .A2(new_n473), .A3(new_n470), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n473), .B1(new_n465), .B2(new_n470), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n483), .A2(new_n484), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n998), .B(G40), .C1(new_n999), .C2(new_n486), .ZN(new_n1000));
  XOR2_X1   g575(.A(KEYINPUT111), .B(G1384), .Z(new_n1001));
  NAND2_X1  g576(.A1(new_n885), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1000), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(G1996), .A3(new_n808), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n1007), .B(KEYINPUT112), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n779), .B(G2067), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n1005), .ZN(new_n1010));
  INV_X1    g585(.A(G1996), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1005), .A2(new_n1011), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1008), .B(new_n1010), .C1(new_n808), .C2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n734), .ZN(new_n1014));
  OR3_X1    g589(.A1(new_n1013), .A2(new_n1014), .A3(new_n732), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n889), .A2(new_n784), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1006), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1005), .B1(new_n1009), .B2(new_n808), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1018), .B(KEYINPUT126), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n1012), .B(KEYINPUT46), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g596(.A(new_n1021), .B(KEYINPUT47), .Z(new_n1022));
  XNOR2_X1  g597(.A(new_n732), .B(new_n1014), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1013), .B1(new_n1005), .B2(new_n1023), .ZN(new_n1024));
  NOR3_X1   g599(.A1(new_n1006), .A2(G1986), .A3(G290), .ZN(new_n1025));
  XNOR2_X1  g600(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n1025), .B(new_n1026), .ZN(new_n1027));
  AOI211_X1 g602(.A(new_n1017), .B(new_n1022), .C1(new_n1024), .C2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1000), .ZN(new_n1029));
  NOR2_X1   g604(.A1(G164), .A2(G1384), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G1976), .ZN(new_n1032));
  NOR2_X1   g607(.A1(G288), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT52), .B1(G288), .B2(new_n1032), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1031), .A2(G8), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1030), .ZN(new_n1037));
  OAI21_X1  g612(.A(G8), .B1(new_n1000), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT52), .B1(new_n1038), .B2(new_n1033), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G1981), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n608), .A2(new_n1041), .A3(new_n612), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT115), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n608), .A2(new_n1044), .A3(new_n1041), .A4(new_n612), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n610), .B1(new_n1047), .B2(new_n603), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(new_n1047), .B2(new_n603), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(G1981), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1046), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT49), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1051), .A2(KEYINPUT117), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n1043), .A2(new_n1045), .B1(G1981), .B2(new_n1049), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1054), .B1(new_n1055), .B2(KEYINPUT49), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1038), .B1(KEYINPUT49), .B2(new_n1055), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1040), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n1060));
  INV_X1    g635(.A(G1384), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n885), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1029), .A2(new_n744), .A3(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1030), .A2(KEYINPUT45), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n885), .A2(KEYINPUT45), .A3(new_n1001), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n1000), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT113), .B(G1971), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1066), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT114), .ZN(new_n1074));
  NAND2_X1  g649(.A1(G303), .A2(G8), .ZN(new_n1075));
  XOR2_X1   g650(.A(new_n1075), .B(KEYINPUT55), .Z(new_n1076));
  INV_X1    g651(.A(KEYINPUT114), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1066), .B(new_n1077), .C1(new_n1070), .C2(new_n1072), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1074), .A2(G8), .A3(new_n1076), .A4(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1076), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1037), .A2(new_n1003), .ZN(new_n1081));
  NAND4_X1  g656(.A1(G160), .A2(new_n1081), .A3(G40), .A4(new_n1068), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1000), .A2(new_n1064), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1082), .A2(new_n1071), .B1(new_n1083), .B2(new_n744), .ZN(new_n1084));
  INV_X1    g659(.A(G8), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1080), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1059), .A2(new_n1079), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1029), .A2(new_n1065), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n800), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1029), .A2(new_n784), .A3(new_n1030), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1089), .B1(KEYINPUT122), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(KEYINPUT122), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n634), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  XOR2_X1   g669(.A(G299), .B(KEYINPUT57), .Z(new_n1095));
  XOR2_X1   g670(.A(KEYINPUT121), .B(G1956), .Z(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n1000), .B2(new_n1064), .ZN(new_n1097));
  XOR2_X1   g672(.A(KEYINPUT56), .B(G2072), .Z(new_n1098));
  OAI211_X1 g673(.A(new_n1095), .B(new_n1097), .C1(new_n1082), .C2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1094), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1098), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1070), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1095), .B1(new_n1103), .B2(new_n1097), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  XOR2_X1   g680(.A(KEYINPUT58), .B(G1341), .Z(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(new_n1000), .B2(new_n1037), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(new_n1082), .B2(G1996), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1108), .A2(KEYINPUT59), .A3(new_n563), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT59), .B1(new_n1108), .B2(new_n563), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1104), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1112), .A2(KEYINPUT61), .A3(new_n1099), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1114), .B1(new_n1100), .B2(new_n1104), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n1090), .A2(KEYINPUT122), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n633), .A2(KEYINPUT60), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1116), .A2(new_n1092), .A3(new_n1089), .A4(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1111), .A2(new_n1113), .A3(new_n1115), .A4(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT60), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1116), .A2(new_n633), .A3(new_n1092), .A4(new_n1089), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1120), .B1(new_n1094), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1105), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n816), .B1(new_n1000), .B2(new_n1064), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(KEYINPUT123), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT123), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1126), .B(new_n816), .C1(new_n1000), .C2(new_n1064), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT53), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1129), .A2(G2078), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n998), .A2(G40), .A3(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1131), .A2(new_n483), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1132), .A2(new_n1068), .A3(new_n1004), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1129), .B1(new_n1082), .B2(G2078), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1128), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1135), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT125), .B1(new_n1135), .B2(G171), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1030), .A2(KEYINPUT45), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1029), .A2(new_n1081), .A3(new_n1138), .A4(new_n1130), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1134), .A2(new_n1124), .A3(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT54), .B1(new_n1140), .B2(G171), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1137), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT118), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1143), .B1(new_n1088), .B2(G2084), .ZN(new_n1144));
  NAND4_X1  g719(.A1(G160), .A2(new_n1081), .A3(G40), .A4(new_n1138), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n765), .ZN(new_n1146));
  INV_X1    g721(.A(G2084), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1083), .A2(KEYINPUT118), .A3(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1144), .A2(G168), .A3(new_n1146), .A4(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(G8), .ZN(new_n1150));
  AOI21_X1  g725(.A(KEYINPUT118), .B1(new_n1083), .B2(new_n1147), .ZN(new_n1151));
  NOR4_X1   g726(.A1(new_n1000), .A2(new_n1064), .A3(new_n1143), .A4(G2084), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(G168), .B1(new_n1153), .B2(new_n1146), .ZN(new_n1154));
  OAI21_X1  g729(.A(KEYINPUT51), .B1(new_n1150), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT51), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1149), .A2(new_n1156), .A3(G8), .ZN(new_n1157));
  AOI22_X1  g732(.A1(new_n1136), .A2(new_n1142), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT54), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1140), .A2(G171), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1128), .A2(new_n1133), .A3(new_n1134), .A4(G301), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT124), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  AND2_X1   g738(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1159), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1123), .A2(new_n1158), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(KEYINPUT62), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1160), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT62), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1155), .A2(new_n1170), .A3(new_n1157), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1168), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1087), .B1(new_n1166), .B2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1085), .B1(new_n1073), .B2(KEYINPUT114), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1076), .B1(new_n1174), .B2(new_n1078), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1176), .A2(new_n1039), .A3(new_n1036), .ZN(new_n1177));
  OAI21_X1  g752(.A(KEYINPUT119), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n638), .A2(G8), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1179), .B1(new_n1153), .B2(new_n1146), .ZN(new_n1180));
  AND3_X1   g755(.A1(new_n1079), .A2(KEYINPUT63), .A3(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(G8), .B1(new_n1084), .B2(new_n1077), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1078), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1080), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT119), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1184), .A2(new_n1059), .A3(new_n1185), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1178), .A2(new_n1181), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1187), .A2(KEYINPUT120), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT120), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1178), .A2(new_n1181), .A3(new_n1186), .A4(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT63), .ZN(new_n1191));
  INV_X1    g766(.A(new_n1180), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1191), .B1(new_n1087), .B2(new_n1192), .ZN(new_n1193));
  AND3_X1   g768(.A1(new_n1188), .A2(new_n1190), .A3(new_n1193), .ZN(new_n1194));
  NOR2_X1   g769(.A1(G288), .A2(G1976), .ZN(new_n1195));
  AOI22_X1  g770(.A1(new_n1176), .A2(new_n1195), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1196));
  OAI22_X1  g771(.A1(new_n1196), .A2(new_n1038), .B1(new_n1177), .B2(new_n1079), .ZN(new_n1197));
  NOR3_X1   g772(.A1(new_n1173), .A2(new_n1194), .A3(new_n1197), .ZN(new_n1198));
  XOR2_X1   g773(.A(G290), .B(G1986), .Z(new_n1199));
  OAI21_X1  g774(.A(new_n1024), .B1(new_n1006), .B2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1028), .B1(new_n1198), .B2(new_n1200), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g776(.A1(new_n899), .A2(new_n903), .ZN(new_n1203));
  NAND2_X1  g777(.A1(new_n984), .A2(new_n985), .ZN(new_n1204));
  NAND2_X1  g778(.A1(new_n689), .A2(G319), .ZN(new_n1205));
  NOR3_X1   g779(.A1(G229), .A2(G401), .A3(new_n1205), .ZN(new_n1206));
  NAND3_X1  g780(.A1(new_n1203), .A2(new_n1204), .A3(new_n1206), .ZN(G225));
  INV_X1    g781(.A(G225), .ZN(G308));
endmodule


