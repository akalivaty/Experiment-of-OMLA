//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 1 0 0 1 0 1 0 0 1 0 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 1 1 1 1 1 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  OR2_X1    g003(.A1(KEYINPUT75), .A2(KEYINPUT25), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NOR3_X1   g005(.A1(new_n191), .A2(KEYINPUT16), .A3(G140), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G140), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G125), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n191), .A2(G140), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT16), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n193), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(G125), .B(G140), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n192), .B1(new_n202), .B2(KEYINPUT16), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n206));
  INV_X1    g020(.A(G119), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G128), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(KEYINPUT23), .A3(G119), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n208), .B(new_n210), .C1(G119), .C2(new_n209), .ZN(new_n211));
  XNOR2_X1  g025(.A(G119), .B(G128), .ZN(new_n212));
  XOR2_X1   g026(.A(KEYINPUT24), .B(G110), .Z(new_n213));
  AOI22_X1  g027(.A1(new_n211), .A2(G110), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n205), .A2(new_n214), .ZN(new_n215));
  OAI22_X1  g029(.A1(new_n211), .A2(G110), .B1(new_n212), .B2(new_n213), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n202), .A2(new_n200), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n217), .A3(new_n204), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT22), .B(G137), .ZN(new_n220));
  INV_X1    g034(.A(G953), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(G221), .A3(G234), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n220), .B(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n215), .A2(new_n218), .A3(new_n223), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n190), .B1(new_n227), .B2(new_n188), .ZN(new_n228));
  AND4_X1   g042(.A1(new_n188), .A2(new_n225), .A3(new_n226), .A4(new_n190), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n189), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n189), .A2(G902), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n234));
  NAND2_X1  g048(.A1(KEYINPUT11), .A2(G134), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n234), .B1(new_n235), .B2(G137), .ZN(new_n236));
  INV_X1    g050(.A(G137), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n237), .A2(KEYINPUT69), .A3(KEYINPUT11), .A4(G134), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  OR2_X1    g053(.A1(KEYINPUT68), .A2(G134), .ZN(new_n240));
  NAND2_X1  g054(.A1(KEYINPUT68), .A2(G134), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n240), .A2(G137), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(G137), .B1(new_n240), .B2(new_n241), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n239), .B(new_n242), .C1(new_n243), .C2(KEYINPUT11), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G131), .ZN(new_n245));
  AND2_X1   g059(.A1(KEYINPUT68), .A2(G134), .ZN(new_n246));
  NOR2_X1   g060(.A1(KEYINPUT68), .A2(G134), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n237), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT11), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT70), .B(G131), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n250), .A2(new_n251), .A3(new_n239), .A4(new_n242), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n245), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n200), .A2(G143), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(KEYINPUT0), .A2(G128), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT66), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n258), .B1(G143), .B2(new_n200), .ZN(new_n259));
  INV_X1    g073(.A(G143), .ZN(new_n260));
  NOR3_X1   g074(.A1(new_n260), .A2(KEYINPUT66), .A3(G146), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n255), .B(new_n257), .C1(new_n259), .C2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n200), .A2(G143), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT65), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n265), .B1(new_n200), .B2(G143), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n260), .A2(KEYINPUT65), .A3(G146), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n264), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n269));
  NOR2_X1   g083(.A1(KEYINPUT0), .A2(G128), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AND3_X1   g085(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n262), .B1(new_n268), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n253), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT2), .ZN(new_n278));
  INV_X1    g092(.A(G113), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n278), .A2(new_n279), .A3(KEYINPUT71), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n281), .B1(KEYINPUT2), .B2(G113), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(KEYINPUT2), .A2(G113), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n207), .A2(G116), .ZN(new_n286));
  INV_X1    g100(.A(G116), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G119), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n280), .A2(new_n282), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT72), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n286), .A2(new_n288), .A3(new_n284), .ZN(new_n293));
  NOR3_X1   g107(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n286), .A2(new_n288), .A3(new_n284), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT72), .B1(new_n295), .B2(new_n283), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n290), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n209), .A2(KEYINPUT1), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n255), .B(new_n299), .C1(new_n259), .C2(new_n261), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n209), .B1(new_n263), .B2(KEYINPUT1), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n300), .B1(new_n268), .B2(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n237), .A2(G134), .ZN(new_n303));
  OAI21_X1  g117(.A(G131), .B1(new_n243), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n302), .A2(new_n252), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n277), .A2(new_n298), .A3(new_n305), .ZN(new_n306));
  XOR2_X1   g120(.A(KEYINPUT73), .B(KEYINPUT27), .Z(new_n307));
  NOR2_X1   g121(.A1(G237), .A2(G953), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G210), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n307), .B(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT26), .B(G101), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n310), .B(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n306), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n275), .A2(KEYINPUT67), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT67), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n262), .B(new_n315), .C1(new_n268), .C2(new_n274), .ZN(new_n316));
  INV_X1    g130(.A(G131), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n246), .A2(new_n247), .A3(new_n237), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n318), .B1(new_n249), .B2(new_n248), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n317), .B1(new_n319), .B2(new_n239), .ZN(new_n320));
  INV_X1    g134(.A(new_n252), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n314), .B(new_n316), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(KEYINPUT30), .B1(new_n322), .B2(new_n305), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n275), .B1(new_n245), .B2(new_n252), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n302), .A2(new_n252), .A3(new_n304), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT30), .ZN(new_n326));
  NOR3_X1   g140(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n313), .B1(new_n328), .B2(new_n297), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT31), .ZN(new_n330));
  INV_X1    g144(.A(new_n312), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n298), .B1(new_n322), .B2(new_n305), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT28), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n324), .A2(new_n325), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n334), .B1(new_n335), .B2(new_n298), .ZN(new_n336));
  NOR4_X1   g150(.A1(new_n324), .A2(new_n325), .A3(KEYINPUT28), .A4(new_n297), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n333), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AOI22_X1  g152(.A1(new_n329), .A2(new_n330), .B1(new_n331), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT74), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n277), .A2(KEYINPUT30), .A3(new_n305), .ZN(new_n341));
  INV_X1    g155(.A(new_n316), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n260), .A2(KEYINPUT65), .A3(G146), .ZN(new_n343));
  AOI21_X1  g157(.A(KEYINPUT65), .B1(new_n260), .B2(G146), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n263), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n272), .A2(new_n269), .A3(new_n270), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n315), .B1(new_n347), .B2(new_n262), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n342), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n325), .B1(new_n349), .B2(new_n253), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n297), .B(new_n341), .C1(new_n350), .C2(KEYINPUT30), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n331), .B1(new_n298), .B2(new_n335), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n340), .B1(new_n353), .B2(KEYINPUT31), .ZN(new_n354));
  AOI211_X1 g168(.A(KEYINPUT74), .B(new_n330), .C1(new_n351), .C2(new_n352), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n339), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(G472), .A2(G902), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT32), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n297), .B1(new_n324), .B2(new_n325), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT29), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n331), .A2(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n361), .B(new_n363), .C1(new_n336), .C2(new_n337), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n188), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n306), .A2(new_n331), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  AOI22_X1  g182(.A1(new_n338), .A2(new_n312), .B1(new_n368), .B2(new_n351), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n366), .B1(new_n369), .B2(KEYINPUT29), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n356), .A2(new_n360), .B1(new_n370), .B2(G472), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n351), .A2(new_n330), .A3(new_n352), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n306), .A2(KEYINPUT28), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n335), .A2(new_n334), .A3(new_n298), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n332), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n372), .B1(new_n312), .B2(new_n375), .ZN(new_n376));
  NOR3_X1   g190(.A1(new_n323), .A2(new_n327), .A3(new_n298), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT31), .B1(new_n377), .B2(new_n313), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(KEYINPUT74), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n353), .A2(new_n340), .A3(KEYINPUT31), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n376), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n359), .B1(new_n381), .B2(new_n358), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n233), .B1(new_n371), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(G214), .B1(G237), .B2(G902), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n221), .A2(G952), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n386), .B1(G234), .B2(G237), .ZN(new_n387));
  XOR2_X1   g201(.A(KEYINPUT21), .B(G898), .Z(new_n388));
  XNOR2_X1  g202(.A(new_n388), .B(KEYINPUT94), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  AOI211_X1 g204(.A(new_n188), .B(new_n221), .C1(G234), .C2(G237), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n387), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n292), .B1(new_n291), .B2(new_n293), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n295), .A2(KEYINPUT72), .A3(new_n283), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G104), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n396), .A2(G107), .ZN(new_n397));
  INV_X1    g211(.A(G107), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(G104), .ZN(new_n399));
  OAI21_X1  g213(.A(G101), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT3), .B1(new_n396), .B2(G107), .ZN(new_n401));
  AOI21_X1  g215(.A(G101), .B1(new_n396), .B2(G107), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT3), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(new_n398), .A3(G104), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n401), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n400), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n286), .A2(new_n288), .A3(KEYINPUT5), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n408), .B(G113), .C1(KEYINPUT5), .C2(new_n286), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n395), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n396), .A2(G107), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n401), .A2(new_n404), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G101), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(KEYINPUT4), .A3(new_n405), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(KEYINPUT76), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT76), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n405), .A2(KEYINPUT4), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n416), .B1(new_n417), .B2(new_n413), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n413), .A2(KEYINPUT4), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n297), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n410), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT6), .ZN(new_n424));
  XNOR2_X1  g238(.A(G110), .B(G122), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n425), .B(KEYINPUT78), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n423), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n426), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n428), .B(new_n410), .C1(new_n419), .C2(new_n422), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT6), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n414), .A2(KEYINPUT76), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n417), .A2(new_n416), .A3(new_n413), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(new_n297), .A3(new_n421), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n428), .B1(new_n434), .B2(new_n410), .ZN(new_n435));
  OAI211_X1 g249(.A(KEYINPUT79), .B(new_n427), .C1(new_n430), .C2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n423), .A2(new_n426), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT79), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n437), .A2(new_n438), .A3(KEYINPUT6), .A4(new_n429), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n275), .A2(G125), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n300), .B(new_n191), .C1(new_n268), .C2(new_n301), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n221), .A2(G224), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n443), .B(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n440), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(G210), .B1(G237), .B2(G902), .ZN(new_n448));
  XOR2_X1   g262(.A(new_n426), .B(KEYINPUT8), .Z(new_n449));
  INV_X1    g263(.A(new_n410), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n407), .B1(new_n395), .B2(new_n409), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n444), .A2(KEYINPUT7), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n442), .A2(KEYINPUT80), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n441), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n442), .A2(KEYINPUT80), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n453), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT81), .ZN(new_n458));
  OAI21_X1  g272(.A(KEYINPUT7), .B1(new_n444), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n459), .B1(new_n458), .B2(new_n444), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n441), .A2(new_n442), .A3(new_n460), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n452), .A2(new_n457), .A3(KEYINPUT82), .A4(new_n461), .ZN(new_n462));
  AND2_X1   g276(.A1(new_n462), .A2(new_n429), .ZN(new_n463));
  INV_X1    g277(.A(new_n461), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n395), .A2(new_n409), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n406), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n410), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n464), .B1(new_n467), .B2(new_n449), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n457), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT82), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(G902), .B1(new_n463), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n447), .A2(new_n448), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n448), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n445), .B1(new_n436), .B2(new_n439), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n462), .A2(new_n429), .ZN(new_n476));
  AOI21_X1  g290(.A(KEYINPUT82), .B1(new_n468), .B2(new_n457), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n188), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n474), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  AOI211_X1 g293(.A(new_n385), .B(new_n392), .C1(new_n473), .C2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT13), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n481), .B1(new_n209), .B2(G143), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n260), .A2(KEYINPUT13), .A3(G128), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n209), .A2(G143), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n482), .A2(new_n483), .A3(KEYINPUT90), .A4(new_n484), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n485), .B(G134), .C1(KEYINPUT90), .C2(new_n483), .ZN(new_n486));
  XOR2_X1   g300(.A(G116), .B(G122), .Z(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(G107), .ZN(new_n488));
  XNOR2_X1  g302(.A(G116), .B(G122), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n398), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n240), .A2(new_n241), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n260), .A2(G128), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n484), .ZN(new_n494));
  OR2_X1    g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n486), .A2(new_n491), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT91), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n486), .A2(new_n491), .A3(KEYINPUT91), .A4(new_n495), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n492), .B(new_n494), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n287), .A2(KEYINPUT14), .A3(G122), .ZN(new_n501));
  OAI211_X1 g315(.A(G107), .B(new_n501), .C1(new_n487), .C2(KEYINPUT14), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n500), .A2(new_n490), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n498), .A2(new_n499), .A3(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(KEYINPUT9), .B(G234), .ZN(new_n505));
  NOR3_X1   g319(.A1(new_n505), .A2(new_n187), .A3(G953), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(KEYINPUT92), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n498), .A2(new_n507), .A3(new_n499), .A4(new_n503), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(new_n188), .A3(new_n510), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n511), .A2(KEYINPUT93), .ZN(new_n512));
  INV_X1    g326(.A(G478), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n513), .A2(KEYINPUT15), .ZN(new_n514));
  OR2_X1    g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n511), .A2(KEYINPUT93), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n514), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  XOR2_X1   g332(.A(KEYINPUT70), .B(G131), .Z(new_n519));
  AND3_X1   g333(.A1(new_n308), .A2(G143), .A3(G214), .ZN(new_n520));
  AOI21_X1  g334(.A(G143), .B1(new_n308), .B2(G214), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT17), .ZN(new_n523));
  INV_X1    g337(.A(G237), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n524), .A2(new_n221), .A3(G214), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n260), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n308), .A2(G143), .A3(G214), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n526), .A2(new_n527), .A3(new_n251), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n522), .A2(new_n523), .A3(new_n528), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n519), .B(KEYINPUT17), .C1(new_n520), .C2(new_n521), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n529), .A2(new_n201), .A3(new_n204), .A4(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(KEYINPUT83), .B1(new_n526), .B2(new_n527), .ZN(new_n532));
  AND2_X1   g346(.A1(KEYINPUT18), .A2(G131), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT84), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n197), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n202), .A2(KEYINPUT84), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n536), .A2(new_n537), .A3(KEYINPUT85), .A4(G146), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n195), .A2(new_n196), .A3(KEYINPUT84), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT84), .B1(new_n195), .B2(new_n196), .ZN(new_n540));
  NOR3_X1   g354(.A1(new_n539), .A2(new_n540), .A3(new_n200), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT85), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n217), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n534), .B(new_n538), .C1(new_n541), .C2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n526), .A2(KEYINPUT83), .A3(new_n527), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n532), .B1(new_n545), .B2(new_n533), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n531), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  XOR2_X1   g361(.A(G113), .B(G122), .Z(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT87), .B(G104), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n548), .B(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT89), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n188), .B1(new_n547), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n545), .A2(new_n533), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n520), .A2(new_n521), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n555), .B1(KEYINPUT83), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n536), .A2(new_n537), .A3(G146), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n558), .A2(new_n542), .A3(new_n217), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n557), .A2(new_n559), .A3(new_n534), .A4(new_n538), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n552), .B1(new_n560), .B2(new_n531), .ZN(new_n561));
  OAI21_X1  g375(.A(G475), .B1(new_n554), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n547), .A2(new_n550), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT88), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n536), .A2(new_n537), .A3(KEYINPUT19), .ZN(new_n565));
  OR3_X1    g379(.A1(new_n197), .A2(KEYINPUT86), .A3(KEYINPUT19), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT86), .B1(new_n197), .B2(KEYINPUT19), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n565), .A2(new_n566), .A3(new_n200), .A4(new_n567), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n522), .A2(new_n528), .B1(new_n203), .B2(G146), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n550), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n560), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n563), .A2(new_n564), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT20), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n547), .A2(new_n550), .B1(new_n560), .B2(new_n570), .ZN(new_n574));
  NOR2_X1   g388(.A1(G475), .A2(G902), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n572), .A2(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AND4_X1   g390(.A1(KEYINPUT88), .A2(new_n574), .A3(new_n573), .A4(new_n575), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n562), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n518), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(G469), .ZN(new_n580));
  XNOR2_X1  g394(.A(G110), .B(G140), .ZN(new_n581));
  INV_X1    g395(.A(G227), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n582), .A2(G953), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n581), .B(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n420), .A2(new_n275), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n433), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT77), .ZN(new_n588));
  INV_X1    g402(.A(new_n301), .ZN(new_n589));
  OAI21_X1  g403(.A(KEYINPUT66), .B1(new_n260), .B2(G146), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n258), .A2(new_n200), .A3(G143), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n254), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g406(.A1(new_n345), .A2(new_n589), .B1(new_n592), .B2(new_n299), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n400), .A2(new_n405), .A3(KEYINPUT10), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n588), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n302), .A2(new_n407), .A3(KEYINPUT77), .A4(KEYINPUT10), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n255), .B1(new_n259), .B2(new_n261), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n589), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n300), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT10), .B1(new_n600), .B2(new_n407), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n587), .A2(new_n597), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n253), .ZN(new_n604));
  INV_X1    g418(.A(new_n253), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n587), .A2(new_n605), .A3(new_n597), .A4(new_n602), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n585), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n302), .A2(new_n407), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n406), .B1(new_n599), .B2(new_n300), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n253), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(KEYINPUT12), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT12), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n253), .B(new_n612), .C1(new_n608), .C2(new_n609), .ZN(new_n613));
  AND4_X1   g427(.A1(new_n606), .A2(new_n585), .A3(new_n611), .A4(new_n613), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n580), .B(new_n188), .C1(new_n607), .C2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n580), .A2(new_n188), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n606), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n611), .A2(new_n613), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n584), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n604), .A2(new_n606), .A3(new_n585), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n620), .A2(G469), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n615), .A2(new_n617), .A3(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(G221), .B1(new_n505), .B2(G902), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n383), .A2(new_n480), .A3(new_n579), .A4(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT95), .B(G101), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G3));
  INV_X1    g442(.A(G472), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n629), .B1(new_n356), .B2(new_n188), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n381), .A2(new_n358), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n233), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n633), .A2(new_n624), .A3(new_n623), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(new_n635), .B(KEYINPUT96), .Z(new_n636));
  NOR2_X1   g450(.A1(new_n513), .A2(G902), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n509), .A2(KEYINPUT33), .A3(new_n510), .ZN(new_n638));
  AOI21_X1  g452(.A(KEYINPUT33), .B1(new_n509), .B2(new_n510), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT97), .B(G478), .Z(new_n641));
  NAND2_X1  g455(.A1(new_n511), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n578), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n480), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n636), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT34), .B(G104), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G6));
  NAND2_X1  g464(.A1(new_n574), .A2(new_n575), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT20), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n562), .A2(KEYINPUT98), .ZN(new_n653));
  OR2_X1    g467(.A1(new_n562), .A2(KEYINPUT98), .ZN(new_n654));
  AND4_X1   g468(.A1(new_n518), .A2(new_n652), .A3(new_n653), .A4(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n636), .A2(new_n480), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT35), .B(G107), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G9));
  NOR2_X1   g472(.A1(new_n224), .A2(KEYINPUT36), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n219), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n231), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n230), .A2(new_n661), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n623), .A2(new_n624), .A3(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n480), .A2(new_n632), .A3(new_n579), .A4(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT37), .B(G110), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G12));
  INV_X1    g480(.A(new_n360), .ZN(new_n667));
  OAI22_X1  g481(.A1(new_n375), .A2(new_n331), .B1(new_n377), .B2(new_n367), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n365), .B1(new_n668), .B2(new_n362), .ZN(new_n669));
  OAI22_X1  g483(.A1(new_n381), .A2(new_n667), .B1(new_n629), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(KEYINPUT32), .B1(new_n356), .B2(new_n357), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n663), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n385), .B1(new_n473), .B2(new_n479), .ZN(new_n674));
  INV_X1    g488(.A(new_n518), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n387), .B(KEYINPUT99), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(G900), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n677), .B1(new_n678), .B2(new_n391), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n652), .A2(new_n653), .A3(new_n654), .A4(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n675), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n674), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n673), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G128), .ZN(G30));
  NAND2_X1  g500(.A1(new_n473), .A2(new_n479), .ZN(new_n687));
  XOR2_X1   g501(.A(new_n687), .B(KEYINPUT38), .Z(new_n688));
  AND2_X1   g502(.A1(new_n518), .A2(new_n578), .ZN(new_n689));
  INV_X1    g503(.A(new_n662), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n689), .A2(new_n384), .A3(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(new_n679), .B(KEYINPUT39), .Z(new_n693));
  NAND2_X1  g507(.A1(new_n625), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT40), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n368), .A2(new_n361), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n188), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n331), .B1(new_n351), .B2(new_n306), .ZN(new_n699));
  OAI21_X1  g513(.A(G472), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n700), .B(KEYINPUT100), .Z(new_n701));
  NAND2_X1  g515(.A1(new_n356), .A2(new_n360), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n701), .A2(new_n382), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n692), .A2(new_n696), .A3(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT101), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n692), .A2(new_n696), .A3(KEYINPUT101), .A4(new_n703), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G143), .ZN(G45));
  NAND3_X1  g523(.A1(new_n578), .A2(new_n643), .A3(new_n680), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n674), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(KEYINPUT102), .B1(new_n672), .B2(new_n712), .ZN(new_n713));
  AOI211_X1 g527(.A(new_n385), .B(new_n710), .C1(new_n473), .C2(new_n479), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n371), .A2(new_n382), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT102), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n714), .A2(new_n715), .A3(new_n716), .A4(new_n663), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G146), .ZN(G48));
  OAI21_X1  g533(.A(new_n188), .B1(new_n607), .B2(new_n614), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(G469), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n721), .A2(new_n624), .A3(new_n615), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n715), .A2(new_n633), .A3(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n646), .ZN(new_n724));
  XOR2_X1   g538(.A(KEYINPUT41), .B(G113), .Z(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G15));
  NAND2_X1  g540(.A1(new_n480), .A2(new_n655), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(new_n287), .ZN(G18));
  NOR2_X1   g543(.A1(new_n690), .A2(new_n392), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n579), .B(new_n730), .C1(new_n670), .C2(new_n671), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n674), .A2(new_n722), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT103), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n674), .A2(KEYINPUT103), .A3(new_n722), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n731), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(new_n207), .ZN(G21));
  INV_X1    g551(.A(new_n630), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n361), .B1(new_n336), .B2(new_n337), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n331), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n378), .A2(new_n740), .A3(new_n372), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n357), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT104), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n741), .A2(KEYINPUT104), .A3(new_n357), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n738), .A2(new_n633), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n392), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n674), .A2(new_n747), .A3(new_n689), .A4(new_n722), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  XOR2_X1   g563(.A(new_n749), .B(G122), .Z(G24));
  NAND2_X1  g564(.A1(new_n744), .A2(new_n745), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n751), .A2(new_n630), .A3(new_n690), .ZN(new_n752));
  AND4_X1   g566(.A1(KEYINPUT103), .A2(new_n687), .A3(new_n722), .A4(new_n384), .ZN(new_n753));
  AOI21_X1  g567(.A(KEYINPUT103), .B1(new_n674), .B2(new_n722), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n711), .B(new_n752), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G125), .ZN(G27));
  NAND2_X1  g570(.A1(new_n382), .A2(new_n702), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT107), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n370), .A2(G472), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT107), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n382), .A2(new_n760), .A3(new_n702), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n758), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT105), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n763), .B1(new_n620), .B2(new_n621), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n621), .A2(new_n763), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n764), .A2(new_n765), .A3(new_n580), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n615), .A2(new_n617), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n624), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n473), .A2(new_n384), .A3(new_n479), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT42), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n710), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n762), .A2(new_n633), .A3(new_n770), .A4(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n383), .A2(new_n770), .A3(new_n711), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT106), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n383), .A2(new_n770), .A3(KEYINPUT106), .A4(new_n711), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n771), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n773), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G131), .ZN(G33));
  NAND3_X1  g594(.A1(new_n383), .A2(new_n770), .A3(new_n682), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G134), .ZN(G36));
  INV_X1    g596(.A(KEYINPUT45), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n764), .A2(new_n765), .A3(new_n783), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n620), .A2(new_n621), .ZN(new_n785));
  OAI21_X1  g599(.A(G469), .B1(new_n785), .B2(KEYINPUT45), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(new_n616), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n788), .A2(KEYINPUT46), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n615), .B1(new_n788), .B2(KEYINPUT46), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n624), .B(new_n693), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT108), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n791), .B(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n578), .B1(new_n640), .B2(new_n642), .ZN(new_n794));
  AND2_X1   g608(.A1(KEYINPUT109), .A2(KEYINPUT43), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(KEYINPUT109), .A2(KEYINPUT43), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n794), .B1(new_n797), .B2(new_n795), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT110), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n632), .A2(new_n690), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n796), .A2(KEYINPUT110), .A3(new_n798), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT44), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n806), .A2(new_n807), .A3(new_n769), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n793), .A2(new_n808), .ZN(new_n809));
  XOR2_X1   g623(.A(KEYINPUT111), .B(G137), .Z(new_n810));
  XNOR2_X1  g624(.A(new_n809), .B(new_n810), .ZN(G39));
  OR4_X1    g625(.A1(new_n715), .A2(new_n633), .A3(new_n710), .A4(new_n769), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n624), .B1(new_n789), .B2(new_n790), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT47), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI211_X1 g629(.A(KEYINPUT47), .B(new_n624), .C1(new_n789), .C2(new_n790), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n812), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(new_n194), .ZN(G42));
  OAI22_X1  g632(.A1(new_n723), .A2(new_n646), .B1(new_n746), .B2(new_n748), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n819), .A2(new_n736), .A3(new_n728), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n644), .B1(new_n675), .B2(new_n578), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n480), .A2(new_n632), .A3(new_n634), .A4(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n626), .A2(new_n664), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n751), .A2(new_n630), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n770), .A2(new_n824), .A3(new_n662), .A4(new_n711), .ZN(new_n825));
  INV_X1    g639(.A(new_n769), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n518), .A2(new_n681), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n715), .A2(new_n826), .A3(new_n663), .A4(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n825), .A2(new_n781), .A3(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n823), .A2(new_n829), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n779), .A2(new_n820), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(KEYINPUT112), .B1(new_n662), .B2(new_n679), .ZN(new_n832));
  OR3_X1    g646(.A1(new_n662), .A2(KEYINPUT112), .A3(new_n679), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n768), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n674), .A2(new_n689), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n703), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n718), .A2(new_n685), .A3(new_n755), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT52), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n734), .A2(new_n735), .ZN(new_n839));
  NOR4_X1   g653(.A1(new_n751), .A2(new_n630), .A3(new_n690), .A4(new_n710), .ZN(new_n840));
  AOI22_X1  g654(.A1(new_n839), .A2(new_n840), .B1(new_n673), .B2(new_n684), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT52), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n841), .A2(new_n842), .A3(new_n718), .A4(new_n836), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n755), .A2(new_n685), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n844), .B1(new_n845), .B2(KEYINPUT52), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n831), .A2(new_n838), .A3(new_n843), .A4(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n838), .A2(new_n843), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n779), .A2(new_n820), .A3(new_n830), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n844), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n851), .A2(KEYINPUT54), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n838), .A2(new_n843), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n845), .A2(KEYINPUT52), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n844), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n854), .A2(new_n831), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n853), .B1(new_n857), .B2(new_n850), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n852), .A2(new_n858), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n826), .A2(new_n722), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n676), .B1(new_n796), .B2(new_n798), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XOR2_X1   g676(.A(new_n862), .B(KEYINPUT115), .Z(new_n863));
  AND2_X1   g677(.A1(new_n762), .A2(new_n633), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT48), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n861), .A2(new_n633), .A3(new_n824), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n867), .B1(new_n734), .B2(new_n735), .ZN(new_n868));
  INV_X1    g682(.A(new_n703), .ZN(new_n869));
  AND4_X1   g683(.A1(new_n387), .A2(new_n869), .A3(new_n633), .A4(new_n860), .ZN(new_n870));
  AOI211_X1 g684(.A(new_n386), .B(new_n868), .C1(new_n870), .C2(new_n645), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n866), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n578), .A2(new_n643), .ZN(new_n873));
  AOI22_X1  g687(.A1(new_n863), .A2(new_n752), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n688), .A2(new_n385), .A3(new_n722), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n867), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT50), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n878), .A2(KEYINPUT51), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n867), .A2(new_n769), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n815), .A2(new_n816), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n721), .A2(new_n615), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n882), .A2(new_n624), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n880), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n872), .B1(new_n879), .B2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT113), .ZN(new_n886));
  OAI22_X1  g700(.A1(new_n881), .A2(new_n886), .B1(new_n624), .B2(new_n882), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT113), .B1(new_n815), .B2(new_n816), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n880), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OR2_X1    g703(.A1(new_n889), .A2(KEYINPUT114), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(KEYINPUT114), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n890), .A2(new_n878), .A3(new_n891), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n859), .B(new_n885), .C1(new_n892), .C2(KEYINPUT51), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n893), .B1(G952), .B2(G953), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n882), .A2(KEYINPUT49), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n794), .A2(new_n633), .A3(new_n384), .A4(new_n624), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n882), .A2(KEYINPUT49), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n688), .A2(new_n869), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n894), .A2(new_n899), .ZN(G75));
  AND2_X1   g714(.A1(new_n847), .A2(new_n850), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n901), .A2(new_n188), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(G210), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n440), .A2(new_n446), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n904), .A2(new_n475), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT55), .ZN(new_n906));
  XOR2_X1   g720(.A(KEYINPUT116), .B(KEYINPUT56), .Z(new_n907));
  AND3_X1   g721(.A1(new_n903), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT56), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n906), .B1(new_n903), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n221), .A2(G952), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n908), .A2(new_n910), .A3(new_n911), .ZN(G51));
  NAND2_X1  g726(.A1(new_n901), .A2(new_n853), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT117), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n851), .A2(KEYINPUT54), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n851), .A2(KEYINPUT117), .A3(KEYINPUT54), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n616), .B(KEYINPUT57), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(new_n607), .B2(new_n614), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n902), .A2(new_n787), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n911), .B1(new_n920), .B2(new_n921), .ZN(G54));
  NAND3_X1  g736(.A1(new_n902), .A2(KEYINPUT58), .A3(G475), .ZN(new_n923));
  INV_X1    g737(.A(new_n574), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n923), .A2(new_n924), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n925), .A2(new_n926), .A3(new_n911), .ZN(G60));
  OR2_X1    g741(.A1(new_n638), .A2(new_n639), .ZN(new_n928));
  NAND2_X1  g742(.A1(G478), .A2(G902), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT59), .Z(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n916), .A2(new_n928), .A3(new_n917), .A4(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n911), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n931), .B1(new_n852), .B2(new_n858), .ZN(new_n935));
  INV_X1    g749(.A(new_n928), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT118), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n935), .A2(KEYINPUT118), .A3(new_n936), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n934), .A2(new_n937), .A3(new_n938), .ZN(G63));
  XNOR2_X1  g753(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n940));
  NAND2_X1  g754(.A1(G217), .A2(G902), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT60), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(KEYINPUT119), .B1(new_n851), .B2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT119), .ZN(new_n945));
  AOI211_X1 g759(.A(new_n945), .B(new_n942), .C1(new_n847), .C2(new_n850), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n227), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n911), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n660), .B1(new_n944), .B2(new_n946), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n940), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n945), .B1(new_n901), .B2(new_n942), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n851), .A2(KEYINPUT119), .A3(new_n943), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n952), .A2(new_n948), .A3(new_n953), .ZN(new_n954));
  AND4_X1   g768(.A1(new_n933), .A2(new_n954), .A3(new_n950), .A4(new_n940), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n951), .A2(new_n955), .ZN(G66));
  INV_X1    g770(.A(G224), .ZN(new_n957));
  OAI21_X1  g771(.A(G953), .B1(new_n390), .B2(new_n957), .ZN(new_n958));
  NOR4_X1   g772(.A1(new_n823), .A2(new_n819), .A3(new_n736), .A4(new_n728), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n958), .B1(new_n959), .B2(G953), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n436), .B(new_n439), .C1(G898), .C2(new_n221), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(G69));
  NAND3_X1  g776(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n328), .B(new_n963), .Z(new_n964));
  AOI21_X1  g778(.A(new_n817), .B1(new_n793), .B2(new_n808), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n841), .A2(new_n718), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n793), .A2(new_n835), .A3(new_n864), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n779), .A2(new_n781), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT124), .Z(new_n970));
  AOI21_X1  g784(.A(G953), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n221), .A2(G900), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n964), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n966), .A2(new_n706), .A3(new_n707), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(KEYINPUT62), .ZN(new_n975));
  INV_X1    g789(.A(new_n694), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n976), .A2(new_n383), .A3(new_n826), .A4(new_n821), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n975), .A2(new_n965), .A3(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT122), .ZN(new_n979));
  OAI21_X1  g793(.A(KEYINPUT121), .B1(new_n974), .B2(KEYINPUT62), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT121), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT62), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n708), .A2(new_n981), .A3(new_n982), .A4(new_n966), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n978), .A2(new_n979), .A3(new_n980), .A4(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n980), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n975), .A2(new_n965), .A3(new_n977), .ZN(new_n986));
  OAI21_X1  g800(.A(KEYINPUT122), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(G953), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n973), .B1(new_n988), .B2(new_n964), .ZN(new_n989));
  OAI21_X1  g803(.A(G953), .B1(new_n582), .B2(new_n678), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT123), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(new_n991), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n973), .B(new_n993), .C1(new_n988), .C2(new_n964), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n992), .A2(new_n994), .ZN(G72));
  NOR2_X1   g809(.A1(new_n377), .A2(new_n367), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n968), .A2(new_n959), .A3(new_n970), .ZN(new_n998));
  NAND2_X1  g812(.A1(G472), .A2(G902), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT63), .Z(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT125), .Z(new_n1001));
  AOI21_X1  g815(.A(new_n997), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n857), .A2(new_n850), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT127), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1000), .ZN(new_n1005));
  NOR3_X1   g819(.A1(new_n996), .A2(new_n699), .A3(new_n1005), .ZN(new_n1006));
  XOR2_X1   g820(.A(new_n1006), .B(KEYINPUT126), .Z(new_n1007));
  AND3_X1   g821(.A1(new_n1003), .A2(new_n1004), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1004), .B1(new_n1003), .B2(new_n1007), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n933), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n984), .A2(new_n987), .A3(new_n959), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(new_n1001), .ZN(new_n1012));
  AOI211_X1 g826(.A(new_n1002), .B(new_n1010), .C1(new_n1012), .C2(new_n699), .ZN(G57));
endmodule


