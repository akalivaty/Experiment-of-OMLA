//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0 1 0 0 1 0 0 0 1 1 0 0 1 1 0 0 0 0 1 1 1 1 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n569, new_n571,
    new_n572, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1163, new_n1164, new_n1165;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  XNOR2_X1  g031(.A(KEYINPUT3), .B(G2104), .ZN(new_n457));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G137), .ZN(new_n461));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n463), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  AND3_X1   g047(.A1(new_n461), .A2(new_n470), .A3(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n460), .A2(G136), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n467), .A2(new_n458), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  OR2_X1    g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n477), .B(G2104), .C1(G112), .C2(new_n458), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n474), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G162));
  INV_X1    g055(.A(KEYINPUT70), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT67), .ZN(new_n484));
  OAI21_X1  g059(.A(G2105), .B1(new_n484), .B2(G114), .ZN(new_n485));
  INV_X1    g060(.A(G114), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(KEYINPUT67), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n483), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n464), .A2(new_n466), .A3(G126), .A4(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n458), .ZN(new_n491));
  XOR2_X1   g066(.A(KEYINPUT69), .B(KEYINPUT4), .Z(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n457), .A2(G138), .A3(new_n458), .A4(new_n495), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n490), .A2(KEYINPUT68), .B1(new_n493), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n488), .A2(new_n498), .A3(new_n489), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n481), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n489), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n458), .B1(KEYINPUT67), .B2(new_n486), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n484), .A2(G114), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n482), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT68), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n493), .A2(new_n496), .ZN(new_n506));
  AND4_X1   g081(.A1(new_n481), .A2(new_n505), .A3(new_n499), .A4(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n500), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G651), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n512), .A2(KEYINPUT71), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(KEYINPUT71), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n513), .A2(new_n514), .B1(KEYINPUT6), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n519), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G543), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n520), .A2(new_n522), .B1(new_n519), .B2(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n516), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G88), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n510), .A2(new_n517), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n523), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n527), .A2(new_n515), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n526), .A2(new_n528), .ZN(G166));
  INV_X1    g104(.A(new_n517), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G51), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n523), .B(KEYINPUT73), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n532), .A2(G63), .A3(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT74), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  INV_X1    g112(.A(G89), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n524), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(KEYINPUT75), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n541));
  OAI211_X1 g116(.A(new_n537), .B(new_n541), .C1(new_n538), .C2(new_n524), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n534), .B1(new_n540), .B2(new_n542), .ZN(G168));
  NAND2_X1  g118(.A1(new_n530), .A2(G52), .ZN(new_n544));
  INV_X1    g119(.A(new_n524), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G90), .ZN(new_n546));
  AND3_X1   g121(.A1(new_n544), .A2(new_n546), .A3(KEYINPUT76), .ZN(new_n547));
  AOI21_X1  g122(.A(KEYINPUT76), .B1(new_n544), .B2(new_n546), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n532), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n515), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n549), .A2(new_n551), .ZN(G171));
  NAND2_X1  g127(.A1(new_n532), .A2(G56), .ZN(new_n553));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G651), .ZN(new_n556));
  INV_X1    g131(.A(G43), .ZN(new_n557));
  INV_X1    g132(.A(G81), .ZN(new_n558));
  OAI22_X1  g133(.A1(new_n557), .A2(new_n517), .B1(new_n524), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT77), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n515), .B1(new_n553), .B2(new_n554), .ZN(new_n564));
  NOR3_X1   g139(.A1(new_n564), .A2(new_n559), .A3(new_n562), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  AND3_X1   g143(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G36), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n569), .A2(new_n572), .ZN(G188));
  NAND3_X1  g148(.A1(new_n516), .A2(G53), .A3(G543), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT9), .ZN(new_n575));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n520), .A2(new_n522), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n519), .A2(G543), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(G65), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n576), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n545), .A2(G91), .B1(G651), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n575), .A2(new_n582), .ZN(G299));
  INV_X1    g158(.A(G171), .ZN(G301));
  INV_X1    g159(.A(G168), .ZN(G286));
  INV_X1    g160(.A(G166), .ZN(G303));
  AOI22_X1  g161(.A1(G49), .A2(new_n530), .B1(new_n545), .B2(G87), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n532), .A2(G74), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n515), .B2(new_n588), .ZN(G288));
  NAND2_X1  g164(.A1(new_n545), .A2(G86), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n590), .A2(KEYINPUT78), .ZN(new_n591));
  INV_X1    g166(.A(G48), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n523), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n593));
  OAI22_X1  g168(.A1(new_n517), .A2(new_n592), .B1(new_n515), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n590), .A2(KEYINPUT78), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n591), .A2(new_n595), .A3(new_n596), .ZN(G305));
  AND2_X1   g172(.A1(new_n532), .A2(G60), .ZN(new_n598));
  AND2_X1   g173(.A1(G72), .A2(G543), .ZN(new_n599));
  OAI21_X1  g174(.A(G651), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(G47), .A2(new_n530), .B1(new_n545), .B2(G85), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n600), .A2(new_n601), .ZN(new_n605));
  OR2_X1    g180(.A1(new_n604), .A2(new_n605), .ZN(G290));
  XOR2_X1   g181(.A(KEYINPUT80), .B(KEYINPUT10), .Z(new_n607));
  NAND3_X1  g182(.A1(new_n545), .A2(G92), .A3(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n607), .ZN(new_n609));
  INV_X1    g184(.A(G92), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n524), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(G54), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n523), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n614));
  OAI22_X1  g189(.A1(new_n517), .A2(new_n613), .B1(new_n515), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G171), .B2(new_n618), .ZN(G284));
  XNOR2_X1  g195(.A(G284), .B(KEYINPUT81), .ZN(G321));
  NAND2_X1  g196(.A1(G299), .A2(new_n618), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G168), .B2(new_n618), .ZN(G297));
  XNOR2_X1  g198(.A(G297), .B(KEYINPUT82), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n616), .B1(new_n625), .B2(G860), .ZN(G148));
  AOI21_X1  g201(.A(KEYINPUT77), .B1(new_n556), .B2(new_n560), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n627), .A2(new_n565), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(new_n618), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n617), .A2(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n618), .B2(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT83), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g208(.A1(new_n460), .A2(G135), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n475), .A2(G123), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n458), .A2(G111), .ZN(new_n636));
  OAI21_X1  g211(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n634), .B(new_n635), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT84), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(G2096), .Z(new_n643));
  NAND2_X1  g218(.A1(new_n457), .A2(new_n471), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT12), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT13), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2100), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n643), .A2(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT85), .B(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2427), .B(G2430), .Z(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(KEYINPUT14), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT16), .B(G1341), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G1348), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n658), .B(new_n660), .ZN(new_n661));
  OAI21_X1  g236(.A(G14), .B1(new_n655), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n662), .B1(new_n655), .B2(new_n661), .ZN(G401));
  XOR2_X1   g238(.A(G2072), .B(G2078), .Z(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT18), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n667), .B(KEYINPUT86), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(new_n666), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n666), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n664), .B(KEYINPUT17), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n670), .A2(new_n665), .A3(new_n666), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n669), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2096), .B(G2100), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT87), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n676), .B(new_n678), .ZN(G227));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  XOR2_X1   g256(.A(G1956), .B(G2474), .Z(new_n682));
  XOR2_X1   g257(.A(G1961), .B(G1966), .Z(new_n683));
  OR2_X1    g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n683), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n681), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n681), .A2(new_n686), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT20), .ZN(new_n689));
  OAI211_X1 g264(.A(new_n685), .B(new_n687), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(new_n689), .B2(new_n688), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT88), .ZN(new_n692));
  INV_X1    g267(.A(G1991), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G1996), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n695), .A2(new_n696), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  OR3_X1    g275(.A1(new_n697), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n697), .B2(new_n698), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(G229));
  MUX2_X1   g278(.A(G6), .B(G305), .S(G16), .Z(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT32), .B(G1981), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(G16), .A2(G23), .ZN(new_n707));
  INV_X1    g282(.A(G288), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(G16), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT33), .B(G1976), .Z(new_n710));
  AOI22_X1  g285(.A1(new_n704), .A2(new_n705), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G22), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G166), .B2(new_n712), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(G1971), .Z(new_n715));
  OR2_X1    g290(.A1(new_n709), .A2(new_n710), .ZN(new_n716));
  NAND4_X1  g291(.A1(new_n706), .A2(new_n711), .A3(new_n715), .A4(new_n716), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT34), .Z(new_n718));
  NAND2_X1  g293(.A1(new_n712), .A2(G24), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n604), .A2(new_n605), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(new_n712), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G1986), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n721), .A2(G1986), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n460), .A2(G131), .B1(new_n475), .B2(G119), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT89), .ZN(new_n725));
  NOR3_X1   g300(.A1(new_n725), .A2(G95), .A3(G2105), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(G95), .B2(G2105), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n727), .B(G2104), .C1(G107), .C2(new_n458), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n724), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  MUX2_X1   g304(.A(G25), .B(new_n729), .S(G29), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT90), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT35), .B(G1991), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n718), .A2(new_n722), .A3(new_n723), .A4(new_n733), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT36), .Z(new_n735));
  NOR2_X1   g310(.A1(G5), .A2(G16), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT95), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G301), .B2(new_n712), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT96), .B(G1961), .Z(new_n739));
  NOR2_X1   g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT26), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G105), .B2(new_n471), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n475), .A2(G129), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n460), .A2(G141), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G29), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G29), .B2(G32), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT27), .B(G1996), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT93), .B(KEYINPUT24), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G34), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n752), .A2(G29), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G160), .B2(G29), .ZN(new_n754));
  OAI22_X1  g329(.A1(new_n749), .A2(new_n750), .B1(G2084), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n471), .A2(G103), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(KEYINPUT25), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT25), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n471), .A2(new_n758), .A3(G103), .ZN(new_n759));
  INV_X1    g334(.A(G139), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n757), .B(new_n759), .C1(new_n459), .C2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(G115), .A2(G2104), .ZN(new_n762));
  INV_X1    g337(.A(G127), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n467), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n761), .B1(G2105), .B2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G29), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n766), .B2(G33), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n755), .B1(G2072), .B2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(G2090), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n766), .A2(G35), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G162), .B2(new_n766), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT29), .Z(new_n774));
  OAI21_X1  g349(.A(new_n770), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(G140), .ZN(new_n776));
  OR3_X1    g351(.A1(new_n459), .A2(KEYINPUT91), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(KEYINPUT91), .B1(new_n459), .B2(new_n776), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n475), .A2(G128), .ZN(new_n779));
  OR2_X1    g354(.A1(G104), .A2(G2105), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n780), .B(G2104), .C1(G116), .C2(new_n458), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n777), .A2(new_n778), .A3(new_n779), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n782), .A2(G29), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n784));
  NAND2_X1  g359(.A1(new_n766), .A2(G26), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G2067), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n774), .A2(new_n771), .ZN(new_n789));
  NOR4_X1   g364(.A1(new_n740), .A2(new_n775), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n642), .ZN(new_n791));
  AOI22_X1  g366(.A1(new_n791), .A2(G29), .B1(G2084), .B2(new_n754), .ZN(new_n792));
  INV_X1    g367(.A(G28), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n793), .A2(KEYINPUT30), .ZN(new_n794));
  AOI21_X1  g369(.A(G29), .B1(new_n793), .B2(KEYINPUT30), .ZN(new_n795));
  OR2_X1    g370(.A1(KEYINPUT31), .A2(G11), .ZN(new_n796));
  NAND2_X1  g371(.A1(KEYINPUT31), .A2(G11), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n794), .A2(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n792), .B(new_n798), .C1(new_n769), .C2(G2072), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n749), .A2(new_n750), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT94), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n712), .A2(G4), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n616), .B2(new_n712), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n803), .A2(G1348), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n803), .A2(G1348), .ZN(new_n805));
  NOR4_X1   g380(.A1(new_n799), .A2(new_n801), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT23), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n712), .A2(G20), .ZN(new_n808));
  AOI211_X1 g383(.A(new_n807), .B(new_n808), .C1(G299), .C2(G16), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n807), .B2(new_n808), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT98), .B(G1956), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(G27), .A2(G29), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G164), .B2(G29), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT97), .B(G2078), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n790), .A2(new_n806), .A3(new_n812), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(G168), .A2(G16), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G16), .B2(G21), .ZN(new_n819));
  INV_X1    g394(.A(G1966), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n738), .B2(new_n739), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n712), .A2(G19), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(new_n567), .B2(new_n712), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n824), .A2(G1341), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(G1341), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n819), .A2(new_n820), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n822), .A2(new_n825), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  NOR3_X1   g403(.A1(new_n735), .A2(new_n817), .A3(new_n828), .ZN(G311));
  INV_X1    g404(.A(G311), .ZN(G150));
  AOI22_X1  g405(.A1(new_n532), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n831), .A2(new_n515), .ZN(new_n832));
  INV_X1    g407(.A(G55), .ZN(new_n833));
  INV_X1    g408(.A(G93), .ZN(new_n834));
  OAI22_X1  g409(.A1(new_n833), .A2(new_n517), .B1(new_n524), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(G860), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT37), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n628), .A2(new_n836), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n836), .A2(new_n561), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT39), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n616), .A2(G559), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT38), .Z(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(new_n837), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n844), .A2(new_n846), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n839), .B1(new_n848), .B2(new_n849), .ZN(G145));
  NAND2_X1  g425(.A1(new_n460), .A2(G142), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n475), .A2(G130), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n458), .A2(G118), .ZN(new_n853));
  OAI21_X1  g428(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n851), .B(new_n852), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n765), .B(new_n855), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n782), .B(new_n645), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n490), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(new_n506), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n858), .B(new_n860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(new_n729), .Z(new_n862));
  XNOR2_X1  g437(.A(new_n642), .B(G160), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n746), .B(new_n479), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(G37), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n866), .B1(new_n865), .B2(new_n862), .ZN(new_n867));
  XNOR2_X1  g442(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(G395));
  NAND2_X1  g444(.A1(G290), .A2(new_n708), .ZN(new_n870));
  OR2_X1    g445(.A1(G305), .A2(G166), .ZN(new_n871));
  NAND2_X1  g446(.A1(G305), .A2(G166), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n720), .A2(G288), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n870), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n873), .B1(new_n870), .B2(new_n874), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT42), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n843), .B(new_n630), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n616), .B(G299), .Z(new_n880));
  OR2_X1    g455(.A1(new_n880), .A2(KEYINPUT41), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(KEYINPUT41), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n884), .B1(new_n880), .B2(new_n879), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n878), .A2(new_n885), .ZN(new_n886));
  AND2_X1   g461(.A1(new_n886), .A2(KEYINPUT100), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n878), .A2(new_n885), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(new_n886), .B2(KEYINPUT100), .ZN(new_n889));
  OAI21_X1  g464(.A(G868), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(KEYINPUT101), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT101), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n892), .B(G868), .C1(new_n887), .C2(new_n889), .ZN(new_n893));
  INV_X1    g468(.A(new_n836), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(new_n618), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n891), .A2(new_n893), .A3(new_n895), .ZN(G295));
  NAND3_X1  g471(.A1(new_n891), .A2(new_n893), .A3(new_n895), .ZN(G331));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n898));
  OR2_X1    g473(.A1(new_n547), .A2(new_n548), .ZN(new_n899));
  INV_X1    g474(.A(new_n551), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n899), .A2(G286), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(G168), .B1(new_n549), .B2(new_n551), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n903), .B1(new_n840), .B2(new_n842), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n567), .A2(new_n894), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n905), .A2(new_n841), .A3(new_n902), .A4(new_n901), .ZN(new_n906));
  AOI22_X1  g481(.A1(new_n881), .A2(new_n882), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n904), .A2(new_n906), .A3(KEYINPUT102), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT102), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n903), .B(new_n910), .C1(new_n840), .C2(new_n842), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n898), .B(new_n908), .C1(new_n912), .C2(new_n880), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n870), .A2(new_n874), .ZN(new_n914));
  INV_X1    g489(.A(new_n873), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n870), .A2(new_n873), .A3(new_n874), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n916), .A2(KEYINPUT104), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(KEYINPUT104), .B1(new_n916), .B2(new_n917), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n880), .B1(new_n909), .B2(new_n911), .ZN(new_n921));
  OAI21_X1  g496(.A(KEYINPUT103), .B1(new_n921), .B2(new_n907), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n913), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  NOR3_X1   g498(.A1(new_n921), .A2(new_n877), .A3(new_n907), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n924), .A2(G37), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n909), .A2(new_n883), .A3(new_n911), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n904), .A2(new_n906), .ZN(new_n930));
  OAI22_X1  g505(.A1(new_n929), .A2(KEYINPUT105), .B1(new_n880), .B2(new_n930), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n929), .A2(KEYINPUT105), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n920), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n933), .A2(new_n925), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n928), .B(KEYINPUT44), .C1(new_n927), .C2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n933), .A2(new_n925), .A3(new_n927), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n937), .B1(new_n926), .B2(new_n927), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n933), .A2(new_n927), .A3(new_n925), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n927), .B1(new_n923), .B2(new_n925), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n936), .B(new_n939), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n935), .B1(new_n940), .B2(new_n944), .ZN(G397));
  XOR2_X1   g520(.A(new_n782), .B(G2067), .Z(new_n946));
  INV_X1    g521(.A(G1996), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n746), .B(new_n947), .ZN(new_n948));
  OR2_X1    g523(.A1(new_n729), .A2(new_n732), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n729), .A2(new_n732), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n946), .A2(new_n948), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  XOR2_X1   g526(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(G1384), .B1(new_n859), .B2(new_n506), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n953), .B1(new_n954), .B2(KEYINPUT107), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n955), .B1(KEYINPUT107), .B2(new_n954), .ZN(new_n956));
  AND4_X1   g531(.A1(G40), .A2(new_n461), .A3(new_n470), .A4(new_n472), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n951), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(G290), .B(G1986), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n960), .B1(new_n961), .B2(new_n959), .ZN(new_n962));
  XOR2_X1   g537(.A(new_n962), .B(KEYINPUT109), .Z(new_n963));
  OAI21_X1  g538(.A(new_n957), .B1(KEYINPUT45), .B2(new_n954), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n505), .A2(new_n499), .A3(new_n506), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT70), .ZN(new_n966));
  INV_X1    g541(.A(G1384), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n505), .A2(new_n499), .A3(new_n506), .A4(new_n481), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n966), .A2(new_n967), .A3(new_n968), .A4(new_n952), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n964), .B1(new_n969), .B2(KEYINPUT114), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT114), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n508), .A2(new_n971), .A3(new_n967), .A4(new_n952), .ZN(new_n972));
  AOI21_X1  g547(.A(G1966), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n974), .A2(KEYINPUT111), .A3(KEYINPUT50), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT111), .B1(new_n974), .B2(KEYINPUT50), .ZN(new_n976));
  INV_X1    g551(.A(new_n954), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n957), .B1(new_n977), .B2(KEYINPUT50), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n975), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G2084), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n973), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(G286), .A2(KEYINPUT118), .A3(G8), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT118), .ZN(new_n983));
  INV_X1    g558(.A(G8), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n983), .B1(G168), .B2(new_n984), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  OR2_X1    g561(.A1(new_n981), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n986), .B1(new_n981), .B2(new_n984), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT119), .B1(new_n988), .B2(KEYINPUT51), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n969), .A2(KEYINPUT114), .ZN(new_n990));
  INV_X1    g565(.A(new_n964), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n969), .A2(KEYINPUT114), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n820), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n974), .A2(KEYINPUT50), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT111), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n974), .A2(KEYINPUT111), .A3(KEYINPUT50), .ZN(new_n998));
  INV_X1    g573(.A(new_n978), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n997), .A2(new_n980), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n984), .B1(new_n994), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n982), .A2(new_n985), .ZN(new_n1002));
  OAI211_X1 g577(.A(KEYINPUT119), .B(KEYINPUT51), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n1004), .B(new_n986), .C1(new_n981), .C2(new_n984), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n987), .B1(new_n989), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT120), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT62), .ZN(new_n1010));
  OAI211_X1 g585(.A(KEYINPUT120), .B(new_n987), .C1(new_n989), .C2(new_n1006), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT123), .ZN(new_n1013));
  INV_X1    g588(.A(new_n957), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1014), .A2(new_n977), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1015), .A2(new_n984), .ZN(new_n1016));
  INV_X1    g591(.A(G1976), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1016), .A2(new_n1017), .A3(G288), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1016), .B(new_n1021), .C1(G288), .C2(new_n1017), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1020), .B(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n595), .A2(new_n590), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(G1981), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1025), .B1(G305), .B2(G1981), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT49), .ZN(new_n1027));
  OR2_X1    g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AOI211_X1 g603(.A(new_n984), .B(new_n1015), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1023), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n978), .B1(new_n995), .B2(new_n996), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n998), .ZN(new_n1032));
  OR3_X1    g607(.A1(new_n1032), .A2(KEYINPUT112), .A3(G2090), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n954), .A2(KEYINPUT45), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n957), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1035), .B1(new_n974), .B2(new_n953), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1036), .A2(G1971), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT110), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n1037), .B(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT112), .B1(new_n1032), .B2(G2090), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1033), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(G303), .A2(G8), .ZN(new_n1042));
  XOR2_X1   g617(.A(new_n1042), .B(KEYINPUT55), .Z(new_n1043));
  NAND3_X1  g618(.A1(new_n1041), .A2(G8), .A3(new_n1043), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1030), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1043), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT50), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n508), .A2(new_n1047), .A3(new_n967), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1014), .B1(KEYINPUT50), .B2(new_n977), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1050), .A2(G2090), .ZN(new_n1051));
  OAI21_X1  g626(.A(G8), .B1(new_n1051), .B2(new_n1037), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1046), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(G1961), .B1(new_n1031), .B2(new_n998), .ZN(new_n1054));
  INV_X1    g629(.A(G2078), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT53), .B1(new_n1036), .B2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n970), .A2(new_n972), .A3(KEYINPUT53), .A4(new_n1055), .ZN(new_n1058));
  AOI21_X1  g633(.A(G301), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1045), .A2(new_n1053), .A3(new_n1059), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1012), .A2(new_n1013), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1013), .B1(new_n1012), .B2(new_n1060), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1010), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1063));
  NOR3_X1   g638(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1030), .A2(G8), .A3(new_n1043), .A4(new_n1041), .ZN(new_n1065));
  AOI211_X1 g640(.A(G1976), .B(G288), .C1(new_n1029), .C2(new_n1028), .ZN(new_n1066));
  NOR2_X1   g641(.A1(G305), .A2(G1981), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1016), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1065), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT63), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1041), .A2(G8), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1070), .B1(new_n1071), .B2(new_n1046), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1045), .A2(G168), .A3(new_n1072), .A4(new_n1001), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1069), .B1(new_n1073), .B2(KEYINPUT63), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1001), .A2(G168), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1075), .B1(new_n1045), .B2(new_n1072), .ZN(new_n1076));
  INV_X1    g651(.A(G1956), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1050), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n1079));
  NAND2_X1  g654(.A1(G299), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n575), .A2(new_n582), .A3(KEYINPUT57), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  XOR2_X1   g657(.A(KEYINPUT56), .B(G2072), .Z(new_n1083));
  XNOR2_X1  g658(.A(new_n1083), .B(KEYINPUT115), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1036), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1078), .A2(new_n1082), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT116), .ZN(new_n1087));
  NOR3_X1   g662(.A1(new_n1014), .A2(new_n977), .A3(G2067), .ZN(new_n1088));
  INV_X1    g663(.A(G1348), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1088), .B1(new_n1032), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1087), .B1(new_n1090), .B2(new_n617), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1036), .A2(new_n1084), .ZN(new_n1092));
  AOI21_X1  g667(.A(G1956), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1080), .B(new_n1081), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1091), .A2(new_n1094), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n1090), .A2(new_n1087), .A3(new_n617), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1086), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n617), .A2(KEYINPUT60), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1090), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n1100));
  XNOR2_X1  g675(.A(KEYINPUT58), .B(G1341), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1015), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1102), .B1(new_n1036), .B2(new_n947), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1100), .B1(new_n1103), .B2(new_n628), .ZN(new_n1104));
  OR3_X1    g679(.A1(new_n1103), .A2(new_n628), .A3(new_n1100), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1099), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1090), .A2(new_n617), .ZN(new_n1107));
  AOI211_X1 g682(.A(new_n616), .B(new_n1088), .C1(new_n1032), .C2(new_n1089), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT60), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1094), .A2(new_n1086), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT61), .B1(new_n1111), .B2(KEYINPUT117), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT117), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n1114));
  AOI211_X1 g689(.A(new_n1113), .B(new_n1114), .C1(new_n1094), .C2(new_n1086), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1097), .B1(new_n1110), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT54), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1055), .A2(KEYINPUT53), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1119), .B1(new_n1014), .B2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1121), .B(new_n1034), .C1(new_n1120), .C2(new_n1014), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1122), .A2(new_n956), .ZN(new_n1123));
  NOR4_X1   g698(.A1(new_n1054), .A2(new_n1123), .A3(new_n1056), .A4(G171), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1118), .B1(new_n1059), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(KEYINPUT122), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1127), .B(new_n1118), .C1(new_n1059), .C2(new_n1124), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1057), .A2(G301), .A3(new_n1058), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1054), .A2(new_n1123), .A3(new_n1056), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1130), .B(KEYINPUT54), .C1(G301), .C2(new_n1131), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1117), .A2(new_n1129), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1076), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1045), .A2(new_n1053), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1074), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n963), .B1(new_n1064), .B2(new_n1137), .ZN(new_n1138));
  OR2_X1    g713(.A1(G290), .A2(G1986), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT48), .ZN(new_n1140));
  OR3_X1    g715(.A1(new_n1139), .A2(new_n1140), .A3(new_n958), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1140), .B1(new_n1139), .B2(new_n958), .ZN(new_n1142));
  XOR2_X1   g717(.A(new_n960), .B(KEYINPUT125), .Z(new_n1143));
  AND3_X1   g718(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n959), .A2(KEYINPUT46), .A3(new_n947), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT46), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(new_n958), .B2(G1996), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n946), .A2(new_n747), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1145), .B(new_n1147), .C1(new_n958), .C2(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n1149), .B(KEYINPUT124), .ZN(new_n1150));
  XOR2_X1   g725(.A(new_n1150), .B(KEYINPUT47), .Z(new_n1151));
  NAND2_X1  g726(.A1(new_n946), .A2(new_n948), .ZN(new_n1152));
  OAI22_X1  g727(.A1(new_n1152), .A2(new_n949), .B1(G2067), .B2(new_n782), .ZN(new_n1153));
  AOI211_X1 g728(.A(new_n1144), .B(new_n1151), .C1(new_n959), .C2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1138), .A2(new_n1154), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g730(.A(G319), .ZN(new_n1157));
  NOR2_X1   g731(.A1(G227), .A2(new_n1157), .ZN(new_n1158));
  XOR2_X1   g732(.A(new_n1158), .B(KEYINPUT126), .Z(new_n1159));
  NOR2_X1   g733(.A1(new_n1159), .A2(G401), .ZN(new_n1160));
  AND4_X1   g734(.A1(new_n701), .A2(new_n867), .A3(new_n702), .A4(new_n1160), .ZN(new_n1161));
  NAND2_X1  g735(.A1(new_n1161), .A2(new_n938), .ZN(G225));
  NAND2_X1  g736(.A1(G225), .A2(KEYINPUT127), .ZN(new_n1163));
  INV_X1    g737(.A(KEYINPUT127), .ZN(new_n1164));
  NAND3_X1  g738(.A1(new_n1161), .A2(new_n938), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1165), .ZN(G308));
endmodule


