//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 0 0 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 0 1 0 0 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n562, new_n564, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n630,
    new_n633, new_n635, new_n636, new_n637, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1234, new_n1235, new_n1236, new_n1237;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n461), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND3_X1   g044(.A1(new_n461), .A2(KEYINPUT68), .A3(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(KEYINPUT68), .B1(new_n461), .B2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G101), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n463), .A2(new_n465), .ZN(new_n475));
  INV_X1    g050(.A(G137), .ZN(new_n476));
  NOR3_X1   g051(.A1(new_n475), .A2(new_n476), .A3(G2105), .ZN(new_n477));
  OR3_X1    g052(.A1(new_n474), .A2(KEYINPUT69), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g053(.A(KEYINPUT69), .B1(new_n474), .B2(new_n477), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n469), .B1(new_n478), .B2(new_n479), .ZN(G160));
  INV_X1    g055(.A(KEYINPUT70), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n475), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n463), .A2(new_n465), .A3(KEYINPUT70), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n482), .A2(G2105), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n461), .A3(new_n483), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n486), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT4), .B1(new_n494), .B2(new_n462), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(new_n466), .B2(G126), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(KEYINPUT71), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(new_n463), .A3(new_n465), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  AOI21_X1  g075(.A(G2105), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n466), .A2(KEYINPUT4), .A3(new_n498), .ZN(new_n503));
  NAND2_X1  g078(.A1(G102), .A2(G2104), .ZN(new_n504));
  AOI21_X1  g079(.A(G2105), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n502), .A2(new_n505), .ZN(G164));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G651), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n508), .A2(new_n510), .A3(new_n516), .A4(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n516), .A2(new_n518), .A3(G543), .ZN(new_n521));
  INV_X1    g096(.A(G50), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n515), .A2(new_n523), .ZN(G166));
  AND4_X1   g099(.A1(new_n508), .A2(new_n510), .A3(new_n516), .A4(new_n518), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT7), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n528), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n525), .A2(G89), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT73), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n521), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n516), .A2(new_n518), .A3(KEYINPUT73), .A4(G543), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n532), .A2(G51), .A3(new_n533), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n508), .A2(new_n510), .A3(KEYINPUT72), .ZN(new_n535));
  AOI21_X1  g110(.A(KEYINPUT72), .B1(new_n508), .B2(new_n510), .ZN(new_n536));
  OAI211_X1 g111(.A(G63), .B(G651), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  AND3_X1   g112(.A1(new_n530), .A2(new_n534), .A3(new_n537), .ZN(G168));
  OAI21_X1  g113(.A(G64), .B1(new_n535), .B2(new_n536), .ZN(new_n539));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n514), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT74), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n532), .A2(new_n533), .ZN(new_n543));
  XNOR2_X1  g118(.A(KEYINPUT75), .B(G90), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n543), .A2(G52), .B1(new_n525), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n542), .A2(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  NAND3_X1  g122(.A1(new_n532), .A2(G43), .A3(new_n533), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n525), .A2(G81), .ZN(new_n549));
  AND2_X1   g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT72), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n511), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n508), .A2(new_n510), .A3(KEYINPUT72), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n551), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  OAI21_X1  g132(.A(G651), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n550), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  AND3_X1   g136(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G36), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(G188));
  NAND4_X1  g141(.A1(new_n516), .A2(new_n518), .A3(G53), .A4(G543), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT9), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  XOR2_X1   g144(.A(KEYINPUT77), .B(G65), .Z(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n570), .B2(new_n511), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G651), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n573));
  AND3_X1   g148(.A1(new_n525), .A2(new_n573), .A3(G91), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n573), .B1(new_n525), .B2(G91), .ZN(new_n575));
  OAI211_X1 g150(.A(new_n568), .B(new_n572), .C1(new_n574), .C2(new_n575), .ZN(G299));
  INV_X1    g151(.A(G168), .ZN(G286));
  XNOR2_X1  g152(.A(G166), .B(KEYINPUT78), .ZN(G303));
  INV_X1    g153(.A(G74), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n553), .A2(new_n579), .A3(new_n554), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G651), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n521), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n525), .A2(G87), .B1(new_n584), .B2(G49), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n580), .A2(KEYINPUT79), .A3(G651), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n583), .A2(new_n585), .A3(new_n586), .ZN(G288));
  AND3_X1   g162(.A1(new_n508), .A2(new_n510), .A3(G61), .ZN(new_n588));
  INV_X1    g163(.A(G73), .ZN(new_n589));
  OAI21_X1  g164(.A(KEYINPUT80), .B1(new_n589), .B2(new_n507), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT80), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n591), .A2(G73), .A3(G543), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n588), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(KEYINPUT81), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n525), .A2(G86), .B1(new_n584), .B2(G48), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT81), .ZN(new_n597));
  OAI211_X1 g172(.A(new_n597), .B(G651), .C1(new_n588), .C2(new_n593), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT82), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n595), .A2(new_n596), .A3(KEYINPUT82), .A4(new_n598), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(G305));
  OAI21_X1  g178(.A(G60), .B1(new_n535), .B2(new_n536), .ZN(new_n604));
  AND2_X1   g179(.A1(G72), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G651), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT83), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n543), .A2(G47), .B1(G85), .B2(new_n525), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n607), .A2(KEYINPUT83), .A3(G651), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(G290));
  NAND2_X1  g188(.A1(G301), .A2(G868), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT84), .Z(new_n615));
  INV_X1    g190(.A(G92), .ZN(new_n616));
  XNOR2_X1  g191(.A(KEYINPUT85), .B(KEYINPUT10), .ZN(new_n617));
  OR3_X1    g192(.A1(new_n519), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n532), .A2(G54), .A3(new_n533), .ZN(new_n619));
  NAND2_X1  g194(.A1(G79), .A2(G543), .ZN(new_n620));
  INV_X1    g195(.A(G66), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n511), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G651), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n617), .B1(new_n519), .B2(new_n616), .ZN(new_n624));
  NAND4_X1  g199(.A1(new_n618), .A2(new_n619), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n615), .B1(G868), .B2(new_n626), .ZN(G284));
  OAI21_X1  g202(.A(new_n615), .B1(G868), .B2(new_n626), .ZN(G321));
  INV_X1    g203(.A(G868), .ZN(new_n629));
  NAND2_X1  g204(.A1(G299), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(new_n629), .B2(G168), .ZN(G297));
  OAI21_X1  g206(.A(new_n630), .B1(new_n629), .B2(G168), .ZN(G280));
  INV_X1    g207(.A(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n626), .B1(new_n633), .B2(G860), .ZN(G148));
  NAND2_X1  g209(.A1(new_n559), .A2(new_n629), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n625), .A2(G559), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT86), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n635), .B1(new_n637), .B2(new_n629), .ZN(G323));
  XNOR2_X1  g213(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g214(.A(new_n466), .B1(new_n471), .B2(new_n470), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT12), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT13), .Z(new_n642));
  OR2_X1    g217(.A1(new_n642), .A2(G2100), .ZN(new_n643));
  OR2_X1    g218(.A1(G99), .A2(G2105), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n644), .B(G2104), .C1(G111), .C2(new_n461), .ZN(new_n645));
  INV_X1    g220(.A(G123), .ZN(new_n646));
  INV_X1    g221(.A(G135), .ZN(new_n647));
  OAI221_X1 g222(.A(new_n645), .B1(new_n484), .B2(new_n646), .C1(new_n647), .C2(new_n487), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(G2096), .Z(new_n649));
  NAND2_X1  g224(.A1(new_n642), .A2(G2100), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n643), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT87), .ZN(G156));
  XOR2_X1   g227(.A(KEYINPUT88), .B(G2438), .Z(new_n653));
  XNOR2_X1  g228(.A(G2427), .B(G2430), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(KEYINPUT15), .B(G2435), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(KEYINPUT14), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  INV_X1    g237(.A(new_n660), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n657), .A2(KEYINPUT14), .A3(new_n663), .ZN(new_n664));
  AND3_X1   g239(.A1(new_n661), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n662), .B1(new_n661), .B2(new_n664), .ZN(new_n666));
  XOR2_X1   g241(.A(G1341), .B(G1348), .Z(new_n667));
  OR3_X1    g242(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT89), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(G14), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n665), .A2(new_n666), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n671), .B1(new_n673), .B2(new_n667), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(G401));
  XOR2_X1   g251(.A(G2084), .B(G2090), .Z(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G2067), .B(G2678), .Z(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G2072), .B(G2078), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n678), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT90), .Z(new_n683));
  XOR2_X1   g258(.A(new_n681), .B(KEYINPUT17), .Z(new_n684));
  OAI21_X1  g259(.A(new_n683), .B1(new_n679), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n680), .A2(new_n681), .A3(new_n677), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT18), .Z(new_n687));
  NAND3_X1  g262(.A1(new_n684), .A2(new_n679), .A3(new_n677), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n685), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G2096), .B(G2100), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(G227));
  XOR2_X1   g267(.A(G1956), .B(G2474), .Z(new_n693));
  XOR2_X1   g268(.A(G1961), .B(G1966), .Z(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1971), .B(G1976), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT19), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n693), .A2(new_n694), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT20), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n699), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n696), .A2(new_n698), .A3(new_n700), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n703), .B(new_n704), .C1(new_n702), .C2(new_n701), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(G1991), .B(G1996), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G1981), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G1986), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n707), .B(new_n710), .ZN(G229));
  INV_X1    g286(.A(KEYINPUT95), .ZN(new_n712));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G23), .ZN(new_n714));
  INV_X1    g289(.A(G288), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n713), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT94), .B(KEYINPUT33), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G1976), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n716), .B(new_n718), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n713), .A2(G6), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G305), .B2(G16), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT32), .B(G1981), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT93), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n515), .A2(new_n523), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G16), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n713), .A2(G22), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(G1971), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n721), .A2(new_n723), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n719), .A2(new_n724), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n712), .B1(new_n732), .B2(KEYINPUT34), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n732), .A2(new_n712), .A3(KEYINPUT34), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT34), .ZN(new_n736));
  INV_X1    g311(.A(new_n732), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n734), .A2(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT36), .ZN(new_n739));
  INV_X1    g314(.A(G29), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G25), .ZN(new_n741));
  AND3_X1   g316(.A1(new_n463), .A2(new_n465), .A3(KEYINPUT70), .ZN(new_n742));
  AOI21_X1  g317(.A(KEYINPUT70), .B1(new_n463), .B2(new_n465), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g319(.A1(new_n744), .A2(KEYINPUT91), .A3(G119), .A4(G2105), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n482), .A2(G119), .A3(G2105), .A4(new_n483), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT91), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n749));
  INV_X1    g324(.A(G107), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n749), .B1(new_n750), .B2(G2105), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT92), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n744), .A2(G131), .A3(new_n461), .ZN(new_n754));
  NAND4_X1  g329(.A1(new_n745), .A2(new_n748), .A3(new_n753), .A4(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n741), .B1(new_n756), .B2(new_n740), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT35), .B(G1991), .Z(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  OR2_X1    g334(.A1(G16), .A2(G24), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G290), .B2(new_n713), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(G1986), .Z(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n738), .A2(new_n739), .A3(new_n759), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n737), .A2(new_n736), .ZN(new_n765));
  INV_X1    g340(.A(new_n735), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n759), .B(new_n765), .C1(new_n766), .C2(new_n733), .ZN(new_n767));
  OAI21_X1  g342(.A(KEYINPUT36), .B1(new_n767), .B2(new_n762), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n713), .A2(G4), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n626), .B2(new_n713), .ZN(new_n771));
  INV_X1    g346(.A(G1348), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n713), .A2(G19), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n560), .B2(new_n713), .ZN(new_n775));
  MUX2_X1   g350(.A(new_n774), .B(new_n775), .S(KEYINPUT96), .Z(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(G1341), .Z(new_n777));
  NAND2_X1  g352(.A1(G164), .A2(G29), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G27), .B2(G29), .ZN(new_n779));
  INV_X1    g354(.A(G2078), .ZN(new_n780));
  INV_X1    g355(.A(G2072), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT97), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G29), .B2(G33), .ZN(new_n783));
  OR3_X1    g358(.A1(new_n782), .A2(G29), .A3(G33), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n785), .A2(KEYINPUT98), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(KEYINPUT98), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT25), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(G115), .A2(G2104), .ZN(new_n791));
  INV_X1    g366(.A(G127), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n475), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n793), .A2(G2105), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n482), .A2(G139), .A3(new_n461), .A4(new_n483), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n786), .A2(KEYINPUT25), .A3(new_n787), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n790), .A2(new_n794), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n783), .B(new_n784), .C1(new_n797), .C2(new_n740), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n779), .A2(new_n780), .B1(new_n781), .B2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT30), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n740), .B1(new_n800), .B2(G28), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(KEYINPUT102), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n800), .A2(G28), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n801), .A2(KEYINPUT102), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  AND3_X1   g380(.A1(new_n777), .A2(new_n799), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(G168), .A2(G16), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G16), .B2(G21), .ZN(new_n808));
  INV_X1    g383(.A(G1966), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n779), .A2(new_n780), .ZN(new_n811));
  INV_X1    g386(.A(G11), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n812), .A2(KEYINPUT31), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n798), .A2(new_n781), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n812), .A2(KEYINPUT31), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n648), .B2(new_n740), .ZN(new_n816));
  NOR4_X1   g391(.A1(new_n811), .A2(new_n813), .A3(new_n814), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n713), .A2(G5), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G171), .B2(new_n713), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(G1961), .Z(new_n820));
  NAND4_X1  g395(.A1(new_n806), .A2(new_n810), .A3(new_n817), .A4(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT103), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n740), .A2(G35), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n492), .A2(G29), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n822), .B2(new_n823), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT29), .Z(new_n826));
  INV_X1    g401(.A(G2090), .ZN(new_n827));
  INV_X1    g402(.A(G2084), .ZN(new_n828));
  AND2_X1   g403(.A1(KEYINPUT24), .A2(G34), .ZN(new_n829));
  NOR2_X1   g404(.A1(KEYINPUT24), .A2(G34), .ZN(new_n830));
  NOR3_X1   g405(.A1(new_n829), .A2(new_n830), .A3(G29), .ZN(new_n831));
  INV_X1    g406(.A(G160), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n831), .B1(new_n832), .B2(G29), .ZN(new_n833));
  OAI22_X1  g408(.A1(new_n826), .A2(new_n827), .B1(new_n828), .B2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(G105), .ZN(new_n835));
  OAI21_X1  g410(.A(KEYINPUT99), .B1(new_n472), .B2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT99), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n837), .B(G105), .C1(new_n470), .C2(new_n471), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n744), .A2(G129), .A3(G2105), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n744), .A2(G141), .A3(new_n461), .ZN(new_n841));
  NAND3_X1  g416(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT26), .Z(new_n843));
  NAND4_X1  g418(.A1(new_n839), .A2(new_n840), .A3(new_n841), .A4(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(G29), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(G29), .B2(G32), .ZN(new_n847));
  XOR2_X1   g422(.A(KEYINPUT27), .B(G1996), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT100), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT101), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n834), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n833), .A2(new_n828), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n740), .A2(G26), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n485), .A2(G128), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n488), .A2(G140), .ZN(new_n856));
  OR2_X1    g431(.A1(G104), .A2(G2105), .ZN(new_n857));
  OAI211_X1 g432(.A(new_n857), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n855), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n854), .B1(new_n859), .B2(G29), .ZN(new_n860));
  MUX2_X1   g435(.A(new_n854), .B(new_n860), .S(KEYINPUT28), .Z(new_n861));
  INV_X1    g436(.A(G2067), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(G299), .A2(G16), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n713), .A2(KEYINPUT23), .A3(G20), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT23), .ZN(new_n866));
  INV_X1    g441(.A(G20), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n866), .B1(new_n867), .B2(G16), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n864), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(G1956), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n863), .A2(new_n870), .ZN(new_n871));
  OAI22_X1  g446(.A1(new_n847), .A2(new_n849), .B1(new_n809), .B2(new_n808), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n872), .B1(new_n826), .B2(new_n827), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n852), .A2(new_n853), .A3(new_n871), .A4(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n821), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n769), .A2(new_n773), .A3(new_n875), .ZN(G150));
  NAND2_X1  g451(.A1(G150), .A2(KEYINPUT104), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT104), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n769), .A2(new_n878), .A3(new_n773), .A4(new_n875), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(G311));
  NAND3_X1  g455(.A1(new_n532), .A2(G55), .A3(new_n533), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n525), .A2(G93), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(G67), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(new_n553), .B2(new_n554), .ZN(new_n885));
  NAND2_X1  g460(.A1(G80), .A2(G543), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(G651), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(G860), .ZN(new_n890));
  XOR2_X1   g465(.A(new_n890), .B(KEYINPUT37), .Z(new_n891));
  OAI21_X1  g466(.A(G67), .B1(new_n535), .B2(new_n536), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n514), .B1(new_n892), .B2(new_n886), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n881), .A2(new_n882), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n550), .B(new_n558), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(G56), .B1(new_n535), .B2(new_n536), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n514), .B1(new_n896), .B2(new_n556), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n548), .A2(new_n549), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n883), .B(new_n888), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT39), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n626), .A2(G559), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT38), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n901), .B(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n891), .B1(new_n904), .B2(G860), .ZN(G145));
  XNOR2_X1  g480(.A(G160), .B(new_n492), .ZN(new_n906));
  XOR2_X1   g481(.A(new_n906), .B(new_n648), .Z(new_n907));
  NAND2_X1  g482(.A1(new_n859), .A2(G164), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n839), .A2(new_n841), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n909), .A2(new_n797), .A3(new_n840), .A4(new_n843), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n504), .B1(new_n499), .B2(new_n500), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(new_n461), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n912), .B1(new_n501), .B2(new_n496), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n913), .A2(new_n855), .A3(new_n856), .A4(new_n858), .ZN(new_n914));
  INV_X1    g489(.A(new_n797), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n844), .ZN(new_n916));
  AND4_X1   g491(.A1(new_n908), .A2(new_n910), .A3(new_n914), .A4(new_n916), .ZN(new_n917));
  AOI22_X1  g492(.A1(new_n916), .A2(new_n910), .B1(new_n908), .B2(new_n914), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n744), .A2(new_n920), .A3(G142), .A4(new_n461), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n482), .A2(G142), .A3(new_n461), .A4(new_n483), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(KEYINPUT105), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n744), .A2(G130), .A3(G2105), .ZN(new_n924));
  OR2_X1    g499(.A1(G106), .A2(G2105), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n925), .B(G2104), .C1(G118), .C2(new_n461), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n921), .A2(new_n923), .A3(new_n924), .A4(new_n926), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n754), .A2(new_n753), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n927), .A2(new_n928), .A3(new_n748), .A4(new_n745), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n924), .A2(new_n926), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n755), .A2(new_n930), .A3(new_n923), .A4(new_n921), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n929), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n932), .B1(new_n929), .B2(new_n931), .ZN(new_n934));
  NOR3_X1   g509(.A1(new_n933), .A2(new_n934), .A3(new_n641), .ZN(new_n935));
  INV_X1    g510(.A(new_n641), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n929), .A2(new_n931), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT106), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n929), .A2(new_n931), .A3(new_n932), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI211_X1 g515(.A(KEYINPUT107), .B(new_n919), .C1(new_n935), .C2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n641), .B1(new_n933), .B2(new_n934), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n938), .A2(new_n936), .A3(new_n939), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n917), .A2(new_n918), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n942), .A2(new_n943), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT107), .B1(new_n947), .B2(new_n919), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n907), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT108), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n945), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n947), .A2(new_n919), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n907), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n947), .A2(new_n950), .A3(new_n919), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(G37), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n949), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g534(.A1(new_n889), .A2(new_n629), .ZN(new_n960));
  XOR2_X1   g535(.A(new_n637), .B(new_n900), .Z(new_n961));
  AND2_X1   g536(.A1(new_n626), .A2(G299), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n626), .A2(G299), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT41), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT41), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n966), .B1(new_n962), .B2(new_n963), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n961), .A2(new_n968), .ZN(new_n969));
  XOR2_X1   g544(.A(new_n969), .B(KEYINPUT109), .Z(new_n970));
  OAI21_X1  g545(.A(new_n970), .B1(new_n964), .B2(new_n961), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT110), .ZN(new_n972));
  NAND2_X1  g547(.A1(G305), .A2(G166), .ZN(new_n973));
  NAND2_X1  g548(.A1(G290), .A2(new_n715), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n601), .A2(new_n725), .A3(new_n602), .ZN(new_n975));
  NAND4_X1  g550(.A1(G288), .A2(new_n610), .A3(new_n611), .A4(new_n612), .ZN(new_n976));
  AND4_X1   g551(.A1(new_n973), .A2(new_n974), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  AOI22_X1  g552(.A1(new_n973), .A2(new_n975), .B1(new_n974), .B2(new_n976), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n972), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n973), .A2(new_n975), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n974), .A2(new_n976), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n973), .A2(new_n974), .A3(new_n975), .A4(new_n976), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n982), .A2(KEYINPUT110), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n979), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT42), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n982), .A2(new_n983), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n986), .B1(KEYINPUT42), .B2(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n971), .B(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n960), .B1(new_n989), .B2(new_n629), .ZN(G295));
  OAI21_X1  g565(.A(new_n960), .B1(new_n989), .B2(new_n629), .ZN(G331));
  INV_X1    g566(.A(KEYINPUT111), .ZN(new_n992));
  NOR2_X1   g567(.A1(G168), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n993), .B1(new_n542), .B2(new_n545), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n527), .A2(new_n529), .ZN(new_n996));
  INV_X1    g571(.A(G89), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n996), .B1(new_n519), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G63), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n999), .B1(new_n553), .B2(new_n554), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n998), .B1(new_n1000), .B2(G651), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT112), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n1001), .A2(new_n992), .A3(new_n1002), .A4(new_n534), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n530), .A2(new_n534), .A3(new_n537), .A4(new_n992), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT112), .ZN(new_n1005));
  AND2_X1   g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1006), .A2(new_n900), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1008), .B1(new_n895), .B2(new_n899), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n995), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1006), .A2(new_n900), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1008), .A2(new_n895), .A3(new_n899), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1011), .A2(new_n994), .A3(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1010), .A2(new_n968), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1015));
  INV_X1    g590(.A(new_n964), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT113), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT113), .ZN(new_n1018));
  AOI211_X1 g593(.A(new_n1018), .B(new_n964), .C1(new_n1010), .C2(new_n1013), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n985), .B(new_n1014), .C1(new_n1017), .C2(new_n1019), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n982), .A2(KEYINPUT110), .A3(new_n983), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT110), .B1(new_n982), .B2(new_n983), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n1011), .A2(new_n994), .A3(new_n1012), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n994), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1016), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1014), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(G37), .B1(new_n1023), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1020), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT114), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1020), .A2(new_n1028), .A3(KEYINPUT114), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1031), .A2(KEYINPUT43), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n1010), .A2(new_n968), .A3(new_n1013), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1026), .A2(new_n1018), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1015), .A2(KEYINPUT113), .A3(new_n1016), .ZN(new_n1038));
  AOI221_X4 g613(.A(new_n1036), .B1(new_n984), .B2(new_n979), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n985), .B1(new_n1040), .B2(new_n1014), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT43), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1042), .A2(new_n1043), .A3(new_n957), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1031), .A2(KEYINPUT115), .A3(KEYINPUT43), .A4(new_n1032), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1035), .A2(KEYINPUT44), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n1020), .A2(new_n1028), .A3(new_n1043), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1014), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n1023), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1049), .A2(new_n957), .A3(new_n1020), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1047), .B1(new_n1050), .B2(KEYINPUT43), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1046), .B1(KEYINPUT44), .B2(new_n1051), .ZN(G397));
  OR2_X1    g627(.A1(G290), .A2(G1986), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT117), .ZN(new_n1054));
  NAND2_X1  g629(.A1(G290), .A2(G1986), .ZN(new_n1055));
  XNOR2_X1  g630(.A(new_n1054), .B(new_n1055), .ZN(new_n1056));
  OR2_X1    g631(.A1(G164), .A2(G1384), .ZN(new_n1057));
  XOR2_X1   g632(.A(KEYINPUT116), .B(KEYINPUT45), .Z(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(G160), .A2(G40), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1056), .A2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n859), .B(new_n862), .ZN(new_n1064));
  INV_X1    g639(.A(G1996), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n844), .B(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  XOR2_X1   g642(.A(new_n755), .B(new_n758), .Z(new_n1068));
  OAI21_X1  g643(.A(new_n1062), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AND2_X1   g644(.A1(new_n1063), .A2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(G164), .A2(G1384), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT50), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G40), .ZN(new_n1074));
  AOI211_X1 g649(.A(new_n1074), .B(new_n469), .C1(new_n478), .C2(new_n479), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OR2_X1    g653(.A1(new_n1078), .A2(G1956), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1071), .A2(KEYINPUT45), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1060), .A2(new_n1075), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g657(.A(KEYINPUT56), .B(G2072), .ZN(new_n1083));
  XOR2_X1   g658(.A(new_n1083), .B(KEYINPUT120), .Z(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1079), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n1087));
  NAND2_X1  g662(.A1(G299), .A2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n1089));
  XOR2_X1   g664(.A(new_n1088), .B(new_n1089), .Z(new_n1090));
  OR2_X1    g665(.A1(new_n1086), .A2(new_n1090), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT118), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1093));
  OR3_X1    g668(.A1(new_n1071), .A2(KEYINPUT118), .A3(new_n1072), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n772), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1061), .A2(new_n1057), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n862), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1084), .ZN(new_n1100));
  OAI221_X1 g675(.A(new_n1090), .B1(new_n1081), .B2(new_n1100), .C1(new_n1078), .C2(G1956), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1099), .A2(new_n1101), .A3(new_n626), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT61), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1103), .A2(KEYINPUT123), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(KEYINPUT123), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1101), .A2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1079), .A2(new_n1085), .A3(new_n1090), .A4(new_n1105), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1104), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1110), .A2(KEYINPUT122), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1060), .A2(new_n1065), .A3(new_n1075), .A4(new_n1080), .ZN(new_n1112));
  XOR2_X1   g687(.A(KEYINPUT58), .B(G1341), .Z(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n1061), .B2(new_n1057), .ZN(new_n1114));
  AOI21_X1  g689(.A(KEYINPUT121), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1112), .A2(KEYINPUT121), .A3(new_n1114), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1116), .A2(new_n560), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1110), .A2(KEYINPUT122), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1111), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1111), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1117), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1122), .A2(new_n1115), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1121), .B1(new_n1123), .B2(new_n560), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1109), .B1(new_n1120), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT60), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1099), .A2(new_n1126), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1095), .A2(new_n772), .B1(new_n862), .B2(new_n1097), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT60), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1127), .A2(new_n626), .A3(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1128), .A2(KEYINPUT60), .A3(new_n625), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1091), .B(new_n1102), .C1(new_n1125), .C2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(G8), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1097), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n715), .A2(G1976), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT52), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n599), .B(G1981), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT49), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(new_n1135), .ZN(new_n1141));
  INV_X1    g716(.A(G1976), .ZN(new_n1142));
  AOI21_X1  g717(.A(KEYINPUT52), .B1(G288), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1135), .A2(new_n1136), .A3(new_n1143), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1138), .A2(new_n1141), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(G303), .A2(G8), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(KEYINPUT55), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  OAI22_X1  g723(.A1(new_n1095), .A2(G2090), .B1(new_n1082), .B2(G1971), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1148), .A2(G8), .A3(new_n1149), .ZN(new_n1150));
  AOI22_X1  g725(.A1(new_n1078), .A2(new_n827), .B1(new_n1081), .B2(new_n729), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1147), .B1(new_n1151), .B2(new_n1134), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1145), .A2(new_n1150), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT54), .ZN(new_n1154));
  XOR2_X1   g729(.A(KEYINPUT125), .B(G1961), .Z(new_n1155));
  NAND2_X1  g730(.A1(new_n1095), .A2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1060), .A2(new_n780), .A3(new_n1075), .A4(new_n1080), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT53), .ZN(new_n1158));
  OR2_X1    g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1156), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1161), .A2(G171), .ZN(new_n1162));
  OR2_X1    g737(.A1(new_n1071), .A2(KEYINPUT45), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1071), .A2(new_n1058), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1163), .A2(new_n780), .A3(new_n1075), .A4(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT124), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1158), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1164), .A2(new_n1075), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1071), .A2(KEYINPUT45), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1170), .A2(KEYINPUT124), .A3(new_n780), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1167), .A2(new_n1171), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1095), .A2(new_n1155), .B1(new_n1158), .B2(new_n1157), .ZN(new_n1173));
  AOI21_X1  g748(.A(G301), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1154), .B1(new_n1162), .B2(new_n1174), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1092), .A2(new_n828), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n809), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(G8), .B1(new_n1178), .B2(G286), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(KEYINPUT51), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT51), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1181), .B1(new_n1178), .B2(G286), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1180), .B1(new_n1182), .B2(new_n1179), .ZN(new_n1183));
  AND3_X1   g758(.A1(new_n1153), .A2(new_n1175), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1161), .A2(G171), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1172), .A2(new_n1173), .A3(G301), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1185), .A2(new_n1186), .A3(KEYINPUT54), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n1188));
  XNOR2_X1  g763(.A(new_n1187), .B(new_n1188), .ZN(new_n1189));
  AND3_X1   g764(.A1(new_n1133), .A2(new_n1184), .A3(new_n1189), .ZN(new_n1190));
  AOI211_X1 g765(.A(new_n1134), .B(G286), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1191));
  NAND4_X1  g766(.A1(new_n1145), .A2(new_n1150), .A3(new_n1152), .A4(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT63), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1149), .A2(G8), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1193), .B1(new_n1195), .B2(new_n1147), .ZN(new_n1196));
  NAND4_X1  g771(.A1(new_n1196), .A2(new_n1150), .A3(new_n1145), .A4(new_n1191), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1141), .A2(new_n1142), .A3(new_n715), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1198), .B1(G1981), .B2(new_n599), .ZN(new_n1199));
  AOI22_X1  g774(.A1(new_n1194), .A2(new_n1197), .B1(new_n1135), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1183), .A2(KEYINPUT62), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT62), .ZN(new_n1202));
  OAI211_X1 g777(.A(new_n1180), .B(new_n1202), .C1(new_n1182), .C2(new_n1179), .ZN(new_n1203));
  NAND4_X1  g778(.A1(new_n1201), .A2(new_n1153), .A3(new_n1174), .A4(new_n1203), .ZN(new_n1204));
  NAND4_X1  g779(.A1(new_n1145), .A2(G8), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1200), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1070), .B1(new_n1190), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n756), .A2(new_n758), .ZN(new_n1208));
  OAI22_X1  g783(.A1(new_n1067), .A2(new_n1208), .B1(G2067), .B2(new_n859), .ZN(new_n1209));
  AND2_X1   g784(.A1(new_n1209), .A2(new_n1062), .ZN(new_n1210));
  INV_X1    g785(.A(new_n1062), .ZN(new_n1211));
  AOI21_X1  g786(.A(new_n1211), .B1(new_n845), .B2(new_n1064), .ZN(new_n1212));
  AND3_X1   g787(.A1(new_n1062), .A2(KEYINPUT46), .A3(new_n1065), .ZN(new_n1213));
  AOI21_X1  g788(.A(KEYINPUT46), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1214));
  NOR3_X1   g789(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  XNOR2_X1  g790(.A(new_n1215), .B(KEYINPUT47), .ZN(new_n1216));
  NOR2_X1   g791(.A1(new_n1211), .A2(new_n1053), .ZN(new_n1217));
  XOR2_X1   g792(.A(new_n1217), .B(KEYINPUT48), .Z(new_n1218));
  AOI211_X1 g793(.A(new_n1210), .B(new_n1216), .C1(new_n1069), .C2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1207), .A2(new_n1219), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g795(.A1(G229), .A2(new_n459), .ZN(new_n1222));
  INV_X1    g796(.A(new_n1222), .ZN(new_n1223));
  NAND2_X1  g797(.A1(new_n1050), .A2(KEYINPUT43), .ZN(new_n1224));
  INV_X1    g798(.A(new_n1047), .ZN(new_n1225));
  AOI21_X1  g799(.A(new_n1223), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g800(.A(G227), .B1(new_n670), .B2(new_n674), .ZN(new_n1227));
  AND2_X1   g801(.A1(new_n958), .A2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g802(.A(KEYINPUT127), .B1(new_n1226), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g803(.A1(new_n958), .A2(new_n1227), .ZN(new_n1230));
  INV_X1    g804(.A(KEYINPUT127), .ZN(new_n1231));
  NOR4_X1   g805(.A1(new_n1051), .A2(new_n1230), .A3(new_n1231), .A4(new_n1223), .ZN(new_n1232));
  NOR2_X1   g806(.A1(new_n1229), .A2(new_n1232), .ZN(G308));
  AOI21_X1  g807(.A(new_n1043), .B1(new_n1042), .B2(new_n957), .ZN(new_n1234));
  OAI211_X1 g808(.A(new_n1222), .B(new_n1228), .C1(new_n1234), .C2(new_n1047), .ZN(new_n1235));
  NAND2_X1  g809(.A1(new_n1235), .A2(new_n1231), .ZN(new_n1236));
  NAND3_X1  g810(.A1(new_n1226), .A2(KEYINPUT127), .A3(new_n1228), .ZN(new_n1237));
  NAND2_X1  g811(.A1(new_n1236), .A2(new_n1237), .ZN(G225));
endmodule


