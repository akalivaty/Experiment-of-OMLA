//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 0 1 0 1 1 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 0 0 0 0 0 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955;
  INV_X1    g000(.A(G15gat), .ZN(new_n202));
  INV_X1    g001(.A(G22gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G15gat), .A2(G22gat), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT16), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(G8gat), .B1(new_n206), .B2(G1gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT16), .ZN(new_n208));
  INV_X1    g007(.A(new_n205), .ZN(new_n209));
  NOR2_X1   g008(.A1(G15gat), .A2(G22gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G1gat), .ZN(new_n212));
  INV_X1    g011(.A(G8gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n207), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n204), .A2(new_n205), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  OR2_X1    g016(.A1(new_n217), .A2(KEYINPUT90), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n217), .A2(KEYINPUT90), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n207), .A2(new_n220), .A3(new_n214), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT21), .ZN(new_n223));
  NAND2_X1  g022(.A1(G71gat), .A2(G78gat), .ZN(new_n224));
  XOR2_X1   g023(.A(new_n224), .B(KEYINPUT96), .Z(new_n225));
  OR2_X1    g024(.A1(G71gat), .A2(G78gat), .ZN(new_n226));
  INV_X1    g025(.A(G64gat), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n227), .A2(G57gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n227), .A2(G57gat), .ZN(new_n229));
  OAI22_X1  g028(.A1(new_n228), .A2(new_n229), .B1(KEYINPUT96), .B2(KEYINPUT9), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n225), .A2(new_n226), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT9), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n224), .B1(new_n226), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT97), .B(G57gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n234), .A2(new_n227), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n233), .B1(new_n235), .B2(new_n228), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n231), .A2(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n222), .B1(new_n223), .B2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n238), .B(G183gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(G231gat), .A2(G233gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G127gat), .B(G155gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(G211gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n241), .B(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n237), .A2(new_n223), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n245), .B(new_n246), .Z(new_n247));
  XNOR2_X1  g046(.A(new_n244), .B(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G43gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(G50gat), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT15), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n249), .A2(G50gat), .ZN(new_n253));
  NOR3_X1   g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G29gat), .ZN(new_n255));
  INV_X1    g054(.A(G36gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(new_n256), .A3(KEYINPUT14), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT14), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n258), .B1(G29gat), .B2(G36gat), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT89), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n257), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G29gat), .A2(G36gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n260), .B1(new_n257), .B2(new_n259), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n254), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT17), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n252), .B1(new_n251), .B2(new_n253), .ZN(new_n267));
  INV_X1    g066(.A(new_n253), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n268), .A2(new_n250), .A3(KEYINPUT15), .ZN(new_n269));
  AND2_X1   g068(.A1(new_n257), .A2(new_n259), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n267), .A2(new_n269), .A3(new_n270), .A4(new_n262), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n265), .A2(new_n266), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n266), .B1(new_n265), .B2(new_n271), .ZN(new_n274));
  XOR2_X1   g073(.A(G99gat), .B(G106gat), .Z(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(G85gat), .A2(G92gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT98), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT98), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n279), .A2(G85gat), .A3(G92gat), .ZN(new_n280));
  AND3_X1   g079(.A1(new_n278), .A2(new_n280), .A3(KEYINPUT7), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT7), .B1(new_n278), .B2(new_n280), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G99gat), .A2(G106gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT99), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT99), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n286), .A2(G99gat), .A3(G106gat), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n285), .A2(new_n287), .A3(KEYINPUT8), .ZN(new_n288));
  INV_X1    g087(.A(G85gat), .ZN(new_n289));
  INV_X1    g088(.A(G92gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n276), .B1(new_n283), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT7), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n279), .B1(G85gat), .B2(G92gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n277), .A2(KEYINPUT98), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n278), .A2(new_n280), .A3(KEYINPUT7), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n297), .A2(new_n291), .A3(new_n288), .A4(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n299), .A2(new_n275), .ZN(new_n300));
  OAI22_X1  g099(.A1(new_n273), .A2(new_n274), .B1(new_n293), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n300), .A2(new_n293), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n265), .A2(new_n271), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n301), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  XOR2_X1   g105(.A(G190gat), .B(G218gat), .Z(new_n307));
  XOR2_X1   g106(.A(new_n306), .B(new_n307), .Z(new_n308));
  XNOR2_X1  g107(.A(G134gat), .B(G162gat), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n309), .B(new_n310), .ZN(new_n311));
  OR3_X1    g110(.A1(new_n308), .A2(KEYINPUT100), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n308), .A2(new_n311), .ZN(new_n313));
  INV_X1    g112(.A(new_n307), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n306), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT100), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n312), .A2(new_n313), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n248), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G120gat), .B(G148gat), .ZN(new_n319));
  INV_X1    g118(.A(G176gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n319), .B(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(G204gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n321), .B(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT101), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n299), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n283), .A2(new_n292), .A3(KEYINPUT101), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n276), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT102), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n300), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT101), .B1(new_n283), .B2(new_n292), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n288), .A2(new_n291), .ZN(new_n332));
  NOR4_X1   g131(.A1(new_n332), .A2(new_n281), .A3(new_n282), .A4(new_n325), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n275), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT102), .ZN(new_n335));
  INV_X1    g134(.A(new_n237), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n330), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n237), .B1(new_n300), .B2(new_n293), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G230gat), .A2(G233gat), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT103), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT103), .ZN(new_n343));
  AOI211_X1 g142(.A(new_n343), .B(new_n340), .C1(new_n337), .C2(new_n338), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT10), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n337), .A2(new_n346), .A3(new_n338), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n303), .A2(KEYINPUT10), .A3(new_n336), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n340), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n324), .B1(new_n345), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n341), .B1(new_n347), .B2(new_n348), .ZN(new_n353));
  NOR3_X1   g152(.A1(new_n353), .A2(new_n342), .A3(new_n344), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT104), .B1(new_n354), .B2(new_n324), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n341), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(new_n343), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n339), .A2(KEYINPUT103), .A3(new_n341), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n350), .A2(new_n357), .A3(new_n324), .A4(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT104), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n352), .B1(new_n355), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT1), .ZN(new_n363));
  INV_X1    g162(.A(G120gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n364), .A2(G113gat), .ZN(new_n365));
  INV_X1    g164(.A(G113gat), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n366), .A2(G120gat), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n363), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  OR2_X1    g167(.A1(G127gat), .A2(G134gat), .ZN(new_n369));
  INV_X1    g168(.A(G134gat), .ZN(new_n370));
  XOR2_X1   g169(.A(KEYINPUT72), .B(G127gat), .Z(new_n371));
  OAI211_X1 g170(.A(new_n368), .B(new_n369), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  XOR2_X1   g171(.A(G141gat), .B(G148gat), .Z(new_n373));
  INV_X1    g172(.A(G155gat), .ZN(new_n374));
  INV_X1    g173(.A(G162gat), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT2), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G155gat), .B(G162gat), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(G127gat), .A2(G134gat), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT1), .B1(new_n369), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT73), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n383), .B1(new_n366), .B2(G120gat), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n364), .A2(KEYINPUT73), .A3(G113gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n382), .B1(new_n386), .B2(new_n365), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n373), .A2(new_n378), .A3(new_n376), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n372), .A2(new_n380), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT4), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n389), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT4), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n380), .A2(new_n388), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT3), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n372), .A2(new_n387), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT3), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n380), .A2(new_n397), .A3(new_n388), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n395), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(G225gat), .A2(G233gat), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n389), .A2(new_n401), .ZN(new_n402));
  AND4_X1   g201(.A1(new_n391), .A2(new_n393), .A3(new_n399), .A4(new_n402), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n372), .A2(new_n387), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n380), .A2(new_n388), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n401), .B1(new_n406), .B2(new_n392), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT5), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n393), .A2(new_n399), .A3(new_n391), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n401), .A2(KEYINPUT5), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  OAI22_X1  g210(.A1(new_n403), .A2(new_n408), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G1gat), .B(G29gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n413), .B(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(G57gat), .B(G85gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n412), .A2(KEYINPUT6), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n412), .A2(new_n418), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT6), .ZN(new_n421));
  OAI221_X1 g220(.A(new_n417), .B1(new_n409), .B2(new_n411), .C1(new_n403), .C2(new_n408), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT85), .ZN(new_n424));
  XNOR2_X1  g223(.A(G8gat), .B(G36gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(new_n227), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(new_n290), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(G183gat), .A2(G190gat), .ZN(new_n429));
  INV_X1    g228(.A(G169gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n320), .ZN(new_n431));
  NOR3_X1   g230(.A1(new_n431), .A2(KEYINPUT70), .A3(KEYINPUT26), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT70), .ZN(new_n433));
  NOR2_X1   g232(.A1(G169gat), .A2(G176gat), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT26), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OR2_X1    g235(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(G169gat), .A2(G176gat), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n438), .B1(new_n434), .B2(new_n435), .ZN(new_n439));
  OAI211_X1 g238(.A(KEYINPUT71), .B(new_n429), .C1(new_n437), .C2(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(KEYINPUT27), .B(G183gat), .ZN(new_n441));
  INV_X1    g240(.A(G190gat), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(KEYINPUT28), .A3(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT69), .B(G183gat), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT27), .ZN(new_n445));
  OR2_X1    g244(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n446));
  AOI21_X1  g245(.A(G190gat), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n443), .B1(new_n447), .B2(KEYINPUT28), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT71), .ZN(new_n449));
  NOR3_X1   g248(.A1(new_n432), .A2(new_n439), .A3(new_n436), .ZN(new_n450));
  INV_X1    g249(.A(new_n429), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n440), .A2(new_n448), .A3(new_n452), .ZN(new_n453));
  XOR2_X1   g252(.A(KEYINPUT69), .B(G183gat), .Z(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n442), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT24), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n429), .A2(new_n456), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n457), .A2(KEYINPUT68), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(KEYINPUT68), .ZN(new_n459));
  OR2_X1    g258(.A1(new_n456), .A2(KEYINPUT67), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n456), .A2(KEYINPUT67), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n429), .A3(new_n461), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n455), .A2(new_n458), .A3(new_n459), .A4(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT65), .B(KEYINPUT23), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(new_n431), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n434), .A2(KEYINPUT23), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n438), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n468), .B(KEYINPUT66), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT25), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n451), .A2(KEYINPUT24), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n429), .A2(new_n456), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n471), .B(new_n472), .C1(G183gat), .C2(G190gat), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT25), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(new_n474), .A3(new_n465), .ZN(new_n475));
  XOR2_X1   g274(.A(new_n467), .B(KEYINPUT64), .Z(new_n476));
  INV_X1    g275(.A(new_n438), .ZN(new_n477));
  OR3_X1    g276(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n453), .A2(new_n470), .A3(new_n478), .ZN(new_n479));
  XOR2_X1   g278(.A(KEYINPUT77), .B(KEYINPUT29), .Z(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(G226gat), .A2(G233gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NOR3_X1   g283(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n485));
  XOR2_X1   g284(.A(new_n468), .B(KEYINPUT66), .Z(new_n486));
  NAND3_X1  g285(.A1(new_n486), .A2(new_n463), .A3(new_n465), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n485), .B1(new_n487), .B2(KEYINPUT25), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n483), .B1(new_n488), .B2(new_n453), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(G211gat), .A2(G218gat), .ZN(new_n491));
  INV_X1    g290(.A(G211gat), .ZN(new_n492));
  INV_X1    g291(.A(G218gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT22), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n491), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(G197gat), .B(G204gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n498), .B(KEYINPUT76), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(KEYINPUT22), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n500), .A2(new_n491), .A3(new_n494), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n484), .A2(new_n490), .A3(new_n503), .ZN(new_n504));
  OR2_X1    g303(.A1(new_n499), .A2(new_n502), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT29), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n479), .A2(new_n506), .B1(G226gat), .B2(G233gat), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n505), .B1(new_n507), .B2(new_n489), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n428), .B1(new_n509), .B2(KEYINPUT38), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT85), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n420), .A2(new_n422), .A3(new_n511), .A4(new_n421), .ZN(new_n512));
  AND4_X1   g311(.A1(new_n419), .A2(new_n424), .A3(new_n510), .A4(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT37), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n509), .A2(new_n514), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT38), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n484), .A2(new_n490), .A3(new_n505), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT86), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n484), .A2(new_n490), .A3(KEYINPUT86), .A4(new_n505), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n503), .B1(new_n507), .B2(new_n489), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT37), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT38), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n525), .A2(new_n526), .A3(new_n427), .A4(new_n515), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n513), .A2(new_n518), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT78), .B1(new_n509), .B2(new_n428), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT78), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n504), .A2(new_n508), .A3(new_n530), .A4(new_n427), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT79), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n533), .A2(KEYINPUT30), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n509), .A2(new_n428), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(KEYINPUT30), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n509), .A2(new_n533), .A3(KEYINPUT30), .A4(new_n428), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n532), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n409), .A2(new_n401), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n406), .A2(new_n392), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n540), .B(KEYINPUT39), .C1(new_n401), .C2(new_n541), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n542), .B(new_n417), .C1(KEYINPUT39), .C2(new_n540), .ZN(new_n543));
  NOR2_X1   g342(.A1(KEYINPUT84), .A2(KEYINPUT40), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n543), .B(new_n544), .Z(new_n545));
  NAND3_X1  g344(.A1(new_n539), .A2(new_n420), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n398), .A2(new_n481), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n547), .A2(KEYINPUT81), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT81), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n549), .B1(new_n398), .B2(new_n481), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n503), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT82), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n397), .B1(new_n503), .B2(KEYINPUT29), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(new_n394), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT82), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n555), .B(new_n503), .C1(new_n548), .C2(new_n550), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n552), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(G228gat), .ZN(new_n558));
  INV_X1    g357(.A(G233gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n505), .A2(new_n481), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n405), .B1(new_n562), .B2(new_n397), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n503), .A2(new_n547), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n564), .B1(new_n558), .B2(new_n559), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(G22gat), .B1(new_n561), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(G78gat), .B(G106gat), .Z(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT31), .ZN(new_n571));
  INV_X1    g370(.A(G50gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT83), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n561), .A2(G22gat), .A3(new_n567), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n569), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n573), .A2(new_n574), .ZN(new_n578));
  AND3_X1   g377(.A1(new_n561), .A2(G22gat), .A3(new_n567), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n578), .B1(new_n579), .B2(new_n568), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n528), .A2(new_n546), .A3(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G15gat), .B(G43gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(G71gat), .B(G99gat), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n583), .B(new_n584), .Z(new_n585));
  NAND2_X1  g384(.A1(G227gat), .A2(G233gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n479), .A2(new_n396), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n488), .A2(new_n404), .A3(new_n453), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n585), .B1(new_n589), .B2(KEYINPUT33), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT32), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n587), .A2(new_n588), .A3(new_n586), .ZN(new_n594));
  INV_X1    g393(.A(new_n586), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT34), .B1(new_n595), .B2(KEYINPUT74), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n594), .B(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n587), .A2(new_n588), .ZN(new_n598));
  AOI221_X4 g397(.A(new_n591), .B1(KEYINPUT33), .B2(new_n585), .C1(new_n598), .C2(new_n595), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n593), .A2(new_n597), .A3(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n594), .B(new_n596), .Z(new_n602));
  NOR2_X1   g401(.A1(new_n590), .A2(new_n592), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n602), .B1(new_n603), .B2(new_n599), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n601), .A2(new_n604), .A3(KEYINPUT36), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n601), .A2(new_n604), .A3(KEYINPUT75), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT75), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n602), .B(new_n607), .C1(new_n603), .C2(new_n599), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n605), .B1(new_n609), .B2(KEYINPUT36), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n582), .A2(new_n610), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n577), .A2(new_n580), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n423), .A2(new_n419), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n532), .A2(new_n537), .A3(new_n613), .A4(new_n538), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n609), .A2(KEYINPUT87), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT35), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n424), .A2(new_n419), .A3(new_n512), .ZN(new_n618));
  AND3_X1   g417(.A1(new_n581), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n539), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT87), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n606), .A2(new_n621), .A3(new_n608), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n616), .A2(new_n619), .A3(new_n620), .A4(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n581), .A2(new_n604), .A3(new_n601), .ZN(new_n624));
  OAI21_X1  g423(.A(KEYINPUT35), .B1(new_n624), .B2(new_n614), .ZN(new_n625));
  AOI22_X1  g424(.A1(new_n611), .A2(new_n615), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT91), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n222), .B(new_n627), .C1(new_n273), .C2(new_n274), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n304), .A2(KEYINPUT17), .ZN(new_n629));
  AOI22_X1  g428(.A1(new_n629), .A2(new_n272), .B1(new_n221), .B2(new_n219), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n265), .A2(new_n271), .ZN(new_n631));
  OAI21_X1  g430(.A(KEYINPUT91), .B1(new_n222), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n628), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(G229gat), .A2(G233gat), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT18), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n635), .B1(KEYINPUT92), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n636), .A2(KEYINPUT92), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n222), .B(new_n631), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n634), .B(KEYINPUT93), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT13), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n633), .A2(new_n639), .A3(new_n637), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n641), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(G113gat), .B(G141gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(G169gat), .B(G197gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT12), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n648), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n654), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n641), .A2(new_n646), .A3(new_n647), .A4(new_n656), .ZN(new_n657));
  AND3_X1   g456(.A1(new_n655), .A2(KEYINPUT94), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT94), .B1(new_n655), .B2(new_n657), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT95), .B1(new_n626), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n623), .A2(new_n625), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n582), .A2(new_n610), .A3(new_n615), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT95), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n665), .A2(new_n666), .A3(new_n660), .ZN(new_n667));
  AOI211_X1 g466(.A(new_n318), .B(new_n362), .C1(new_n662), .C2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n613), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g470(.A1(new_n668), .A2(new_n539), .ZN(new_n672));
  NAND2_X1  g471(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n208), .A2(new_n213), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT42), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n672), .A2(KEYINPUT42), .A3(new_n673), .A4(new_n674), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n677), .B(new_n678), .C1(new_n213), .C2(new_n672), .ZN(G1325gat));
  NAND2_X1  g478(.A1(new_n616), .A2(new_n622), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(G15gat), .B1(new_n668), .B2(new_n681), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n682), .A2(KEYINPUT105), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(KEYINPUT105), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n610), .A2(new_n202), .ZN(new_n685));
  AOI22_X1  g484(.A1(new_n683), .A2(new_n684), .B1(new_n668), .B2(new_n685), .ZN(G1326gat));
  NAND2_X1  g485(.A1(new_n668), .A2(new_n612), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT43), .B(G22gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1327gat));
  NOR2_X1   g488(.A1(new_n248), .A2(new_n362), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n691), .B1(new_n662), .B2(new_n667), .ZN(new_n692));
  INV_X1    g491(.A(new_n317), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n694), .A2(G29gat), .A3(new_n613), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT45), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT45), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n615), .B(KEYINPUT106), .ZN(new_n699));
  AOI22_X1  g498(.A1(new_n611), .A2(new_n699), .B1(new_n623), .B2(new_n625), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n698), .B1(new_n700), .B2(new_n317), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n655), .A2(new_n657), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n665), .A2(KEYINPUT44), .A3(new_n693), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n701), .A2(new_n702), .A3(new_n690), .A4(new_n703), .ZN(new_n704));
  OR2_X1    g503(.A1(new_n704), .A2(new_n613), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n697), .B1(new_n705), .B2(G29gat), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n696), .B1(new_n706), .B2(new_n695), .ZN(G1328gat));
  NOR3_X1   g506(.A1(new_n694), .A2(G36gat), .A3(new_n620), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT46), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(G36gat), .B1(new_n704), .B2(new_n620), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n708), .A2(new_n709), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(G1329gat));
  OAI21_X1  g512(.A(G43gat), .B1(new_n704), .B2(new_n610), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n692), .A2(new_n249), .A3(new_n681), .A4(new_n693), .ZN(new_n715));
  OAI211_X1 g514(.A(new_n714), .B(new_n715), .C1(KEYINPUT107), .C2(KEYINPUT47), .ZN(new_n716));
  NAND2_X1  g515(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(G1330gat));
  INV_X1    g517(.A(KEYINPUT48), .ZN(new_n719));
  OAI21_X1  g518(.A(G50gat), .B1(new_n704), .B2(new_n581), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n692), .A2(new_n572), .A3(new_n612), .A4(new_n693), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT108), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n722), .B1(new_n720), .B2(new_n721), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n719), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n720), .A2(new_n721), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(KEYINPUT108), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n727), .A2(KEYINPUT48), .A3(new_n728), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n725), .A2(new_n729), .ZN(G1331gat));
  NAND2_X1  g529(.A1(new_n359), .A2(new_n360), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n345), .A2(KEYINPUT104), .A3(new_n324), .A4(new_n350), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n351), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NOR4_X1   g532(.A1(new_n700), .A2(new_n702), .A3(new_n318), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n669), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(new_n234), .ZN(G1332gat));
  NAND2_X1  g535(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n734), .A2(new_n539), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT109), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n739), .B(new_n740), .Z(G1333gat));
  XNOR2_X1  g540(.A(new_n680), .B(KEYINPUT110), .ZN(new_n742));
  AOI21_X1  g541(.A(G71gat), .B1(new_n734), .B2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n610), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n744), .A2(G71gat), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n743), .B1(new_n734), .B2(new_n745), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g546(.A1(new_n734), .A2(new_n612), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(G78gat), .ZN(G1335gat));
  INV_X1    g548(.A(new_n248), .ZN(new_n750));
  INV_X1    g549(.A(new_n702), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n701), .A2(new_n362), .A3(new_n703), .A4(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(G85gat), .B1(new_n754), .B2(new_n613), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n611), .A2(new_n699), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n663), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n757), .A2(new_n693), .A3(new_n753), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n362), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n669), .A2(new_n289), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n755), .B1(new_n762), .B2(new_n763), .ZN(G1336gat));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n620), .A2(new_n733), .A3(G92gat), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT111), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(new_n760), .B2(new_n761), .ZN(new_n769));
  OAI21_X1  g568(.A(G92gat), .B1(new_n754), .B2(new_n620), .ZN(new_n770));
  XNOR2_X1  g569(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT112), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n759), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n758), .A2(new_n775), .A3(KEYINPUT51), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n777), .A2(new_n768), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n774), .B1(new_n779), .B2(new_n770), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n765), .B1(new_n773), .B2(new_n780), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n779), .A2(new_n770), .ZN(new_n782));
  OAI211_X1 g581(.A(KEYINPUT114), .B(new_n772), .C1(new_n782), .C2(new_n774), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(G1337gat));
  OAI21_X1  g583(.A(G99gat), .B1(new_n754), .B2(new_n610), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n680), .A2(G99gat), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n762), .B2(new_n786), .ZN(G1338gat));
  NOR2_X1   g586(.A1(new_n581), .A2(G106gat), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n777), .A2(new_n362), .A3(new_n778), .A4(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(G106gat), .B1(new_n754), .B2(new_n581), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT53), .ZN(new_n792));
  XNOR2_X1  g591(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n793));
  INV_X1    g592(.A(new_n788), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n790), .B(new_n793), .C1(new_n762), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n792), .A2(new_n795), .ZN(G1339gat));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n349), .A2(new_n797), .A3(new_n340), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n323), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT116), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n347), .A2(new_n800), .A3(new_n341), .A4(new_n348), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT54), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n347), .A2(new_n341), .A3(new_n348), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n804), .B1(new_n353), .B2(KEYINPUT116), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n799), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  AOI22_X1  g605(.A1(new_n806), .A2(KEYINPUT55), .B1(new_n731), .B2(new_n732), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT117), .B1(new_n806), .B2(KEYINPUT55), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n350), .A2(new_n800), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n802), .B1(new_n811), .B2(new_n804), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n809), .B(new_n810), .C1(new_n812), .C2(new_n799), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n807), .A2(new_n808), .A3(new_n702), .A4(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n633), .ZN(new_n815));
  AOI22_X1  g614(.A1(new_n815), .A2(new_n635), .B1(new_n643), .B2(new_n645), .ZN(new_n816));
  OR2_X1    g615(.A1(new_n816), .A2(new_n653), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n657), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n362), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n693), .B1(new_n814), .B2(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n807), .A2(new_n808), .A3(new_n813), .A4(new_n819), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n822), .A2(new_n317), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n750), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n318), .A2(new_n702), .A3(new_n362), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n624), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n539), .A2(new_n613), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n829), .A2(new_n366), .A3(new_n702), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n824), .A2(new_n826), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n612), .A2(new_n613), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n831), .A2(new_n620), .A3(new_n681), .A4(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(G113gat), .B1(new_n833), .B2(new_n661), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n830), .A2(new_n834), .ZN(G1340gat));
  NAND3_X1  g634(.A1(new_n829), .A2(new_n364), .A3(new_n362), .ZN(new_n836));
  OAI21_X1  g635(.A(G120gat), .B1(new_n833), .B2(new_n733), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(G1341gat));
  NOR3_X1   g637(.A1(new_n833), .A2(new_n371), .A3(new_n750), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n829), .A2(new_n248), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n839), .B1(new_n840), .B2(new_n371), .ZN(G1342gat));
  NAND3_X1  g640(.A1(new_n829), .A2(new_n370), .A3(new_n693), .ZN(new_n842));
  XOR2_X1   g641(.A(new_n842), .B(KEYINPUT56), .Z(new_n843));
  OAI21_X1  g642(.A(G134gat), .B1(new_n833), .B2(new_n317), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(G1343gat));
  NAND2_X1  g644(.A1(new_n806), .A2(KEYINPUT55), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n810), .B1(new_n812), .B2(new_n799), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n731), .A2(new_n732), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n660), .A2(new_n846), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n362), .A2(new_n850), .A3(new_n819), .ZN(new_n851));
  OAI21_X1  g650(.A(KEYINPUT118), .B1(new_n733), .B2(new_n818), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n849), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n317), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n822), .A2(new_n317), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n248), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n612), .B1(new_n856), .B2(new_n825), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(KEYINPUT57), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n610), .A2(new_n828), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n581), .B1(new_n824), .B2(new_n826), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n858), .A2(new_n860), .A3(new_n863), .ZN(new_n864));
  OR3_X1    g663(.A1(new_n864), .A2(KEYINPUT119), .A3(new_n661), .ZN(new_n865));
  OAI21_X1  g664(.A(KEYINPUT119), .B1(new_n864), .B2(new_n661), .ZN(new_n866));
  AND3_X1   g665(.A1(new_n865), .A2(G141gat), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n861), .A2(new_n860), .ZN(new_n868));
  OR3_X1    g667(.A1(new_n868), .A2(G141gat), .A3(new_n661), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT58), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(G141gat), .B1(new_n864), .B2(new_n751), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n872), .A2(new_n869), .ZN(new_n873));
  OAI22_X1  g672(.A1(new_n867), .A2(new_n871), .B1(new_n870), .B2(new_n873), .ZN(G1344gat));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n875), .B(G148gat), .C1(new_n864), .C2(new_n733), .ZN(new_n876));
  XNOR2_X1  g675(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n831), .A2(new_n612), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(KEYINPUT57), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n318), .A2(new_n660), .A3(new_n362), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n862), .B(new_n612), .C1(new_n856), .C2(new_n880), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n879), .A2(new_n362), .A3(new_n860), .A4(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n877), .B1(new_n882), .B2(G148gat), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI211_X1 g684(.A(KEYINPUT121), .B(new_n877), .C1(new_n882), .C2(G148gat), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n876), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n733), .A2(G148gat), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n887), .B1(new_n868), .B2(new_n888), .ZN(G1345gat));
  INV_X1    g688(.A(new_n868), .ZN(new_n890));
  AOI21_X1  g689(.A(G155gat), .B1(new_n890), .B2(new_n248), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n864), .A2(new_n750), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n891), .B1(new_n892), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g692(.A(G162gat), .B1(new_n890), .B2(new_n693), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n864), .A2(new_n375), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n894), .B1(new_n895), .B2(new_n693), .ZN(G1347gat));
  NOR2_X1   g695(.A1(new_n620), .A2(new_n669), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n827), .A2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n899), .A2(new_n430), .A3(new_n702), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n897), .B(KEYINPUT122), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n831), .A2(new_n581), .A3(new_n742), .A4(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(G169gat), .B1(new_n903), .B2(new_n661), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n900), .A2(new_n904), .ZN(G1348gat));
  NOR3_X1   g704(.A1(new_n903), .A2(new_n320), .A3(new_n733), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n899), .A2(new_n362), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(new_n320), .B2(new_n907), .ZN(G1349gat));
  OAI21_X1  g707(.A(new_n444), .B1(new_n903), .B2(new_n750), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n248), .A2(new_n441), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n898), .B2(new_n910), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g711(.A1(new_n899), .A2(new_n442), .A3(new_n693), .ZN(new_n913));
  OAI21_X1  g712(.A(G190gat), .B1(new_n903), .B2(new_n317), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n914), .A2(KEYINPUT61), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n914), .A2(KEYINPUT61), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n913), .B1(new_n915), .B2(new_n916), .ZN(G1351gat));
  NOR2_X1   g716(.A1(new_n901), .A2(new_n744), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n881), .B(new_n918), .C1(new_n862), .C2(new_n861), .ZN(new_n919));
  OAI21_X1  g718(.A(G197gat), .B1(new_n919), .B2(new_n661), .ZN(new_n920));
  AND3_X1   g719(.A1(new_n861), .A2(new_n610), .A3(new_n897), .ZN(new_n921));
  INV_X1    g720(.A(G197gat), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n921), .A2(new_n922), .A3(new_n702), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  XOR2_X1   g723(.A(new_n924), .B(KEYINPUT123), .Z(G1352gat));
  NAND3_X1  g724(.A1(new_n921), .A2(new_n322), .A3(new_n362), .ZN(new_n926));
  XOR2_X1   g725(.A(new_n926), .B(KEYINPUT62), .Z(new_n927));
  INV_X1    g726(.A(KEYINPUT124), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n879), .A2(new_n362), .A3(new_n881), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n322), .B1(new_n930), .B2(new_n918), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n927), .A2(new_n928), .A3(new_n932), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n926), .B(KEYINPUT62), .ZN(new_n934));
  OAI21_X1  g733(.A(KEYINPUT124), .B1(new_n934), .B2(new_n931), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n935), .ZN(G1353gat));
  NAND3_X1  g735(.A1(new_n921), .A2(new_n492), .A3(new_n248), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n879), .A2(new_n248), .A3(new_n881), .A4(new_n918), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n938), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n939));
  AOI21_X1  g738(.A(KEYINPUT63), .B1(new_n938), .B2(G211gat), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI211_X1 g742(.A(KEYINPUT125), .B(new_n937), .C1(new_n939), .C2(new_n940), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1354gat));
  INV_X1    g744(.A(KEYINPUT126), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n919), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n879), .A2(KEYINPUT126), .A3(new_n881), .A4(new_n918), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n947), .A2(new_n693), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(G218gat), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n921), .A2(new_n493), .A3(new_n693), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT127), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n950), .A2(KEYINPUT127), .A3(new_n951), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1355gat));
endmodule


