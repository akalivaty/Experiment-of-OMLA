//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993;
  XNOR2_X1  g000(.A(KEYINPUT2), .B(G113), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT69), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT69), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n189), .A2(new_n191), .A3(G116), .ZN(new_n192));
  OR2_X1    g006(.A1(new_n188), .A2(G116), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(KEYINPUT70), .A3(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  AOI21_X1  g009(.A(KEYINPUT70), .B1(new_n192), .B2(new_n193), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n187), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n192), .A2(new_n193), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(new_n187), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n202));
  AND2_X1   g016(.A1(KEYINPUT0), .A2(G128), .ZN(new_n203));
  NOR2_X1   g017(.A1(KEYINPUT0), .A2(G128), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT64), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G143), .ZN(new_n209));
  AOI21_X1  g023(.A(G146), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(G143), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n202), .B(new_n205), .C1(new_n210), .C2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(G143), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n207), .A2(new_n209), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n203), .B(new_n214), .C1(new_n215), .C2(new_n211), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n212), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT64), .B(G143), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n218), .B1(new_n219), .B2(G146), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n202), .B1(new_n220), .B2(new_n205), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G131), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT11), .ZN(new_n225));
  INV_X1    g039(.A(G137), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n224), .A2(new_n225), .A3(new_n226), .A4(G134), .ZN(new_n227));
  INV_X1    g041(.A(G134), .ZN(new_n228));
  OAI22_X1  g042(.A1(new_n228), .A2(G137), .B1(KEYINPUT66), .B2(KEYINPUT11), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n228), .A2(G137), .B1(KEYINPUT66), .B2(KEYINPUT11), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n223), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  OAI22_X1  g047(.A1(new_n224), .A2(new_n225), .B1(new_n226), .B2(G134), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n234), .B1(new_n229), .B2(new_n227), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(new_n223), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n222), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G128), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(KEYINPUT1), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n214), .B(new_n240), .C1(new_n215), .C2(new_n211), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n212), .B1(new_n215), .B2(new_n211), .ZN(new_n242));
  OR2_X1    g056(.A1(KEYINPUT68), .A2(G128), .ZN(new_n243));
  NAND2_X1  g057(.A1(KEYINPUT68), .A2(G128), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n243), .A2(new_n244), .B1(new_n214), .B2(KEYINPUT1), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n241), .B1(new_n242), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n226), .A2(G134), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n228), .A2(G137), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n223), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n249), .B1(new_n235), .B2(new_n223), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n238), .A2(KEYINPUT30), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n251), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT67), .ZN(new_n254));
  INV_X1    g068(.A(new_n205), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT65), .B1(new_n242), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(new_n213), .A3(new_n216), .ZN(new_n257));
  AND3_X1   g071(.A1(new_n230), .A2(new_n223), .A3(new_n231), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n258), .A2(new_n232), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n254), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n213), .A2(new_n216), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n237), .A2(new_n261), .A3(KEYINPUT67), .A4(new_n256), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n253), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n201), .B(new_n252), .C1(new_n263), .C2(KEYINPUT30), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n251), .B1(new_n257), .B2(new_n259), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(new_n201), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G237), .ZN(new_n268));
  INV_X1    g082(.A(G953), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n268), .A2(new_n269), .A3(G210), .ZN(new_n270));
  XOR2_X1   g084(.A(new_n270), .B(KEYINPUT27), .Z(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT26), .B(G101), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n271), .B(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n264), .A2(new_n267), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT31), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n264), .A2(KEYINPUT31), .A3(new_n267), .A4(new_n274), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n265), .A2(KEYINPUT71), .ZN(new_n280));
  INV_X1    g094(.A(new_n201), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT71), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n282), .B(new_n251), .C1(new_n257), .C2(new_n259), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n280), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT28), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT67), .B1(new_n222), .B2(new_n237), .ZN(new_n287));
  NOR3_X1   g101(.A1(new_n257), .A2(new_n254), .A3(new_n259), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n251), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n266), .B1(new_n289), .B2(new_n201), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n286), .B1(new_n290), .B2(new_n285), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n273), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n279), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(G472), .A2(G902), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(KEYINPUT32), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT32), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n277), .A2(new_n278), .B1(new_n291), .B2(new_n273), .ZN(new_n297));
  INV_X1    g111(.A(new_n294), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n264), .A2(new_n267), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n273), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n286), .B(new_n274), .C1(new_n290), .C2(new_n285), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT29), .ZN(new_n303));
  AND3_X1   g117(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n281), .B1(new_n238), .B2(new_n251), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT28), .B1(new_n305), .B2(new_n266), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n273), .A2(new_n303), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n286), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT72), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G902), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n286), .A2(new_n306), .A3(KEYINPUT72), .A4(new_n307), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(G472), .B1(new_n304), .B2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n295), .A2(new_n299), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G217), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n317), .B1(G234), .B2(new_n311), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT75), .ZN(new_n319));
  XNOR2_X1  g133(.A(G125), .B(G140), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT16), .ZN(new_n321));
  INV_X1    g135(.A(G140), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G125), .ZN(new_n323));
  OR2_X1    g137(.A1(new_n323), .A2(KEYINPUT16), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n321), .A2(G146), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G125), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G140), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n329), .A2(G146), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n189), .A2(new_n191), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n331), .A2(new_n239), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n243), .A2(G119), .A3(new_n244), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT23), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G110), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT23), .ZN(new_n336));
  INV_X1    g150(.A(new_n331), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n336), .B1(new_n337), .B2(G128), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n334), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT24), .B(G110), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n340), .B1(new_n332), .B2(new_n333), .ZN(new_n341));
  AOI211_X1 g155(.A(new_n326), .B(new_n330), .C1(new_n339), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n321), .A2(new_n324), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n211), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n325), .ZN(new_n345));
  OR3_X1    g159(.A1(new_n332), .A2(new_n333), .A3(new_n340), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n335), .B1(new_n334), .B2(new_n338), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n319), .B1(new_n342), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n348), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(new_n346), .A3(new_n345), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n339), .A2(new_n341), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n326), .A2(new_n330), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n352), .A2(new_n355), .A3(KEYINPUT75), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT22), .B(G137), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n269), .A2(G221), .A3(G234), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n357), .B(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n359), .B(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n350), .A2(new_n356), .A3(new_n362), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n352), .A2(new_n355), .A3(KEYINPUT75), .A4(new_n361), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT25), .B1(new_n365), .B2(new_n311), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT25), .ZN(new_n367));
  AOI211_X1 g181(.A(new_n367), .B(G902), .C1(new_n363), .C2(new_n364), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n318), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT76), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT76), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n371), .B(new_n318), .C1(new_n366), .C2(new_n368), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n318), .A2(G902), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n365), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n370), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n316), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(KEYINPUT9), .B(G234), .ZN(new_n377));
  OAI21_X1  g191(.A(G221), .B1(new_n377), .B2(G902), .ZN(new_n378));
  XOR2_X1   g192(.A(new_n378), .B(KEYINPUT77), .Z(new_n379));
  INV_X1    g193(.A(G469), .ZN(new_n380));
  XNOR2_X1  g194(.A(G110), .B(G140), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(KEYINPUT78), .ZN(new_n382));
  AND2_X1   g196(.A1(new_n269), .A2(G227), .ZN(new_n383));
  XOR2_X1   g197(.A(new_n382), .B(new_n383), .Z(new_n384));
  INV_X1    g198(.A(KEYINPUT81), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT80), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT4), .ZN(new_n387));
  INV_X1    g201(.A(G104), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT3), .B1(new_n388), .B2(G107), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT3), .ZN(new_n390));
  INV_X1    g204(.A(G107), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n391), .A3(G104), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n388), .A2(G107), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n389), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT79), .B(G101), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n387), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n389), .A2(new_n392), .A3(new_n393), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G101), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n386), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n395), .A2(new_n392), .A3(new_n389), .A4(new_n393), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n398), .A2(new_n386), .A3(new_n400), .A4(KEYINPUT4), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n398), .A2(KEYINPUT4), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n261), .A2(new_n405), .A3(new_n256), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n385), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT10), .ZN(new_n408));
  INV_X1    g222(.A(new_n241), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT83), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT1), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n410), .B1(new_n210), .B2(new_n411), .ZN(new_n412));
  OAI211_X1 g226(.A(KEYINPUT83), .B(KEYINPUT1), .C1(new_n219), .C2(G146), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(G128), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n214), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n415), .B1(new_n219), .B2(G146), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n409), .B1(new_n414), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n391), .A2(G104), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(new_n393), .A3(KEYINPUT82), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n420), .B(G101), .C1(KEYINPUT82), .C2(new_n419), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n400), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n408), .B1(new_n418), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n422), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(KEYINPUT10), .A3(new_n246), .ZN(new_n425));
  NOR3_X1   g239(.A1(new_n217), .A2(new_n404), .A3(new_n221), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n398), .A2(KEYINPUT4), .A3(new_n400), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT80), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n401), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n426), .A2(new_n429), .A3(KEYINPUT81), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n407), .A2(new_n423), .A3(new_n425), .A4(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(KEYINPUT84), .B1(new_n431), .B2(new_n237), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n426), .A2(new_n429), .A3(KEYINPUT81), .ZN(new_n433));
  AOI21_X1  g247(.A(KEYINPUT81), .B1(new_n426), .B2(new_n429), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n423), .A2(new_n425), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT84), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n435), .A2(new_n436), .A3(new_n437), .A4(new_n259), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n432), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n259), .B1(new_n435), .B2(new_n436), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n384), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n384), .ZN(new_n443));
  OR2_X1    g257(.A1(new_n242), .A2(new_n245), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(new_n241), .A3(new_n422), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n445), .B1(new_n418), .B2(new_n422), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n446), .A2(KEYINPUT12), .A3(new_n237), .ZN(new_n447));
  AOI21_X1  g261(.A(KEYINPUT12), .B1(new_n446), .B2(new_n237), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI211_X1 g263(.A(new_n443), .B(new_n449), .C1(new_n432), .C2(new_n438), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n380), .B(new_n311), .C1(new_n442), .C2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT86), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n439), .A2(new_n384), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n440), .B1(new_n432), .B2(new_n438), .ZN(new_n454));
  OAI22_X1  g268(.A1(new_n453), .A2(new_n449), .B1(new_n454), .B2(new_n384), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT86), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n455), .A2(new_n456), .A3(new_n380), .A4(new_n311), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n449), .B1(new_n432), .B2(new_n438), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n459), .A2(new_n384), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT85), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n453), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n443), .B1(new_n432), .B2(new_n438), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n440), .B1(new_n463), .B2(KEYINPUT85), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n460), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(G469), .B1(new_n465), .B2(G902), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n379), .B1(new_n458), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT90), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n320), .A2(KEYINPUT19), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n320), .A2(KEYINPUT19), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n211), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n268), .A2(new_n269), .A3(G214), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n219), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n268), .A2(new_n269), .A3(G143), .A4(G214), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n473), .A2(new_n223), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n223), .B1(new_n473), .B2(new_n474), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n471), .B(new_n325), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n473), .A2(new_n474), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(KEYINPUT18), .A3(G131), .ZN(new_n479));
  NAND2_X1  g293(.A1(KEYINPUT18), .A2(G131), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n473), .A2(new_n474), .A3(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n320), .B(new_n211), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n479), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT89), .ZN(new_n485));
  XNOR2_X1  g299(.A(G113), .B(G122), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(new_n388), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n484), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n476), .A2(KEYINPUT17), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(new_n344), .A3(new_n325), .ZN(new_n491));
  NOR3_X1   g305(.A1(new_n475), .A2(new_n476), .A3(KEYINPUT17), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n487), .B(new_n483), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n485), .B1(new_n484), .B2(new_n488), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n468), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(G475), .A2(G902), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n484), .A2(new_n488), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(KEYINPUT89), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n499), .A2(KEYINPUT90), .A3(new_n493), .A4(new_n489), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n496), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT20), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n499), .A2(new_n493), .A3(new_n489), .ZN(new_n503));
  NOR3_X1   g317(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n483), .B1(new_n491), .B2(new_n492), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n488), .ZN(new_n508));
  AOI21_X1  g322(.A(G902), .B1(new_n508), .B2(new_n493), .ZN(new_n509));
  INV_X1    g323(.A(G475), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(G116), .B(G122), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT14), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(G122), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n517), .A2(G116), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n391), .B1(new_n518), .B2(KEYINPUT14), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n516), .A2(new_n519), .B1(new_n391), .B2(new_n514), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n243), .A2(G143), .A3(new_n244), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n207), .A2(new_n209), .A3(G128), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n521), .A2(new_n522), .A3(new_n228), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n228), .B1(new_n521), .B2(new_n522), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n520), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n243), .A2(new_n244), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT13), .ZN(new_n528));
  AOI22_X1  g342(.A1(new_n527), .A2(G143), .B1(new_n522), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n219), .A2(KEYINPUT13), .A3(G128), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n228), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n514), .B(new_n391), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n523), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n526), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NOR3_X1   g348(.A1(new_n377), .A2(new_n317), .A3(G953), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n535), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n526), .B(new_n537), .C1(new_n531), .C2(new_n533), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n536), .A2(new_n311), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(G478), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n540), .A2(KEYINPUT15), .ZN(new_n541));
  XOR2_X1   g355(.A(new_n539), .B(new_n541), .Z(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n513), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(G234), .A2(G237), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(G952), .A3(new_n269), .ZN(new_n546));
  XOR2_X1   g360(.A(new_n546), .B(KEYINPUT91), .Z(new_n547));
  AND3_X1   g361(.A1(new_n545), .A2(G902), .A3(G953), .ZN(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT21), .B(G898), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(G214), .B1(G237), .B2(G902), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n404), .B1(new_n197), .B2(new_n200), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n429), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT70), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n198), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n557), .A2(KEYINPUT5), .A3(new_n194), .ZN(new_n558));
  OAI21_X1  g372(.A(G113), .B1(new_n192), .B2(KEYINPUT5), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n199), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n424), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n555), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(G110), .B(G122), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g380(.A1(new_n554), .A2(new_n429), .B1(new_n561), .B2(new_n424), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n564), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n566), .A2(new_n568), .A3(KEYINPUT6), .ZN(new_n569));
  OR3_X1    g383(.A1(new_n567), .A2(KEYINPUT6), .A3(new_n564), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n257), .A2(G125), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n444), .A2(new_n327), .A3(new_n241), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(G224), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n574), .A2(G953), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n573), .B(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n569), .A2(new_n570), .A3(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT87), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n571), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(KEYINPUT7), .B1(new_n574), .B2(G953), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n573), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n580), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n571), .B(new_n572), .C1(new_n578), .C2(new_n582), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n561), .A2(new_n422), .ZN(new_n585));
  XOR2_X1   g399(.A(new_n564), .B(KEYINPUT8), .Z(new_n586));
  AND3_X1   g400(.A1(new_n192), .A2(KEYINPUT5), .A3(new_n193), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n200), .B1(new_n587), .B2(new_n559), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n586), .B1(new_n588), .B2(new_n424), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n567), .A2(new_n564), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(G902), .B1(new_n584), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n577), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(G210), .B1(G237), .B2(G902), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n577), .A2(new_n591), .A3(new_n593), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n553), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT88), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT88), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n551), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n376), .A2(new_n467), .A3(new_n544), .A4(new_n602), .ZN(new_n603));
  XOR2_X1   g417(.A(new_n603), .B(new_n395), .Z(G3));
  AOI21_X1  g418(.A(new_n298), .B1(new_n279), .B2(new_n292), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(G472), .B1(new_n297), .B2(G902), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n608), .A2(new_n375), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n467), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(new_n610), .B(KEYINPUT92), .Z(new_n611));
  NAND2_X1  g425(.A1(new_n311), .A2(G478), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n535), .A2(KEYINPUT94), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n534), .A2(new_n613), .ZN(new_n614));
  OAI221_X1 g428(.A(new_n526), .B1(KEYINPUT94), .B2(new_n535), .C1(new_n531), .C2(new_n533), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n614), .A2(new_n615), .A3(KEYINPUT33), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT33), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n536), .A2(new_n618), .A3(new_n538), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT93), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT93), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n536), .A2(new_n621), .A3(new_n618), .A4(new_n538), .ZN(new_n622));
  AOI211_X1 g436(.A(new_n612), .B(new_n617), .C1(new_n620), .C2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT95), .B(G478), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n539), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT96), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(KEYINPUT96), .B1(new_n539), .B2(new_n624), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g443(.A(KEYINPUT97), .B1(new_n623), .B2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n625), .B(new_n626), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n620), .A2(new_n622), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n632), .A2(G478), .A3(new_n616), .A4(new_n311), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT97), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n631), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n630), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n511), .B1(new_n502), .B2(new_n505), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n551), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n597), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n611), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT34), .B(G104), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  XNOR2_X1  g460(.A(new_n501), .B(KEYINPUT20), .ZN(new_n647));
  XOR2_X1   g461(.A(new_n511), .B(KEYINPUT98), .Z(new_n648));
  AND2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AND4_X1   g463(.A1(new_n543), .A2(new_n649), .A3(new_n641), .A4(new_n597), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n611), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT99), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT35), .B(G107), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  NAND2_X1  g468(.A1(new_n352), .A2(new_n355), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT100), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n361), .A2(KEYINPUT36), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n373), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n370), .A2(new_n372), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n661), .A2(new_n608), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n467), .A2(new_n602), .A3(new_n662), .A4(new_n544), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT37), .B(G110), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G12));
  INV_X1    g479(.A(G900), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n548), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT101), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n547), .ZN(new_n669));
  AND4_X1   g483(.A1(new_n543), .A2(new_n647), .A3(new_n648), .A4(new_n669), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n315), .A2(new_n597), .A3(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n467), .A2(new_n671), .A3(new_n660), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G128), .ZN(G30));
  XNOR2_X1  g487(.A(new_n669), .B(KEYINPUT39), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n467), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT102), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT40), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  NOR4_X1   g493(.A1(new_n660), .A2(new_n638), .A3(new_n542), .A4(new_n553), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n595), .A2(new_n596), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT38), .ZN(new_n682));
  OR2_X1    g496(.A1(new_n305), .A2(new_n266), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n311), .B1(new_n683), .B2(new_n274), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n273), .B1(new_n264), .B2(new_n267), .ZN(new_n685));
  OAI21_X1  g499(.A(G472), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n295), .A2(new_n299), .A3(new_n686), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n680), .A2(new_n682), .A3(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n678), .A2(new_n679), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(new_n215), .ZN(G45));
  AND3_X1   g504(.A1(new_n636), .A2(new_n513), .A3(new_n669), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n315), .A2(new_n597), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n467), .A2(new_n692), .A3(new_n660), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G146), .ZN(G48));
  INV_X1    g508(.A(new_n379), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n311), .B1(new_n442), .B2(new_n450), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(G469), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n458), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT103), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AOI22_X1  g514(.A1(new_n452), .A2(new_n457), .B1(G469), .B2(new_n696), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(KEYINPUT103), .A3(new_n695), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n700), .A2(new_n376), .A3(new_n643), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT41), .B(G113), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G15));
  NAND4_X1  g519(.A1(new_n700), .A2(new_n376), .A3(new_n650), .A4(new_n702), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT104), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G116), .ZN(G18));
  AOI221_X4 g526(.A(new_n379), .B1(G469), .B2(new_n696), .C1(new_n452), .C2(new_n457), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n315), .A2(new_n544), .A3(new_n641), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n713), .A2(new_n714), .A3(new_n597), .A4(new_n660), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G119), .ZN(G21));
  AOI21_X1  g530(.A(new_n274), .B1(new_n286), .B2(new_n306), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n717), .B1(new_n277), .B2(new_n278), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n607), .B1(new_n298), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(KEYINPUT105), .B1(new_n638), .B2(new_n542), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT105), .ZN(new_n721));
  AOI22_X1  g535(.A1(new_n501), .A2(KEYINPUT20), .B1(new_n503), .B2(new_n504), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n721), .B(new_n543), .C1(new_n722), .C2(new_n511), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  NOR4_X1   g538(.A1(new_n719), .A2(new_n724), .A3(new_n375), .A4(new_n642), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n700), .A2(new_n725), .A3(new_n702), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G122), .ZN(G24));
  NAND3_X1  g541(.A1(new_n636), .A2(new_n513), .A3(new_n669), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n719), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n713), .A2(new_n597), .A3(new_n660), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G125), .ZN(G27));
  NAND2_X1  g545(.A1(new_n458), .A2(new_n466), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n595), .A2(new_n552), .A3(new_n596), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT42), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n728), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n732), .A2(new_n695), .A3(new_n734), .A4(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n295), .A2(KEYINPUT108), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n605), .A2(new_n739), .A3(KEYINPUT32), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n738), .A2(new_n299), .A3(new_n314), .A4(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n741), .A2(new_n372), .A3(new_n370), .A4(new_n374), .ZN(new_n742));
  OAI21_X1  g556(.A(KEYINPUT109), .B1(new_n737), .B2(new_n742), .ZN(new_n743));
  AOI211_X1 g557(.A(new_n379), .B(new_n733), .C1(new_n458), .C2(new_n466), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT109), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n299), .A2(new_n314), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n739), .B1(new_n605), .B2(KEYINPUT32), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n375), .B1(new_n748), .B2(new_n740), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n744), .A2(new_n745), .A3(new_n749), .A4(new_n736), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n376), .A2(new_n467), .A3(new_n691), .A4(new_n734), .ZN(new_n751));
  XNOR2_X1  g565(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n751), .A2(KEYINPUT107), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(KEYINPUT107), .B1(new_n751), .B2(new_n752), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n743), .B(new_n750), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G131), .ZN(G33));
  NAND3_X1  g570(.A1(new_n744), .A2(new_n376), .A3(new_n670), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G134), .ZN(G36));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n636), .A2(new_n638), .ZN(new_n760));
  XOR2_X1   g574(.A(new_n760), .B(KEYINPUT43), .Z(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n660), .ZN(new_n762));
  INV_X1    g576(.A(new_n608), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n759), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n761), .A2(KEYINPUT44), .A3(new_n608), .A4(new_n660), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n764), .A2(new_n734), .A3(new_n765), .ZN(new_n766));
  OAI21_X1  g580(.A(G469), .B1(new_n465), .B2(KEYINPUT45), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n767), .B1(KEYINPUT45), .B2(new_n465), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n380), .A2(new_n311), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n770), .A2(KEYINPUT46), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(KEYINPUT46), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n458), .A3(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n766), .A2(new_n773), .A3(new_n695), .A4(new_n674), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G137), .ZN(G39));
  NAND2_X1  g589(.A1(new_n773), .A2(new_n695), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT47), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n773), .A2(KEYINPUT47), .A3(new_n695), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n691), .A2(new_n375), .A3(new_n734), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(new_n316), .A3(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G140), .ZN(G42));
  INV_X1    g597(.A(G952), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT115), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n786));
  AOI211_X1 g600(.A(G953), .B(new_n784), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n547), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n761), .A2(new_n788), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n719), .A2(new_n375), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n791), .A2(new_n598), .A3(new_n698), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n787), .B1(new_n792), .B2(KEYINPUT116), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n793), .B1(KEYINPUT116), .B2(new_n792), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n713), .A2(new_n734), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n789), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(new_n742), .ZN(new_n797));
  XOR2_X1   g611(.A(new_n797), .B(KEYINPUT48), .Z(new_n798));
  NOR4_X1   g612(.A1(new_n795), .A2(new_n375), .A3(new_n547), .A4(new_n687), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT114), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n639), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n794), .A2(new_n798), .A3(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n701), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n778), .B(new_n779), .C1(new_n695), .C2(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n791), .A2(new_n733), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR4_X1   g620(.A1(new_n791), .A2(new_n552), .A3(new_n682), .A4(new_n698), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(KEYINPUT50), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n800), .A2(new_n638), .A3(new_n637), .ZN(new_n809));
  OR3_X1    g623(.A1(new_n796), .A2(new_n661), .A3(new_n719), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n806), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n785), .A2(new_n786), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n802), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI22_X1  g628(.A1(new_n806), .A2(new_n811), .B1(new_n785), .B2(new_n786), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n817));
  AND4_X1   g631(.A1(new_n315), .A2(new_n542), .A3(new_n649), .A4(new_n669), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n744), .B(new_n660), .C1(new_n729), .C2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n757), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n720), .A2(new_n597), .A3(new_n723), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n370), .A2(new_n372), .A3(new_n659), .A4(new_n669), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n732), .A2(new_n823), .A3(new_n695), .A4(new_n687), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n730), .A2(new_n672), .A3(new_n693), .A4(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT52), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n467), .B(new_n660), .C1(new_n671), .C2(new_n692), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n828), .A2(KEYINPUT52), .A3(new_n730), .A4(new_n824), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n820), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n513), .A2(new_n542), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n467), .A2(new_n602), .A3(new_n609), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n663), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT110), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT110), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n663), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n467), .A2(new_n602), .A3(new_n609), .A4(new_n639), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n603), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT111), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n663), .A2(new_n832), .A3(new_n835), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n835), .B1(new_n663), .B2(new_n832), .ZN(new_n842));
  OAI211_X1 g656(.A(KEYINPUT111), .B(new_n839), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n830), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n703), .A2(new_n726), .A3(new_n715), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n846), .B1(new_n708), .B2(new_n710), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n755), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n817), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n827), .A2(new_n829), .ZN(new_n850));
  INV_X1    g664(.A(new_n820), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n839), .B1(new_n841), .B2(new_n842), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT111), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n852), .B1(new_n855), .B2(new_n843), .ZN(new_n856));
  INV_X1    g670(.A(new_n848), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n856), .A2(KEYINPUT53), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n849), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT54), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT112), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n847), .A2(new_n755), .A3(new_n861), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n703), .A2(new_n726), .A3(new_n715), .ZN(new_n863));
  INV_X1    g677(.A(new_n710), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n706), .A2(new_n709), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n743), .A2(new_n750), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n751), .A2(new_n752), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT107), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n751), .A2(KEYINPUT107), .A3(new_n752), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n867), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(KEYINPUT112), .B1(new_n866), .B2(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n856), .A2(KEYINPUT53), .A3(new_n862), .A4(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n874), .A2(new_n849), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n860), .A2(KEYINPUT113), .A3(new_n876), .ZN(new_n877));
  OR2_X1    g691(.A1(new_n876), .A2(KEYINPUT113), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n816), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(G952), .A2(G953), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT117), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n803), .A2(KEYINPUT49), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n636), .A2(new_n638), .A3(new_n695), .A4(new_n552), .ZN(new_n883));
  NOR4_X1   g697(.A1(new_n682), .A2(new_n687), .A3(new_n375), .A4(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT49), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n884), .B1(new_n885), .B2(new_n701), .ZN(new_n886));
  OAI22_X1  g700(.A1(new_n879), .A2(new_n881), .B1(new_n882), .B2(new_n886), .ZN(G75));
  NAND2_X1  g701(.A1(new_n784), .A2(G953), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n888), .B(KEYINPUT118), .Z(new_n889));
  NAND3_X1  g703(.A1(new_n873), .A2(KEYINPUT53), .A3(new_n862), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n890), .A2(new_n845), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT53), .B1(new_n856), .B2(new_n857), .ZN(new_n892));
  OAI211_X1 g706(.A(G210), .B(G902), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT56), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n569), .A2(new_n570), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n895), .B(new_n576), .Z(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT55), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n893), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n897), .B1(new_n893), .B2(new_n894), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n889), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT119), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI211_X1 g716(.A(KEYINPUT119), .B(new_n889), .C1(new_n898), .C2(new_n899), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(G51));
  XOR2_X1   g718(.A(new_n768), .B(KEYINPUT121), .Z(new_n905));
  AOI211_X1 g719(.A(new_n311), .B(new_n905), .C1(new_n874), .C2(new_n849), .ZN(new_n906));
  XNOR2_X1  g720(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(new_n769), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n874), .A2(new_n849), .A3(new_n875), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n875), .B1(new_n874), .B2(new_n849), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n906), .B1(new_n911), .B2(new_n455), .ZN(new_n912));
  INV_X1    g726(.A(new_n889), .ZN(new_n913));
  OAI21_X1  g727(.A(KEYINPUT122), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT122), .ZN(new_n915));
  INV_X1    g729(.A(new_n455), .ZN(new_n916));
  OAI21_X1  g730(.A(KEYINPUT54), .B1(new_n891), .B2(new_n892), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n876), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n916), .B1(new_n918), .B2(new_n908), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n915), .B(new_n889), .C1(new_n919), .C2(new_n906), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n914), .A2(new_n920), .ZN(G54));
  NAND2_X1  g735(.A1(new_n874), .A2(new_n849), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n922), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n496), .A2(new_n500), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  OR2_X1    g739(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n923), .A2(new_n925), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n913), .B1(new_n926), .B2(new_n927), .ZN(G60));
  INV_X1    g742(.A(new_n918), .ZN(new_n929));
  NAND2_X1  g743(.A1(G478), .A2(G902), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT59), .Z(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n632), .A2(new_n616), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n889), .B1(new_n929), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n877), .A2(new_n878), .A3(new_n932), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n632), .A2(new_n616), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(G63));
  NAND2_X1  g751(.A1(G217), .A2(G902), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT60), .Z(new_n939));
  AOI21_X1  g753(.A(new_n365), .B1(new_n922), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n940), .A2(new_n913), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT123), .ZN(new_n942));
  AOI21_X1  g756(.A(KEYINPUT61), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n658), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n922), .A2(new_n939), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n941), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  OAI221_X1 g761(.A(new_n941), .B1(new_n942), .B2(KEYINPUT61), .C1(new_n944), .C2(new_n945), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(G66));
  OAI21_X1  g763(.A(new_n847), .B1(new_n840), .B2(new_n844), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT124), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n269), .ZN(new_n952));
  OAI21_X1  g766(.A(G953), .B1(new_n549), .B2(new_n574), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n895), .B1(G898), .B2(new_n269), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n954), .B(new_n955), .ZN(G69));
  OAI21_X1  g770(.A(new_n252), .B1(new_n263), .B2(KEYINPUT30), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n469), .A2(new_n470), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT125), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n957), .B(new_n959), .ZN(new_n960));
  OAI211_X1 g774(.A(G900), .B(G953), .C1(new_n960), .C2(G227), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n961), .B1(G227), .B2(new_n960), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n828), .A2(new_n730), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n742), .A2(new_n821), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n773), .A2(new_n695), .A3(new_n674), .A4(new_n964), .ZN(new_n965));
  AND4_X1   g779(.A1(new_n757), .A2(new_n774), .A3(new_n963), .A4(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n782), .A2(new_n755), .A3(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(G953), .B1(new_n968), .B2(new_n960), .ZN(new_n969));
  INV_X1    g783(.A(new_n831), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n733), .B1(new_n640), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n676), .A2(new_n376), .A3(new_n971), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n774), .A2(new_n972), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n689), .A2(KEYINPUT62), .A3(new_n963), .ZN(new_n974));
  AOI21_X1  g788(.A(KEYINPUT62), .B1(new_n689), .B2(new_n963), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n782), .B(new_n973), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n960), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n962), .B1(new_n969), .B2(new_n978), .ZN(G72));
  NAND2_X1  g793(.A1(G472), .A2(G902), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT63), .Z(new_n981));
  OAI21_X1  g795(.A(new_n981), .B1(new_n951), .B2(new_n976), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n913), .B1(new_n982), .B2(new_n685), .ZN(new_n983));
  INV_X1    g797(.A(new_n981), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n984), .B1(new_n301), .B2(new_n275), .ZN(new_n985));
  AOI21_X1  g799(.A(KEYINPUT127), .B1(new_n859), .B2(new_n985), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n859), .A2(KEYINPUT127), .A3(new_n985), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n983), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n981), .B1(new_n951), .B2(new_n967), .ZN(new_n989));
  OR2_X1    g803(.A1(new_n989), .A2(KEYINPUT126), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(KEYINPUT126), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n300), .A2(new_n274), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n988), .B1(new_n992), .B2(new_n993), .ZN(G57));
endmodule


