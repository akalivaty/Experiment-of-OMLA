//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 0 0 1 0 1 1 1 0 0 0 0 1 1 1 1 1 0 1 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n631, new_n634, new_n636, new_n637, new_n638, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1211, new_n1212, new_n1213, new_n1214;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  OR4_X1    g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  XNOR2_X1  g033(.A(KEYINPUT3), .B(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G137), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(new_n462));
  AND2_X1   g037(.A1(new_n460), .A2(G2104), .ZN(new_n463));
  AOI22_X1  g038(.A1(new_n459), .A2(new_n462), .B1(new_n463), .B2(G101), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(G125), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n460), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n465), .A2(new_n470), .ZN(G160));
  NOR2_X1   g046(.A1(new_n466), .A2(new_n467), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(new_n460), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G124), .ZN(new_n474));
  OR2_X1    g049(.A1(G100), .A2(G2105), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n475), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n459), .A2(new_n460), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n477), .B1(G136), .B2(new_n479), .ZN(G162));
  INV_X1    g055(.A(KEYINPUT4), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n460), .A2(KEYINPUT66), .A3(G138), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n481), .B1(new_n472), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n459), .A2(G126), .A3(G2105), .ZN(new_n484));
  AND3_X1   g059(.A1(new_n460), .A2(KEYINPUT66), .A3(G138), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n459), .A2(KEYINPUT4), .A3(new_n485), .ZN(new_n486));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G114), .C2(new_n460), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n483), .A2(new_n484), .A3(new_n486), .A4(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G164));
  INV_X1    g065(.A(G62), .ZN(new_n491));
  OR2_X1    g066(.A1(KEYINPUT5), .A2(G543), .ZN(new_n492));
  NAND2_X1  g067(.A1(KEYINPUT5), .A2(G543), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AND2_X1   g069(.A1(G75), .A2(G543), .ZN(new_n495));
  OAI21_X1  g070(.A(G651), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT67), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT6), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(G651), .ZN(new_n499));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(KEYINPUT67), .A3(KEYINPUT6), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n503), .B1(new_n498), .B2(G651), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n502), .A2(G50), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G88), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n498), .A2(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n492), .A2(new_n493), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n502), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  OAI211_X1 g084(.A(new_n496), .B(new_n505), .C1(new_n506), .C2(new_n509), .ZN(G303));
  INV_X1    g085(.A(G303), .ZN(G166));
  OR2_X1    g086(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(KEYINPUT69), .A3(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT69), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  AND3_X1   g094(.A1(new_n514), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n519), .B1(new_n514), .B2(new_n518), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n502), .A2(G89), .A3(new_n508), .A4(new_n507), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n502), .A2(G51), .A3(new_n504), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n522), .A2(new_n526), .ZN(G168));
  AOI22_X1  g102(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(new_n500), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n502), .A2(new_n504), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT70), .B(G52), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AND3_X1   g108(.A1(new_n500), .A2(KEYINPUT67), .A3(KEYINPUT6), .ZN(new_n534));
  AOI21_X1  g109(.A(KEYINPUT67), .B1(new_n500), .B2(KEYINPUT6), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AND2_X1   g111(.A1(KEYINPUT5), .A2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(KEYINPUT5), .A2(G543), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n507), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G90), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n529), .A2(new_n533), .A3(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n537), .A2(new_n538), .ZN(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n500), .B1(new_n547), .B2(KEYINPUT71), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n548), .B1(KEYINPUT71), .B2(new_n547), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n540), .A2(G81), .B1(new_n531), .B2(G43), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  INV_X1    g132(.A(KEYINPUT76), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(KEYINPUT74), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G65), .ZN(new_n562));
  OAI211_X1 g137(.A(new_n560), .B(new_n562), .C1(new_n537), .C2(new_n538), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n563), .A2(KEYINPUT75), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G651), .ZN(new_n566));
  AOI21_X1  g141(.A(KEYINPUT75), .B1(new_n563), .B2(new_n564), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n558), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n563), .A2(new_n564), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n571), .A2(KEYINPUT76), .A3(G651), .A4(new_n565), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g148(.A(KEYINPUT73), .B1(new_n536), .B2(new_n539), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT73), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n502), .A2(new_n575), .A3(new_n508), .A4(new_n507), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(G91), .A3(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(G53), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n578), .A2(KEYINPUT72), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n504), .B(new_n579), .C1(new_n534), .C2(new_n535), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(KEYINPUT9), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT9), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n502), .A2(new_n582), .A3(new_n504), .A4(new_n579), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n577), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n573), .A2(new_n585), .ZN(G299));
  INV_X1    g161(.A(G168), .ZN(G286));
  NAND3_X1  g162(.A1(new_n574), .A2(G87), .A3(new_n576), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n502), .A2(G49), .A3(new_n504), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT77), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n502), .A2(KEYINPUT77), .A3(G49), .A4(new_n504), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(KEYINPUT78), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT78), .ZN(new_n596));
  OAI211_X1 g171(.A(new_n596), .B(G651), .C1(new_n508), .C2(G74), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n588), .A2(new_n593), .A3(new_n598), .ZN(G288));
  NAND2_X1  g174(.A1(G73), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G61), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n545), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n531), .A2(G48), .B1(new_n602), .B2(G651), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n574), .A2(G86), .A3(new_n576), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(G305));
  NAND2_X1  g180(.A1(new_n540), .A2(G85), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n531), .A2(G47), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n606), .B(new_n607), .C1(new_n500), .C2(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n574), .A2(G92), .A3(new_n576), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g188(.A1(new_n574), .A2(KEYINPUT10), .A3(G92), .A4(new_n576), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(G79), .A2(G543), .ZN(new_n616));
  INV_X1    g191(.A(G66), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n545), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G651), .ZN(new_n619));
  INV_X1    g194(.A(G54), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(new_n530), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g197(.A(KEYINPUT79), .B1(new_n615), .B2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT79), .ZN(new_n624));
  AOI211_X1 g199(.A(new_n624), .B(new_n621), .C1(new_n613), .C2(new_n614), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n610), .B1(new_n627), .B2(G868), .ZN(G284));
  OAI21_X1  g203(.A(new_n610), .B1(new_n627), .B2(G868), .ZN(G321));
  INV_X1    g204(.A(G868), .ZN(new_n630));
  NAND2_X1  g205(.A1(G299), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n630), .B2(G168), .ZN(G297));
  OAI21_X1  g207(.A(new_n631), .B1(new_n630), .B2(G168), .ZN(G280));
  INV_X1    g208(.A(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n627), .B1(new_n634), .B2(G860), .ZN(G148));
  OAI21_X1  g210(.A(KEYINPUT80), .B1(new_n552), .B2(G868), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n627), .A2(new_n634), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G868), .ZN(new_n638));
  MUX2_X1   g213(.A(KEYINPUT80), .B(new_n636), .S(new_n638), .Z(G323));
  XNOR2_X1  g214(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g215(.A1(new_n459), .A2(new_n463), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT13), .ZN(new_n643));
  INV_X1    g218(.A(G2100), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n473), .A2(G123), .ZN(new_n647));
  OR3_X1    g222(.A1(new_n460), .A2(KEYINPUT81), .A3(G111), .ZN(new_n648));
  OAI21_X1  g223(.A(KEYINPUT81), .B1(new_n460), .B2(G111), .ZN(new_n649));
  OR2_X1    g224(.A1(G99), .A2(G2105), .ZN(new_n650));
  NAND4_X1  g225(.A1(new_n648), .A2(G2104), .A3(new_n649), .A4(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(G135), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n647), .B(new_n651), .C1(new_n652), .C2(new_n478), .ZN(new_n653));
  INV_X1    g228(.A(G2096), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n645), .A2(new_n646), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT82), .Z(G156));
  INV_X1    g232(.A(KEYINPUT14), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2427), .B(G2438), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2430), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT15), .B(G2435), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n662), .B1(new_n661), .B2(new_n660), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2451), .B(G2454), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT16), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1341), .B(G1348), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n663), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2443), .B(G2446), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(G14), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n668), .A2(new_n669), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(G401));
  XOR2_X1   g248(.A(G2072), .B(G2078), .Z(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT17), .Z(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2067), .B(G2678), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT83), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2084), .B(G2090), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(new_n678), .B2(new_n674), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n679), .B1(KEYINPUT86), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(KEYINPUT86), .B2(new_n682), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n676), .A2(new_n678), .A3(new_n681), .ZN(new_n685));
  NOR3_X1   g260(.A1(new_n678), .A2(new_n674), .A3(new_n680), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT85), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT84), .B(KEYINPUT18), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  OAI211_X1 g265(.A(new_n684), .B(new_n685), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(new_n654), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT87), .B(G2100), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n691), .B(G2096), .ZN(new_n695));
  INV_X1    g270(.A(new_n693), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n694), .A2(new_n697), .ZN(G227));
  XNOR2_X1  g273(.A(G1971), .B(G1976), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT19), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(G1956), .B(G2474), .Z(new_n702));
  XOR2_X1   g277(.A(G1961), .B(G1966), .Z(new_n703));
  AND2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT20), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n702), .A2(new_n703), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  MUX2_X1   g284(.A(new_n709), .B(new_n708), .S(new_n701), .Z(new_n710));
  NOR2_X1   g285(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(G1981), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G1986), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT88), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n712), .A2(G1986), .ZN(new_n717));
  INV_X1    g292(.A(new_n715), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n712), .A2(G1986), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(G1991), .B(G1996), .ZN(new_n721));
  AND3_X1   g296(.A1(new_n716), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n721), .B1(new_n716), .B2(new_n720), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(G229));
  MUX2_X1   g299(.A(G6), .B(G305), .S(G16), .Z(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT32), .B(G1981), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  MUX2_X1   g302(.A(G23), .B(G288), .S(G16), .Z(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT33), .B(G1976), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT90), .B(G16), .Z(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n732), .A2(G22), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G166), .B2(new_n732), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(G1971), .Z(new_n735));
  NAND2_X1  g310(.A1(new_n725), .A2(new_n726), .ZN(new_n736));
  AND4_X1   g311(.A1(new_n727), .A2(new_n730), .A3(new_n735), .A4(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT34), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n479), .A2(G131), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n473), .A2(G119), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n460), .A2(G107), .ZN(new_n743));
  OAI21_X1  g318(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n741), .B(new_n742), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT89), .Z(new_n746));
  MUX2_X1   g321(.A(G25), .B(new_n746), .S(G29), .Z(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT35), .B(G1991), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  MUX2_X1   g324(.A(G24), .B(G290), .S(new_n732), .Z(new_n750));
  XOR2_X1   g325(.A(KEYINPUT91), .B(G1986), .Z(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n739), .A2(new_n740), .A3(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT36), .ZN(new_n755));
  AND3_X1   g330(.A1(new_n754), .A2(KEYINPUT92), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n754), .B1(KEYINPUT92), .B2(new_n755), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n755), .A2(KEYINPUT92), .ZN(new_n759));
  NOR2_X1   g334(.A1(G29), .A2(G35), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G162), .B2(G29), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT29), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(G2090), .Z(new_n763));
  NAND2_X1  g338(.A1(new_n731), .A2(G20), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT101), .Z(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT23), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G16), .B2(G299), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1956), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n763), .A2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(G29), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n770), .A2(G33), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT25), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(G139), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(new_n478), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT97), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n459), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n777), .B1(new_n460), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n771), .B1(new_n779), .B2(G29), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT98), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n780), .A2(new_n781), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n442), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n784), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n786), .A2(G2072), .A3(new_n782), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n770), .A2(G32), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n479), .A2(G141), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT99), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n463), .A2(G105), .ZN(new_n792));
  NAND3_X1  g367(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT26), .ZN(new_n794));
  AOI211_X1 g369(.A(new_n792), .B(new_n794), .C1(G129), .C2(new_n473), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n791), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n789), .B1(new_n796), .B2(new_n770), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT27), .B(G1996), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(G5), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n801), .A2(G16), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G301), .B2(G16), .ZN(new_n803));
  INV_X1    g378(.A(G1961), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n789), .B(new_n798), .C1(new_n796), .C2(new_n770), .ZN(new_n806));
  AND3_X1   g381(.A1(new_n800), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n770), .A2(G27), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G164), .B2(new_n770), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G2078), .ZN(new_n810));
  INV_X1    g385(.A(G2084), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n770), .B1(KEYINPUT24), .B2(G34), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(KEYINPUT24), .B2(G34), .ZN(new_n813));
  INV_X1    g388(.A(G160), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(G29), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n810), .B1(new_n811), .B2(new_n815), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT31), .B(G11), .Z(new_n817));
  INV_X1    g392(.A(G28), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n818), .A2(KEYINPUT30), .ZN(new_n819));
  AOI21_X1  g394(.A(G29), .B1(new_n818), .B2(KEYINPUT30), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n817), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI221_X1 g396(.A(new_n821), .B1(new_n770), .B2(new_n653), .C1(new_n815), .C2(new_n811), .ZN(new_n822));
  INV_X1    g397(.A(new_n803), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n822), .B1(G1961), .B2(new_n823), .ZN(new_n824));
  MUX2_X1   g399(.A(G21), .B(G286), .S(G16), .Z(new_n825));
  INV_X1    g400(.A(G1966), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n807), .A2(new_n816), .A3(new_n824), .A4(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n788), .A2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT100), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n769), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(KEYINPUT100), .B1(new_n788), .B2(new_n828), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n627), .A2(G16), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(G4), .B2(G16), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT93), .B(G1348), .Z(new_n836));
  OR2_X1    g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n836), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n479), .A2(G140), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n473), .A2(G128), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n460), .A2(G116), .ZN(new_n841));
  OAI21_X1  g416(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n839), .B(new_n840), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(G29), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n770), .A2(G26), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT28), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT95), .ZN(new_n848));
  INV_X1    g423(.A(G2067), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n731), .A2(G19), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT94), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n552), .B2(new_n731), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(G1341), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n837), .A2(new_n838), .A3(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT96), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n837), .A2(KEYINPUT96), .A3(new_n838), .A4(new_n855), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n833), .A2(KEYINPUT102), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT102), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n831), .A2(new_n859), .A3(new_n832), .ZN(new_n862));
  INV_X1    g437(.A(new_n858), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI22_X1  g439(.A1(new_n758), .A2(new_n759), .B1(new_n860), .B2(new_n864), .ZN(G311));
  NAND2_X1  g440(.A1(new_n860), .A2(new_n864), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n759), .B1(new_n756), .B2(new_n757), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(G150));
  NOR2_X1   g443(.A1(new_n626), .A2(new_n634), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT38), .ZN(new_n870));
  AOI22_X1  g445(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n871), .A2(new_n500), .ZN(new_n872));
  INV_X1    g447(.A(G93), .ZN(new_n873));
  INV_X1    g448(.A(G55), .ZN(new_n874));
  OAI22_X1  g449(.A1(new_n509), .A2(new_n873), .B1(new_n530), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT103), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n875), .A2(new_n876), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n872), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(new_n551), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n875), .B(new_n876), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n552), .A2(new_n881), .A3(new_n872), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n870), .B(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT39), .ZN(new_n886));
  AOI21_X1  g461(.A(G860), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n887), .B1(new_n886), .B2(new_n885), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n879), .A2(G860), .ZN(new_n889));
  XOR2_X1   g464(.A(new_n889), .B(KEYINPUT37), .Z(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(G145));
  XNOR2_X1  g466(.A(new_n843), .B(G164), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n779), .B(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n796), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n893), .B(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n479), .A2(G142), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n473), .A2(G130), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n460), .A2(G118), .ZN(new_n898));
  OAI21_X1  g473(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n896), .B(new_n897), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(new_n642), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n745), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT104), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n895), .B(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n653), .B(G160), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(G162), .ZN(new_n906));
  AOI21_X1  g481(.A(G37), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n906), .B1(new_n895), .B2(new_n903), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n895), .A2(KEYINPUT105), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n902), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n895), .A2(KEYINPUT105), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n907), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g489(.A1(new_n637), .A2(new_n884), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n627), .A2(new_n883), .A3(new_n634), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n615), .A2(new_n622), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n918), .A2(G299), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(G299), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT41), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n921), .B(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n917), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n915), .A2(new_n921), .A3(new_n916), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n926), .A2(KEYINPUT42), .ZN(new_n927));
  XOR2_X1   g502(.A(G290), .B(G305), .Z(new_n928));
  XNOR2_X1  g503(.A(G288), .B(G166), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n928), .B(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n926), .A2(KEYINPUT42), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n927), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n931), .B1(new_n927), .B2(new_n932), .ZN(new_n934));
  OAI21_X1  g509(.A(G868), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n879), .A2(new_n630), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(G295));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n936), .ZN(G331));
  INV_X1    g513(.A(KEYINPUT106), .ZN(new_n939));
  OAI21_X1  g514(.A(G301), .B1(G168), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(G168), .A2(new_n939), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n880), .A2(new_n882), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n941), .B1(new_n880), .B2(new_n882), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n941), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n883), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n940), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n880), .A2(new_n882), .A3(new_n941), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n944), .A2(new_n949), .A3(new_n920), .A4(new_n919), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n944), .A2(new_n949), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n950), .B1(new_n951), .B2(new_n923), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n931), .ZN(new_n953));
  INV_X1    g528(.A(G37), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n930), .B(new_n950), .C1(new_n951), .C2(new_n923), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n953), .A2(new_n958), .A3(new_n954), .A4(new_n955), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n957), .A2(KEYINPUT107), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n956), .A2(new_n962), .A3(KEYINPUT43), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n960), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n957), .A2(KEYINPUT44), .A3(new_n959), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(G397));
  INV_X1    g541(.A(G1384), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n489), .A2(new_n967), .ZN(new_n968));
  OR2_X1    g543(.A1(new_n968), .A2(KEYINPUT108), .ZN(new_n969));
  INV_X1    g544(.A(G125), .ZN(new_n970));
  OR2_X1    g545(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n971));
  NAND2_X1  g546(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n469), .ZN(new_n974));
  OAI21_X1  g549(.A(G2105), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n975), .A2(new_n976), .A3(G40), .A4(new_n464), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n460), .A2(G101), .A3(G2104), .ZN(new_n978));
  OAI211_X1 g553(.A(G40), .B(new_n978), .C1(new_n472), .C2(new_n461), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT109), .B1(new_n470), .B2(new_n979), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT45), .B1(new_n968), .B2(KEYINPUT108), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n969), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n984));
  OR2_X1    g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n984), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n894), .A2(G1996), .ZN(new_n989));
  OR3_X1    g564(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n988), .B1(new_n987), .B2(new_n989), .ZN(new_n991));
  INV_X1    g566(.A(new_n987), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n843), .B(new_n849), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n993), .B1(new_n894), .B2(G1996), .ZN(new_n994));
  AOI22_X1  g569(.A1(new_n990), .A2(new_n991), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n745), .B(KEYINPUT112), .ZN(new_n996));
  XOR2_X1   g571(.A(new_n996), .B(new_n748), .Z(new_n997));
  OAI21_X1  g572(.A(new_n995), .B1(new_n987), .B2(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(G290), .B(G1986), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n998), .B1(new_n992), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n968), .A2(KEYINPUT50), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT50), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n489), .A2(new_n1002), .A3(new_n967), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n981), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1956), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT57), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n573), .A2(new_n585), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n977), .A2(new_n980), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT45), .B1(new_n489), .B2(new_n967), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n489), .A2(KEYINPUT45), .A3(new_n967), .ZN(new_n1013));
  XNOR2_X1  g588(.A(KEYINPUT56), .B(G2072), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1006), .A2(new_n1007), .A3(new_n1009), .A4(new_n1015), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n981), .A2(new_n967), .A3(new_n849), .A4(new_n489), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1003), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1002), .B1(new_n489), .B2(new_n967), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n1018), .A2(new_n1010), .A3(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1017), .B1(new_n1020), .B2(G1348), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1016), .A2(new_n627), .A3(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1010), .A2(new_n1019), .ZN(new_n1023));
  AOI21_X1  g598(.A(G1956), .B1(new_n1023), .B2(new_n1003), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT45), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n968), .A2(new_n1025), .ZN(new_n1026));
  AND4_X1   g601(.A1(new_n981), .A2(new_n1026), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n573), .A2(new_n585), .A3(new_n1008), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1008), .B1(new_n573), .B2(new_n585), .ZN(new_n1029));
  OAI22_X1  g604(.A1(new_n1024), .A2(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n1022), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT61), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1030), .A2(new_n1016), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1032), .B1(new_n1030), .B2(new_n1016), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1348), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1010), .A2(new_n968), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n1004), .A2(new_n1036), .B1(new_n1037), .B2(new_n849), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1038), .B(KEYINPUT60), .C1(new_n623), .C2(new_n625), .ZN(new_n1039));
  OAI211_X1 g614(.A(KEYINPUT60), .B(new_n1017), .C1(new_n1020), .C2(G1348), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n626), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT60), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1021), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1039), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT119), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT59), .ZN(new_n1046));
  INV_X1    g621(.A(G1996), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n981), .A2(new_n1026), .A3(new_n1047), .A4(new_n1013), .ZN(new_n1048));
  XOR2_X1   g623(.A(KEYINPUT58), .B(G1341), .Z(new_n1049));
  OAI21_X1  g624(.A(new_n1049), .B1(new_n1010), .B2(new_n968), .ZN(new_n1050));
  AOI211_X1 g625(.A(new_n551), .B(new_n1046), .C1(new_n1048), .C2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n552), .ZN(new_n1053));
  XNOR2_X1  g628(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1051), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1044), .A2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1031), .B1(new_n1035), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT120), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT120), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1059), .B(new_n1031), .C1(new_n1035), .C2(new_n1056), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n1061));
  NOR4_X1   g636(.A1(new_n470), .A2(new_n979), .A3(new_n1061), .A4(G2078), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n1013), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1063), .B1(new_n969), .B2(new_n982), .ZN(new_n1064));
  XNOR2_X1  g639(.A(G301), .B(KEYINPUT54), .ZN(new_n1065));
  AOI211_X1 g640(.A(new_n1064), .B(new_n1065), .C1(new_n804), .C2(new_n1004), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n981), .A2(new_n1026), .A3(new_n1013), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1061), .B1(new_n1067), .B2(G2078), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1013), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n1069), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1070), .A2(KEYINPUT53), .A3(new_n443), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1071), .B(new_n1068), .C1(G1961), .C2(new_n1020), .ZN(new_n1072));
  AOI22_X1  g647(.A1(new_n1066), .A2(new_n1068), .B1(new_n1072), .B2(new_n1065), .ZN(new_n1073));
  OAI21_X1  g648(.A(G8), .B1(new_n522), .B2(new_n526), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT121), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT123), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT121), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1077), .B(G8), .C1(new_n522), .C2(new_n526), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1075), .A2(new_n1076), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT51), .ZN(new_n1080));
  INV_X1    g655(.A(G8), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1067), .A2(new_n826), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1023), .A2(new_n811), .A3(new_n1003), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1081), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1080), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(G1966), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1087));
  AND4_X1   g662(.A1(new_n811), .A2(new_n981), .A3(new_n1001), .A4(new_n1003), .ZN(new_n1088));
  OAI21_X1  g663(.A(G8), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1085), .ZN(new_n1090));
  AND2_X1   g665(.A1(new_n1079), .A2(KEYINPUT51), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1086), .A2(new_n1092), .ZN(new_n1093));
  AOI221_X4 g668(.A(KEYINPUT122), .B1(new_n1078), .B2(new_n1075), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n1095));
  OAI22_X1  g670(.A1(new_n1070), .A2(G1966), .B1(new_n1004), .B2(G2084), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1095), .B1(new_n1096), .B2(new_n1085), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1073), .B1(new_n1093), .B2(new_n1098), .ZN(new_n1099));
  OAI22_X1  g674(.A1(new_n1070), .A2(G1971), .B1(new_n1004), .B2(G2090), .ZN(new_n1100));
  NAND2_X1  g675(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(G303), .A2(G8), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1101), .B1(G303), .B2(G8), .ZN(new_n1107));
  OAI21_X1  g682(.A(KEYINPUT114), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(G303), .A2(G8), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(new_n1102), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT114), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1110), .A2(new_n1111), .A3(new_n1105), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1108), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1100), .A2(new_n1113), .A3(G8), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT115), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1100), .A2(new_n1113), .A3(new_n1116), .A4(G8), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(G1976), .ZN(new_n1119));
  NAND2_X1  g694(.A1(G288), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT52), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT117), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n588), .A2(new_n593), .A3(new_n598), .A4(G1976), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1124), .A2(KEYINPUT116), .ZN(new_n1125));
  OAI21_X1  g700(.A(G8), .B1(new_n1010), .B2(new_n968), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1124), .A2(KEYINPUT116), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT117), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1120), .A2(new_n1129), .A3(new_n1121), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1123), .A2(new_n1127), .A3(new_n1128), .A4(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n540), .A2(G86), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n603), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(G1981), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(G305), .B2(G1981), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT49), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1126), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1134), .B(KEYINPUT49), .C1(G1981), .C2(G305), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  OAI221_X1 g715(.A(G8), .B1(new_n1010), .B2(new_n968), .C1(new_n1124), .C2(KEYINPUT116), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1128), .ZN(new_n1142));
  OAI21_X1  g717(.A(KEYINPUT52), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1131), .A2(new_n1140), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1100), .A2(G8), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1110), .A2(new_n1105), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1118), .A2(new_n1145), .A3(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1099), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1058), .A2(new_n1060), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT124), .ZN(new_n1152));
  NOR2_X1   g727(.A1(G288), .A2(G1976), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1140), .A2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(G305), .A2(G1981), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1138), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1156), .B1(new_n1118), .B2(new_n1144), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1089), .A2(G286), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1118), .A2(new_n1145), .A3(new_n1148), .A4(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT63), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT118), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1145), .A2(new_n1162), .A3(new_n1148), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1148), .ZN(new_n1164));
  OAI21_X1  g739(.A(KEYINPUT118), .B1(new_n1164), .B2(new_n1144), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1084), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1166), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1163), .A2(new_n1165), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1157), .B1(new_n1161), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1151), .A2(new_n1152), .A3(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(KEYINPUT62), .B1(new_n1093), .B2(new_n1098), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1096), .A2(new_n1085), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(KEYINPUT122), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1096), .A2(new_n1095), .A3(new_n1085), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT62), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1175), .A2(new_n1176), .A3(new_n1092), .A4(new_n1086), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1171), .A2(new_n1177), .ZN(new_n1178));
  AND2_X1   g753(.A1(new_n1072), .A2(G171), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1118), .A2(new_n1145), .A3(new_n1148), .A4(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(KEYINPUT125), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1180), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT125), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1182), .A2(new_n1183), .A3(new_n1171), .A4(new_n1177), .ZN(new_n1184));
  AND2_X1   g759(.A1(new_n1181), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1170), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1152), .B1(new_n1151), .B2(new_n1169), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1000), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n843), .A2(G2067), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n746), .A2(new_n748), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1189), .B1(new_n995), .B2(new_n1190), .ZN(new_n1191));
  NOR3_X1   g766(.A1(new_n987), .A2(G1986), .A3(G290), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n1192), .B(KEYINPUT48), .ZN(new_n1193));
  OAI22_X1  g768(.A1(new_n1191), .A2(new_n987), .B1(new_n998), .B2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n992), .A2(KEYINPUT46), .A3(new_n1047), .ZN(new_n1195));
  XNOR2_X1  g770(.A(new_n1195), .B(KEYINPUT126), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT127), .ZN(new_n1197));
  AOI21_X1  g772(.A(KEYINPUT46), .B1(new_n992), .B2(new_n1047), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n987), .B1(new_n796), .B2(new_n993), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1196), .A2(new_n1197), .A3(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(new_n1201), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1197), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1203));
  OAI21_X1  g778(.A(KEYINPUT47), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g779(.A(new_n1203), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT47), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1205), .A2(new_n1206), .A3(new_n1201), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1194), .B1(new_n1204), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1188), .A2(new_n1208), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g784(.A(G319), .B1(new_n671), .B2(new_n672), .ZN(new_n1211));
  AOI21_X1  g785(.A(new_n1211), .B1(new_n694), .B2(new_n697), .ZN(new_n1212));
  OAI21_X1  g786(.A(new_n1212), .B1(new_n722), .B2(new_n723), .ZN(new_n1213));
  AOI21_X1  g787(.A(new_n1213), .B1(new_n912), .B2(new_n907), .ZN(new_n1214));
  NAND3_X1  g788(.A1(new_n1214), .A2(new_n963), .A3(new_n960), .ZN(G225));
  INV_X1    g789(.A(G225), .ZN(G308));
endmodule


