

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791;

  NOR2_X1 U376 ( .A1(n422), .A2(n374), .ZN(n373) );
  NAND2_X1 U377 ( .A1(n369), .A2(n383), .ZN(n634) );
  AND2_X1 U378 ( .A1(n597), .A2(n594), .ZN(n612) );
  XNOR2_X1 U379 ( .A(n388), .B(n574), .ZN(n606) );
  OR2_X1 U380 ( .A1(n681), .A2(G902), .ZN(n497) );
  XNOR2_X1 U381 ( .A(G116), .B(G122), .ZN(n541) );
  XNOR2_X1 U382 ( .A(G146), .B(G125), .ZN(n358) );
  XNOR2_X1 U383 ( .A(KEYINPUT78), .B(G122), .ZN(n438) );
  INV_X1 U384 ( .A(G134), .ZN(n538) );
  XNOR2_X2 U385 ( .A(n726), .B(n549), .ZN(n610) );
  XNOR2_X1 U386 ( .A(n356), .B(KEYINPUT84), .ZN(n386) );
  NAND2_X1 U387 ( .A1(n663), .A2(n357), .ZN(n356) );
  NAND2_X1 U388 ( .A1(n371), .A2(n370), .ZN(n357) );
  XNOR2_X2 U389 ( .A(n782), .B(n403), .ZN(n689) );
  XNOR2_X2 U390 ( .A(n394), .B(KEYINPUT39), .ZN(n583) );
  XNOR2_X2 U391 ( .A(KEYINPUT81), .B(KEYINPUT34), .ZN(n570) );
  XNOR2_X2 U392 ( .A(n381), .B(KEYINPUT33), .ZN(n569) );
  XNOR2_X2 U393 ( .A(n456), .B(G902), .ZN(n664) );
  INV_X2 U394 ( .A(KEYINPUT71), .ZN(n399) );
  BUF_X1 U395 ( .A(G113), .Z(n396) );
  AND2_X2 U396 ( .A1(n603), .A2(n604), .ZN(n401) );
  XNOR2_X2 U397 ( .A(G143), .B(G128), .ZN(n540) );
  XNOR2_X2 U398 ( .A(n520), .B(n471), .ZN(n782) );
  XNOR2_X2 U399 ( .A(n406), .B(n455), .ZN(n520) );
  XNOR2_X2 U400 ( .A(n439), .B(G107), .ZN(n502) );
  XNOR2_X2 U401 ( .A(G104), .B(G110), .ZN(n439) );
  NOR2_X1 U402 ( .A1(n553), .A2(n723), .ZN(n554) );
  INV_X1 U403 ( .A(KEYINPUT77), .ZN(n441) );
  NAND2_X1 U404 ( .A1(n421), .A2(KEYINPUT88), .ZN(n420) );
  NAND2_X1 U405 ( .A1(n447), .A2(KEYINPUT44), .ZN(n446) );
  NAND2_X1 U406 ( .A1(n591), .A2(n363), .ZN(n641) );
  XNOR2_X1 U407 ( .A(n675), .B(n676), .ZN(n677) );
  AND2_X1 U408 ( .A1(n419), .A2(n418), .ZN(n417) );
  XNOR2_X1 U409 ( .A(n440), .B(n489), .ZN(n503) );
  XNOR2_X1 U410 ( .A(n442), .B(n441), .ZN(n440) );
  XNOR2_X1 U411 ( .A(KEYINPUT72), .B(G137), .ZN(n471) );
  XNOR2_X2 U412 ( .A(G146), .B(G125), .ZN(n505) );
  BUF_X1 U413 ( .A(n599), .Z(n359) );
  XNOR2_X1 U414 ( .A(n658), .B(n657), .ZN(n428) );
  NAND2_X1 U415 ( .A1(n417), .A2(n413), .ZN(n631) );
  XNOR2_X2 U416 ( .A(n533), .B(n532), .ZN(n577) );
  BUF_X1 U417 ( .A(n408), .Z(n360) );
  BUF_X1 U418 ( .A(n638), .Z(n361) );
  XNOR2_X1 U419 ( .A(n503), .B(n435), .ZN(n408) );
  NAND2_X1 U420 ( .A1(n728), .A2(n380), .ZN(n617) );
  NAND2_X1 U421 ( .A1(n583), .A2(n764), .ZN(n584) );
  AND2_X1 U422 ( .A1(n363), .A2(n728), .ZN(n362) );
  XNOR2_X1 U423 ( .A(n380), .B(KEYINPUT1), .ZN(n363) );
  AND2_X2 U424 ( .A1(n593), .A2(n552), .ZN(n728) );
  XNOR2_X1 U425 ( .A(n631), .B(KEYINPUT1), .ZN(n561) );
  BUF_X1 U426 ( .A(n688), .Z(n696) );
  NAND2_X1 U427 ( .A1(n561), .A2(n728), .ZN(n614) );
  NAND2_X1 U428 ( .A1(n365), .A2(n422), .ZN(n370) );
  XNOR2_X1 U429 ( .A(n400), .B(KEYINPUT74), .ZN(n629) );
  INV_X1 U430 ( .A(KEYINPUT79), .ZN(n374) );
  AND2_X1 U431 ( .A1(n407), .A2(n623), .ZN(n624) );
  XNOR2_X1 U432 ( .A(n476), .B(n475), .ZN(n477) );
  AND2_X1 U433 ( .A1(n448), .A2(n607), .ZN(n609) );
  NAND2_X1 U434 ( .A1(n434), .A2(n433), .ZN(n535) );
  NAND2_X1 U435 ( .A1(n431), .A2(G234), .ZN(n433) );
  NAND2_X1 U436 ( .A1(n432), .A2(KEYINPUT8), .ZN(n434) );
  NOR2_X1 U437 ( .A1(KEYINPUT8), .A2(G953), .ZN(n431) );
  XOR2_X1 U438 ( .A(KEYINPUT70), .B(KEYINPUT10), .Z(n455) );
  INV_X1 U439 ( .A(G140), .ZN(n454) );
  AND2_X1 U440 ( .A1(n425), .A2(n661), .ZN(n424) );
  NAND2_X1 U441 ( .A1(n426), .A2(KEYINPUT88), .ZN(n425) );
  XNOR2_X1 U442 ( .A(n617), .B(n410), .ZN(n409) );
  INV_X1 U443 ( .A(KEYINPUT110), .ZN(n410) );
  XNOR2_X1 U444 ( .A(G128), .B(G119), .ZN(n452) );
  XNOR2_X1 U445 ( .A(n408), .B(n512), .ZN(n674) );
  INV_X2 U446 ( .A(G953), .ZN(n775) );
  XNOR2_X1 U447 ( .A(n459), .B(KEYINPUT25), .ZN(n460) );
  NOR2_X1 U448 ( .A1(n775), .A2(G952), .ZN(n703) );
  NOR2_X1 U449 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U450 ( .A1(n775), .A2(G234), .ZN(n432) );
  NOR2_X1 U451 ( .A1(n373), .A2(n372), .ZN(n371) );
  NOR2_X1 U452 ( .A1(n420), .A2(n374), .ZN(n372) );
  INV_X1 U453 ( .A(n659), .ZN(n426) );
  INV_X1 U454 ( .A(G237), .ZN(n498) );
  NAND2_X1 U455 ( .A1(n416), .A2(n415), .ZN(n414) );
  NOR2_X1 U456 ( .A1(G953), .A2(G237), .ZN(n523) );
  XOR2_X1 U457 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n491) );
  INV_X1 U458 ( .A(G104), .ZN(n517) );
  XNOR2_X1 U459 ( .A(n396), .B(G122), .ZN(n521) );
  XNOR2_X1 U460 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n507) );
  INV_X1 U461 ( .A(KEYINPUT15), .ZN(n456) );
  NAND2_X1 U462 ( .A1(G234), .A2(G237), .ZN(n478) );
  NAND2_X1 U463 ( .A1(n382), .A2(n610), .ZN(n381) );
  XNOR2_X1 U464 ( .A(n614), .B(KEYINPUT107), .ZN(n382) );
  XNOR2_X1 U465 ( .A(n514), .B(n515), .ZN(n712) );
  XNOR2_X1 U466 ( .A(n548), .B(n547), .ZN(n576) );
  NOR2_X1 U467 ( .A1(G902), .A2(n692), .ZN(n548) );
  INV_X1 U468 ( .A(G478), .ZN(n546) );
  XOR2_X1 U469 ( .A(KEYINPUT7), .B(KEYINPUT101), .Z(n542) );
  NOR2_X1 U470 ( .A1(n761), .A2(n629), .ZN(n555) );
  NAND2_X1 U471 ( .A1(n389), .A2(n573), .ZN(n388) );
  XNOR2_X1 U472 ( .A(n488), .B(n487), .ZN(n501) );
  NAND2_X1 U473 ( .A1(n409), .A2(n486), .ZN(n488) );
  XNOR2_X1 U474 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U475 ( .A(n681), .B(KEYINPUT62), .ZN(n682) );
  INV_X1 U476 ( .A(n785), .ZN(n375) );
  XNOR2_X1 U477 ( .A(n502), .B(n436), .ZN(n435) );
  XNOR2_X1 U478 ( .A(n438), .B(n437), .ZN(n436) );
  INV_X1 U479 ( .A(KEYINPUT16), .ZN(n437) );
  XNOR2_X1 U480 ( .A(n405), .B(n404), .ZN(n403) );
  NAND2_X1 U481 ( .A1(n450), .A2(G221), .ZN(n404) );
  XNOR2_X1 U482 ( .A(n453), .B(n451), .ZN(n405) );
  NOR2_X1 U483 ( .A1(n639), .A2(n744), .ZN(n384) );
  INV_X1 U484 ( .A(n734), .ZN(n391) );
  INV_X1 U485 ( .A(n618), .ZN(n392) );
  INV_X1 U486 ( .A(n429), .ZN(n611) );
  INV_X1 U487 ( .A(n703), .ZN(n397) );
  AND2_X1 U488 ( .A1(n568), .A2(n392), .ZN(n364) );
  AND2_X1 U489 ( .A1(n420), .A2(n374), .ZN(n365) );
  NOR2_X1 U490 ( .A1(n715), .A2(n723), .ZN(n366) );
  INV_X1 U491 ( .A(G902), .ZN(n415) );
  XOR2_X1 U492 ( .A(n672), .B(n671), .Z(n367) );
  XNOR2_X1 U493 ( .A(KEYINPUT67), .B(KEYINPUT60), .ZN(n368) );
  XNOR2_X1 U494 ( .A(n369), .B(G131), .ZN(G33) );
  XNOR2_X2 U495 ( .A(n584), .B(KEYINPUT40), .ZN(n369) );
  AND2_X1 U496 ( .A1(n422), .A2(n420), .ZN(n705) );
  XNOR2_X1 U497 ( .A(n705), .B(n375), .ZN(n783) );
  XNOR2_X2 U498 ( .A(n376), .B(n460), .ZN(n593) );
  OR2_X2 U499 ( .A1(n689), .A2(G902), .ZN(n376) );
  XNOR2_X1 U500 ( .A(G143), .B(G128), .ZN(n377) );
  XNOR2_X2 U501 ( .A(n378), .B(n379), .ZN(n562) );
  NOR2_X2 U502 ( .A1(n674), .A2(n664), .ZN(n378) );
  NAND2_X1 U503 ( .A1(n513), .A2(G210), .ZN(n379) );
  INV_X1 U504 ( .A(n593), .ZN(n430) );
  NAND2_X1 U505 ( .A1(n417), .A2(n413), .ZN(n380) );
  NAND2_X1 U506 ( .A1(n688), .A2(G475), .ZN(n673) );
  XNOR2_X1 U507 ( .A(n390), .B(n570), .ZN(n389) );
  AND2_X2 U508 ( .A1(n385), .A2(n709), .ZN(n688) );
  XNOR2_X2 U509 ( .A(n497), .B(G472), .ZN(n726) );
  INV_X1 U510 ( .A(n790), .ZN(n383) );
  XNOR2_X1 U511 ( .A(n384), .B(KEYINPUT42), .ZN(n790) );
  NAND2_X1 U512 ( .A1(n554), .A2(n430), .ZN(n400) );
  NAND2_X1 U513 ( .A1(n386), .A2(n665), .ZN(n385) );
  NAND2_X1 U514 ( .A1(n569), .A2(n568), .ZN(n390) );
  NAND2_X1 U515 ( .A1(n568), .A2(n366), .ZN(n579) );
  NAND2_X1 U516 ( .A1(n568), .A2(n391), .ZN(n616) );
  XNOR2_X2 U517 ( .A(n402), .B(KEYINPUT0), .ZN(n568) );
  AND2_X1 U518 ( .A1(n501), .A2(n500), .ZN(n648) );
  NAND2_X1 U519 ( .A1(n501), .A2(n393), .ZN(n394) );
  AND2_X1 U520 ( .A1(n500), .A2(n712), .ZN(n393) );
  XNOR2_X1 U521 ( .A(n395), .B(n368), .ZN(G60) );
  NAND2_X1 U522 ( .A1(n398), .A2(n397), .ZN(n395) );
  XNOR2_X1 U523 ( .A(n673), .B(n367), .ZN(n398) );
  XNOR2_X2 U524 ( .A(n399), .B(G131), .ZN(n516) );
  XNOR2_X2 U525 ( .A(KEYINPUT109), .B(n556), .ZN(n587) );
  OR2_X2 U526 ( .A1(n577), .A2(n571), .ZN(n551) );
  XNOR2_X1 U527 ( .A(n518), .B(n517), .ZN(n519) );
  NAND2_X1 U528 ( .A1(n401), .A2(n624), .ZN(n443) );
  NOR2_X2 U529 ( .A1(n638), .A2(n567), .ZN(n402) );
  XNOR2_X2 U530 ( .A(n585), .B(KEYINPUT19), .ZN(n638) );
  XNOR2_X2 U531 ( .A(n563), .B(KEYINPUT91), .ZN(n585) );
  XNOR2_X1 U532 ( .A(n505), .B(n454), .ZN(n406) );
  XNOR2_X1 U533 ( .A(n407), .B(G101), .ZN(G3) );
  XNOR2_X2 U534 ( .A(n613), .B(KEYINPUT106), .ZN(n407) );
  XNOR2_X1 U535 ( .A(n360), .B(G101), .ZN(n771) );
  NAND2_X1 U536 ( .A1(n562), .A2(n711), .ZN(n563) );
  XNOR2_X2 U537 ( .A(KEYINPUT68), .B(G101), .ZN(n504) );
  NAND2_X1 U538 ( .A1(n667), .A2(n664), .ZN(n626) );
  XNOR2_X1 U539 ( .A(n411), .B(n625), .ZN(n667) );
  NAND2_X1 U540 ( .A1(n412), .A2(n446), .ZN(n411) );
  NAND2_X1 U541 ( .A1(n443), .A2(n444), .ZN(n412) );
  INV_X1 U542 ( .A(n569), .ZN(n720) );
  XNOR2_X2 U543 ( .A(n516), .B(n538), .ZN(n468) );
  OR2_X1 U544 ( .A1(n697), .A2(n414), .ZN(n413) );
  INV_X1 U545 ( .A(n477), .ZN(n416) );
  NAND2_X1 U546 ( .A1(n477), .A2(G902), .ZN(n418) );
  NAND2_X1 U547 ( .A1(n697), .A2(n477), .ZN(n419) );
  XNOR2_X2 U548 ( .A(n496), .B(n474), .ZN(n697) );
  XNOR2_X2 U549 ( .A(n540), .B(n467), .ZN(n510) );
  INV_X1 U550 ( .A(n428), .ZN(n421) );
  AND2_X2 U551 ( .A1(n423), .A2(n424), .ZN(n422) );
  NAND2_X1 U552 ( .A1(n428), .A2(n427), .ZN(n423) );
  AND2_X1 U553 ( .A1(n659), .A2(n660), .ZN(n427) );
  NAND2_X1 U554 ( .A1(n430), .A2(n723), .ZN(n724) );
  OR2_X1 U555 ( .A1(n610), .A2(n430), .ZN(n429) );
  NAND2_X1 U556 ( .A1(n582), .A2(n430), .ZN(n608) );
  XNOR2_X2 U557 ( .A(G116), .B(G113), .ZN(n442) );
  NAND2_X1 U558 ( .A1(n445), .A2(n624), .ZN(n444) );
  NAND2_X1 U559 ( .A1(n608), .A2(n607), .ZN(n445) );
  NAND2_X1 U560 ( .A1(n609), .A2(n608), .ZN(n447) );
  XNOR2_X1 U561 ( .A(KEYINPUT3), .B(G119), .ZN(n489) );
  XNOR2_X1 U562 ( .A(n520), .B(n519), .ZN(n529) );
  AND2_X1 U563 ( .A1(n606), .A2(n605), .ZN(n448) );
  XOR2_X1 U564 ( .A(n542), .B(n541), .Z(n449) );
  XNOR2_X1 U565 ( .A(n546), .B(KEYINPUT103), .ZN(n547) );
  XNOR2_X1 U566 ( .A(n543), .B(n449), .ZN(n544) );
  XNOR2_X1 U567 ( .A(n545), .B(n544), .ZN(n692) );
  BUF_X1 U568 ( .A(n697), .Z(n700) );
  INV_X1 U569 ( .A(n535), .ZN(n450) );
  XNOR2_X1 U570 ( .A(G110), .B(KEYINPUT24), .ZN(n451) );
  XNOR2_X1 U571 ( .A(n452), .B(KEYINPUT23), .ZN(n453) );
  INV_X1 U572 ( .A(n664), .ZN(n457) );
  NAND2_X1 U573 ( .A1(n457), .A2(G234), .ZN(n458) );
  XNOR2_X1 U574 ( .A(n458), .B(KEYINPUT20), .ZN(n461) );
  AND2_X1 U575 ( .A1(n461), .A2(G217), .ZN(n459) );
  INV_X1 U576 ( .A(n461), .ZN(n463) );
  INV_X1 U577 ( .A(G221), .ZN(n462) );
  OR2_X1 U578 ( .A1(n463), .A2(n462), .ZN(n466) );
  INV_X1 U579 ( .A(KEYINPUT94), .ZN(n464) );
  XNOR2_X1 U580 ( .A(n464), .B(KEYINPUT21), .ZN(n465) );
  XNOR2_X1 U581 ( .A(n466), .B(n465), .ZN(n552) );
  XNOR2_X2 U582 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n467) );
  XNOR2_X2 U583 ( .A(n468), .B(n510), .ZN(n781) );
  XNOR2_X1 U584 ( .A(n504), .B(G146), .ZN(n469) );
  XNOR2_X2 U585 ( .A(n781), .B(n469), .ZN(n496) );
  NAND2_X1 U586 ( .A1(n775), .A2(G227), .ZN(n470) );
  XNOR2_X1 U587 ( .A(n470), .B(G140), .ZN(n472) );
  XNOR2_X1 U588 ( .A(n472), .B(n471), .ZN(n473) );
  XOR2_X1 U589 ( .A(n502), .B(n473), .Z(n474) );
  XNOR2_X1 U590 ( .A(KEYINPUT76), .B(G469), .ZN(n476) );
  INV_X1 U591 ( .A(KEYINPUT75), .ZN(n475) );
  XOR2_X1 U592 ( .A(KEYINPUT14), .B(KEYINPUT93), .Z(n479) );
  XNOR2_X1 U593 ( .A(n479), .B(n478), .ZN(n482) );
  NAND2_X1 U594 ( .A1(G902), .A2(n482), .ZN(n564) );
  NOR2_X1 U595 ( .A1(G900), .A2(n564), .ZN(n480) );
  NAND2_X1 U596 ( .A1(G953), .A2(n480), .ZN(n481) );
  XOR2_X1 U597 ( .A(KEYINPUT108), .B(n481), .Z(n484) );
  NAND2_X1 U598 ( .A1(G952), .A2(n482), .ZN(n743) );
  OR2_X1 U599 ( .A1(n743), .A2(G953), .ZN(n566) );
  INV_X1 U600 ( .A(n566), .ZN(n483) );
  NOR2_X1 U601 ( .A1(n484), .A2(n483), .ZN(n485) );
  XNOR2_X1 U602 ( .A(n485), .B(KEYINPUT82), .ZN(n553) );
  INV_X1 U603 ( .A(n553), .ZN(n486) );
  INV_X1 U604 ( .A(KEYINPUT80), .ZN(n487) );
  XNOR2_X1 U605 ( .A(G137), .B(KEYINPUT5), .ZN(n490) );
  XNOR2_X1 U606 ( .A(n491), .B(n490), .ZN(n493) );
  NAND2_X1 U607 ( .A1(n523), .A2(G210), .ZN(n492) );
  XNOR2_X1 U608 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U609 ( .A(n503), .B(n494), .ZN(n495) );
  XNOR2_X1 U610 ( .A(n496), .B(n495), .ZN(n681) );
  NAND2_X1 U611 ( .A1(n415), .A2(n498), .ZN(n513) );
  NAND2_X1 U612 ( .A1(n513), .A2(G214), .ZN(n711) );
  AND2_X1 U613 ( .A1(n726), .A2(n711), .ZN(n499) );
  XNOR2_X1 U614 ( .A(n499), .B(KEYINPUT30), .ZN(n500) );
  XNOR2_X1 U615 ( .A(n358), .B(n504), .ZN(n509) );
  NAND2_X1 U616 ( .A1(n775), .A2(G224), .ZN(n506) );
  XNOR2_X1 U617 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U618 ( .A(n509), .B(n508), .ZN(n511) );
  XNOR2_X1 U619 ( .A(n510), .B(n511), .ZN(n512) );
  BUF_X1 U620 ( .A(n562), .Z(n514) );
  INV_X1 U621 ( .A(KEYINPUT38), .ZN(n515) );
  XNOR2_X1 U622 ( .A(n516), .B(G143), .ZN(n518) );
  XOR2_X1 U623 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n522) );
  XNOR2_X1 U624 ( .A(n522), .B(n521), .ZN(n527) );
  XOR2_X1 U625 ( .A(KEYINPUT11), .B(KEYINPUT99), .Z(n525) );
  NAND2_X1 U626 ( .A1(G214), .A2(n523), .ZN(n524) );
  XNOR2_X1 U627 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U628 ( .A(n527), .B(n526), .Z(n528) );
  XNOR2_X1 U629 ( .A(n529), .B(n528), .ZN(n672) );
  NOR2_X1 U630 ( .A1(G902), .A2(n672), .ZN(n533) );
  XNOR2_X1 U631 ( .A(KEYINPUT13), .B(KEYINPUT100), .ZN(n531) );
  INV_X1 U632 ( .A(G475), .ZN(n530) );
  INV_X1 U633 ( .A(G217), .ZN(n534) );
  NOR2_X1 U634 ( .A1(n535), .A2(n534), .ZN(n537) );
  XOR2_X1 U635 ( .A(KEYINPUT102), .B(KEYINPUT9), .Z(n536) );
  XNOR2_X1 U636 ( .A(n537), .B(n536), .ZN(n545) );
  XNOR2_X1 U637 ( .A(n538), .B(G107), .ZN(n539) );
  XNOR2_X1 U638 ( .A(n377), .B(n539), .ZN(n543) );
  INV_X1 U639 ( .A(n576), .ZN(n571) );
  AND2_X1 U640 ( .A1(n577), .A2(n571), .ZN(n766) );
  NAND2_X1 U641 ( .A1(n583), .A2(n766), .ZN(n661) );
  XNOR2_X1 U642 ( .A(n661), .B(G134), .ZN(G36) );
  INV_X1 U643 ( .A(KEYINPUT6), .ZN(n549) );
  INV_X1 U644 ( .A(KEYINPUT104), .ZN(n550) );
  XNOR2_X2 U645 ( .A(n551), .B(n550), .ZN(n764) );
  INV_X1 U646 ( .A(n764), .ZN(n761) );
  INV_X1 U647 ( .A(n552), .ZN(n723) );
  NAND2_X1 U648 ( .A1(n610), .A2(n555), .ZN(n556) );
  INV_X1 U649 ( .A(n711), .ZN(n557) );
  NOR2_X1 U650 ( .A1(n363), .A2(n557), .ZN(n558) );
  NAND2_X1 U651 ( .A1(n587), .A2(n558), .ZN(n559) );
  XNOR2_X1 U652 ( .A(n559), .B(KEYINPUT43), .ZN(n560) );
  INV_X1 U653 ( .A(n514), .ZN(n645) );
  NAND2_X1 U654 ( .A1(n560), .A2(n645), .ZN(n659) );
  XNOR2_X1 U655 ( .A(n659), .B(G140), .ZN(G42) );
  INV_X1 U656 ( .A(G898), .ZN(n774) );
  NAND2_X1 U657 ( .A1(G953), .A2(n774), .ZN(n770) );
  OR2_X1 U658 ( .A1(n564), .A2(n770), .ZN(n565) );
  AND2_X1 U659 ( .A1(n566), .A2(n565), .ZN(n567) );
  INV_X1 U660 ( .A(n577), .ZN(n572) );
  NAND2_X1 U661 ( .A1(n572), .A2(n571), .ZN(n646) );
  INV_X1 U662 ( .A(n646), .ZN(n573) );
  INV_X1 U663 ( .A(KEYINPUT35), .ZN(n574) );
  BUF_X2 U664 ( .A(n606), .Z(n599) );
  XNOR2_X1 U665 ( .A(G122), .B(KEYINPUT126), .ZN(n575) );
  XNOR2_X1 U666 ( .A(n359), .B(n575), .ZN(G24) );
  NAND2_X1 U667 ( .A1(n577), .A2(n576), .ZN(n715) );
  INV_X1 U668 ( .A(KEYINPUT22), .ZN(n578) );
  XNOR2_X2 U669 ( .A(n579), .B(n578), .ZN(n597) );
  INV_X1 U670 ( .A(n363), .ZN(n594) );
  INV_X1 U671 ( .A(n726), .ZN(n628) );
  NAND2_X1 U672 ( .A1(n612), .A2(n628), .ZN(n581) );
  INV_X1 U673 ( .A(KEYINPUT66), .ZN(n580) );
  XNOR2_X1 U674 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U675 ( .A(n608), .B(G110), .ZN(G12) );
  BUF_X1 U676 ( .A(n585), .Z(n586) );
  NAND2_X1 U677 ( .A1(n587), .A2(n586), .ZN(n590) );
  INV_X1 U678 ( .A(KEYINPUT90), .ZN(n588) );
  XNOR2_X1 U679 ( .A(n588), .B(KEYINPUT36), .ZN(n589) );
  XNOR2_X1 U680 ( .A(n590), .B(n589), .ZN(n591) );
  XOR2_X1 U681 ( .A(G125), .B(KEYINPUT37), .Z(n592) );
  XNOR2_X1 U682 ( .A(n641), .B(n592), .ZN(G27) );
  OR2_X1 U683 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U684 ( .A1(n610), .A2(n595), .ZN(n596) );
  NAND2_X1 U685 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U686 ( .A(n598), .B(KEYINPUT32), .ZN(n607) );
  XNOR2_X1 U687 ( .A(n607), .B(G119), .ZN(G21) );
  INV_X1 U688 ( .A(n599), .ZN(n600) );
  NAND2_X1 U689 ( .A1(n600), .A2(KEYINPUT69), .ZN(n604) );
  INV_X1 U690 ( .A(KEYINPUT69), .ZN(n605) );
  AND2_X1 U691 ( .A1(n606), .A2(n605), .ZN(n602) );
  INV_X1 U692 ( .A(KEYINPUT44), .ZN(n601) );
  NAND2_X1 U693 ( .A1(n602), .A2(n601), .ZN(n603) );
  NAND2_X1 U694 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U695 ( .A1(n362), .A2(n726), .ZN(n734) );
  XOR2_X1 U696 ( .A(KEYINPUT97), .B(KEYINPUT31), .Z(n615) );
  XNOR2_X1 U697 ( .A(n616), .B(n615), .ZN(n767) );
  OR2_X1 U698 ( .A1(n617), .A2(n726), .ZN(n618) );
  OR2_X1 U699 ( .A1(n767), .A2(n364), .ZN(n622) );
  INV_X1 U700 ( .A(KEYINPUT105), .ZN(n620) );
  INV_X1 U701 ( .A(n766), .ZN(n757) );
  AND2_X1 U702 ( .A1(n761), .A2(n757), .ZN(n619) );
  XNOR2_X1 U703 ( .A(n620), .B(n619), .ZN(n717) );
  XNOR2_X1 U704 ( .A(n717), .B(KEYINPUT83), .ZN(n621) );
  NAND2_X1 U705 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U706 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n625) );
  XNOR2_X1 U707 ( .A(n626), .B(KEYINPUT85), .ZN(n663) );
  NAND2_X1 U708 ( .A1(n712), .A2(n711), .ZN(n716) );
  NOR2_X1 U709 ( .A1(n716), .A2(n715), .ZN(n627) );
  XNOR2_X1 U710 ( .A(n627), .B(KEYINPUT41), .ZN(n744) );
  NOR2_X1 U711 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U712 ( .A(KEYINPUT28), .B(n630), .ZN(n632) );
  NAND2_X1 U713 ( .A1(n632), .A2(n380), .ZN(n639) );
  INV_X1 U714 ( .A(KEYINPUT46), .ZN(n633) );
  XNOR2_X1 U715 ( .A(n634), .B(n633), .ZN(n654) );
  INV_X1 U716 ( .A(n717), .ZN(n643) );
  NOR2_X1 U717 ( .A1(KEYINPUT83), .A2(KEYINPUT47), .ZN(n635) );
  NAND2_X1 U718 ( .A1(n643), .A2(n635), .ZN(n637) );
  NAND2_X1 U719 ( .A1(n717), .A2(KEYINPUT83), .ZN(n636) );
  NAND2_X1 U720 ( .A1(n637), .A2(n636), .ZN(n640) );
  NOR2_X1 U721 ( .A1(n639), .A2(n361), .ZN(n756) );
  NAND2_X1 U722 ( .A1(n640), .A2(n756), .ZN(n642) );
  NAND2_X1 U723 ( .A1(n642), .A2(n641), .ZN(n652) );
  NAND2_X1 U724 ( .A1(n756), .A2(n643), .ZN(n644) );
  NAND2_X1 U725 ( .A1(n644), .A2(KEYINPUT47), .ZN(n650) );
  NOR2_X1 U726 ( .A1(n646), .A2(n645), .ZN(n647) );
  AND2_X1 U727 ( .A1(n648), .A2(n647), .ZN(n760) );
  INV_X1 U728 ( .A(n760), .ZN(n649) );
  NAND2_X1 U729 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U730 ( .A1(n654), .A2(n653), .ZN(n658) );
  XNOR2_X1 U731 ( .A(KEYINPUT89), .B(KEYINPUT48), .ZN(n656) );
  INV_X1 U732 ( .A(KEYINPUT73), .ZN(n655) );
  XNOR2_X1 U733 ( .A(n656), .B(n655), .ZN(n657) );
  INV_X1 U734 ( .A(KEYINPUT88), .ZN(n660) );
  NAND2_X1 U735 ( .A1(n664), .A2(KEYINPUT2), .ZN(n665) );
  NAND2_X1 U736 ( .A1(n705), .A2(KEYINPUT2), .ZN(n666) );
  XNOR2_X1 U737 ( .A(n666), .B(KEYINPUT87), .ZN(n669) );
  BUF_X1 U738 ( .A(n667), .Z(n668) );
  NAND2_X1 U739 ( .A1(n669), .A2(n668), .ZN(n709) );
  XNOR2_X1 U740 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n670) );
  XNOR2_X1 U741 ( .A(n670), .B(KEYINPUT59), .ZN(n671) );
  NAND2_X1 U742 ( .A1(n688), .A2(G210), .ZN(n678) );
  BUF_X1 U743 ( .A(n674), .Z(n675) );
  XOR2_X1 U744 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n676) );
  XNOR2_X1 U745 ( .A(n678), .B(n677), .ZN(n679) );
  NOR2_X2 U746 ( .A1(n679), .A2(n703), .ZN(n680) );
  XNOR2_X1 U747 ( .A(n680), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U748 ( .A1(n688), .A2(G472), .ZN(n683) );
  XNOR2_X1 U749 ( .A(n683), .B(n682), .ZN(n684) );
  NOR2_X2 U750 ( .A1(n684), .A2(n703), .ZN(n687) );
  XNOR2_X1 U751 ( .A(KEYINPUT111), .B(KEYINPUT63), .ZN(n685) );
  XNOR2_X1 U752 ( .A(n685), .B(KEYINPUT92), .ZN(n686) );
  XNOR2_X1 U753 ( .A(n687), .B(n686), .ZN(G57) );
  NAND2_X1 U754 ( .A1(n696), .A2(G217), .ZN(n690) );
  XNOR2_X1 U755 ( .A(n690), .B(n689), .ZN(n691) );
  NOR2_X1 U756 ( .A1(n691), .A2(n703), .ZN(G66) );
  NAND2_X1 U757 ( .A1(n696), .A2(G478), .ZN(n694) );
  XOR2_X1 U758 ( .A(n692), .B(KEYINPUT123), .Z(n693) );
  XNOR2_X1 U759 ( .A(n694), .B(n693), .ZN(n695) );
  NOR2_X1 U760 ( .A1(n695), .A2(n703), .ZN(G63) );
  NAND2_X1 U761 ( .A1(n696), .A2(G469), .ZN(n702) );
  XOR2_X1 U762 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n698) );
  XNOR2_X1 U763 ( .A(n698), .B(KEYINPUT120), .ZN(n699) );
  XNOR2_X1 U764 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U765 ( .A(n702), .B(n701), .ZN(n704) );
  NOR2_X1 U766 ( .A1(n704), .A2(n703), .ZN(G54) );
  NAND2_X1 U767 ( .A1(n705), .A2(n668), .ZN(n707) );
  INV_X1 U768 ( .A(KEYINPUT2), .ZN(n706) );
  NAND2_X1 U769 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U770 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U771 ( .A(n710), .B(KEYINPUT86), .ZN(n750) );
  NOR2_X1 U772 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U773 ( .A(n713), .B(KEYINPUT116), .ZN(n714) );
  NOR2_X1 U774 ( .A1(n715), .A2(n714), .ZN(n719) );
  NOR2_X1 U775 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U776 ( .A1(n719), .A2(n718), .ZN(n721) );
  NOR2_X1 U777 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U778 ( .A(KEYINPUT117), .B(n722), .Z(n739) );
  XNOR2_X1 U779 ( .A(n724), .B(KEYINPUT49), .ZN(n725) );
  NOR2_X1 U780 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U781 ( .A(KEYINPUT113), .B(n727), .Z(n733) );
  XOR2_X1 U782 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n730) );
  NOR2_X1 U783 ( .A1(n363), .A2(n728), .ZN(n729) );
  XOR2_X1 U784 ( .A(n730), .B(n729), .Z(n731) );
  XNOR2_X1 U785 ( .A(KEYINPUT114), .B(n731), .ZN(n732) );
  NAND2_X1 U786 ( .A1(n733), .A2(n732), .ZN(n735) );
  NAND2_X1 U787 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U788 ( .A(KEYINPUT51), .B(n736), .ZN(n737) );
  NOR2_X1 U789 ( .A1(n744), .A2(n737), .ZN(n738) );
  NOR2_X1 U790 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U791 ( .A(n740), .B(KEYINPUT118), .ZN(n741) );
  XNOR2_X1 U792 ( .A(KEYINPUT52), .B(n741), .ZN(n742) );
  NOR2_X1 U793 ( .A1(n743), .A2(n742), .ZN(n746) );
  NOR2_X1 U794 ( .A1(n744), .A2(n720), .ZN(n745) );
  NOR2_X1 U795 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U796 ( .A(KEYINPUT119), .B(n747), .ZN(n748) );
  NOR2_X1 U797 ( .A1(n748), .A2(G953), .ZN(n749) );
  NAND2_X1 U798 ( .A1(n750), .A2(n749), .ZN(n751) );
  XOR2_X1 U799 ( .A(KEYINPUT53), .B(n751), .Z(G75) );
  NAND2_X1 U800 ( .A1(n364), .A2(n764), .ZN(n752) );
  XNOR2_X1 U801 ( .A(n752), .B(G104), .ZN(G6) );
  XOR2_X1 U802 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n754) );
  NAND2_X1 U803 ( .A1(n364), .A2(n766), .ZN(n753) );
  XNOR2_X1 U804 ( .A(n754), .B(n753), .ZN(n755) );
  XNOR2_X1 U805 ( .A(G107), .B(n755), .ZN(G9) );
  INV_X1 U806 ( .A(n756), .ZN(n762) );
  NOR2_X1 U807 ( .A1(n762), .A2(n757), .ZN(n759) );
  XNOR2_X1 U808 ( .A(G128), .B(KEYINPUT29), .ZN(n758) );
  XNOR2_X1 U809 ( .A(n759), .B(n758), .ZN(G30) );
  XOR2_X1 U810 ( .A(G143), .B(n760), .Z(G45) );
  NOR2_X1 U811 ( .A1(n762), .A2(n761), .ZN(n763) );
  XOR2_X1 U812 ( .A(G146), .B(n763), .Z(G48) );
  NAND2_X1 U813 ( .A1(n767), .A2(n764), .ZN(n765) );
  XNOR2_X1 U814 ( .A(n396), .B(n765), .ZN(G15) );
  NAND2_X1 U815 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U816 ( .A(n768), .B(KEYINPUT112), .ZN(n769) );
  XNOR2_X1 U817 ( .A(G116), .B(n769), .ZN(G18) );
  NAND2_X1 U818 ( .A1(n771), .A2(n770), .ZN(n780) );
  NAND2_X1 U819 ( .A1(G953), .A2(G224), .ZN(n772) );
  XOR2_X1 U820 ( .A(KEYINPUT61), .B(n772), .Z(n773) );
  NOR2_X1 U821 ( .A1(n774), .A2(n773), .ZN(n778) );
  NAND2_X1 U822 ( .A1(n668), .A2(n775), .ZN(n776) );
  XOR2_X1 U823 ( .A(KEYINPUT124), .B(n776), .Z(n777) );
  NOR2_X1 U824 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U825 ( .A(n780), .B(n779), .ZN(G69) );
  XNOR2_X1 U826 ( .A(n781), .B(n782), .ZN(n785) );
  NOR2_X1 U827 ( .A1(n783), .A2(G953), .ZN(n784) );
  XNOR2_X1 U828 ( .A(n784), .B(KEYINPUT125), .ZN(n789) );
  XOR2_X1 U829 ( .A(G227), .B(n785), .Z(n786) );
  NAND2_X1 U830 ( .A1(n786), .A2(G900), .ZN(n787) );
  NAND2_X1 U831 ( .A1(n787), .A2(G953), .ZN(n788) );
  NAND2_X1 U832 ( .A1(n789), .A2(n788), .ZN(G72) );
  XNOR2_X1 U833 ( .A(G137), .B(KEYINPUT127), .ZN(n791) );
  XNOR2_X1 U834 ( .A(n791), .B(n790), .ZN(G39) );
endmodule

