//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 1 1 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n825, new_n826, new_n828, new_n829,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952;
  INV_X1    g000(.A(KEYINPUT82), .ZN(new_n202));
  XNOR2_X1  g001(.A(G1gat), .B(G29gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT0), .ZN(new_n204));
  XNOR2_X1  g003(.A(G57gat), .B(G85gat), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  NAND2_X1  g005(.A1(G225gat), .A2(G233gat), .ZN(new_n207));
  INV_X1    g006(.A(G155gat), .ZN(new_n208));
  INV_X1    g007(.A(G162gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT2), .B1(new_n208), .B2(new_n209), .ZN(new_n213));
  XNOR2_X1  g012(.A(G141gat), .B(G148gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n213), .B1(new_n214), .B2(KEYINPUT72), .ZN(new_n215));
  INV_X1    g014(.A(G148gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G141gat), .ZN(new_n217));
  INV_X1    g016(.A(G141gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G148gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT72), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n212), .B1(new_n215), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT73), .B(G141gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n217), .B1(new_n224), .B2(new_n216), .ZN(new_n225));
  INV_X1    g024(.A(new_n212), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(new_n226), .A3(new_n213), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n223), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G120gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G113gat), .ZN(new_n230));
  INV_X1    g029(.A(G113gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G120gat), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT1), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(G127gat), .B(G134gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT68), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n234), .A2(new_n235), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n233), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G134gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n239), .A2(G127gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n233), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT67), .B(G134gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G127gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n238), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n228), .A2(new_n245), .A3(KEYINPUT4), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT4), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n234), .B(new_n235), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n248), .A2(new_n233), .B1(new_n243), .B2(new_n241), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n223), .A2(new_n227), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n247), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT74), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n223), .A2(new_n227), .A3(KEYINPUT74), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n254), .A2(KEYINPUT3), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n223), .A2(new_n227), .A3(new_n257), .ZN(new_n258));
  AND2_X1   g057(.A1(new_n258), .A2(new_n249), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n252), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n254), .A2(new_n255), .A3(new_n249), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT75), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n262), .B1(new_n228), .B2(new_n245), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n207), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n254), .A2(new_n262), .A3(new_n255), .A4(new_n249), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n207), .A2(new_n260), .B1(new_n267), .B2(KEYINPUT5), .ZN(new_n268));
  AND2_X1   g067(.A1(new_n246), .A2(new_n251), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n256), .A2(new_n259), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(new_n270), .A3(new_n207), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT5), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n206), .B1(new_n268), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT6), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n267), .A2(KEYINPUT5), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(new_n271), .ZN(new_n277));
  INV_X1    g076(.A(new_n206), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n260), .A2(KEYINPUT5), .A3(new_n207), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n274), .A2(new_n275), .A3(new_n280), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n277), .A2(KEYINPUT6), .A3(new_n278), .A4(new_n279), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G226gat), .A2(G233gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(G169gat), .A2(G176gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT23), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT23), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n287), .B1(G169gat), .B2(G176gat), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n286), .B1(new_n288), .B2(new_n285), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT25), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(G183gat), .A2(G190gat), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n293), .B1(KEYINPUT65), .B2(KEYINPUT24), .ZN(new_n294));
  AND2_X1   g093(.A1(KEYINPUT65), .A2(KEYINPUT24), .ZN(new_n295));
  OAI221_X1 g094(.A(new_n292), .B1(G183gat), .B2(G190gat), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n292), .B1(G183gat), .B2(G190gat), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n298), .B1(new_n301), .B2(new_n289), .ZN(new_n302));
  INV_X1    g101(.A(G183gat), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT27), .B1(new_n303), .B2(KEYINPUT66), .ZN(new_n304));
  INV_X1    g103(.A(G190gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT27), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G183gat), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n304), .B(new_n305), .C1(KEYINPUT66), .C2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT28), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT27), .B(G183gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n311), .A2(KEYINPUT28), .A3(new_n305), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G169gat), .ZN(new_n314));
  INV_X1    g113(.A(G176gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT26), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n316), .B1(new_n317), .B2(new_n285), .ZN(new_n318));
  OAI21_X1  g117(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n318), .A2(new_n319), .B1(G183gat), .B2(G190gat), .ZN(new_n320));
  AOI22_X1  g119(.A1(new_n297), .A2(new_n302), .B1(new_n313), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n284), .B1(new_n321), .B2(KEYINPUT29), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n313), .A2(new_n320), .ZN(new_n323));
  OAI221_X1 g122(.A(new_n286), .B1(new_n288), .B2(new_n285), .C1(new_n299), .C2(new_n300), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n324), .A2(new_n298), .B1(new_n291), .B2(new_n296), .ZN(new_n325));
  OAI211_X1 g124(.A(G226gat), .B(G233gat), .C1(new_n323), .C2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G197gat), .B(G204gat), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT22), .ZN(new_n329));
  INV_X1    g128(.A(G211gat), .ZN(new_n330));
  INV_X1    g129(.A(G218gat), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(G211gat), .B(G218gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n327), .A2(new_n335), .ZN(new_n336));
  XOR2_X1   g135(.A(G8gat), .B(G36gat), .Z(new_n337));
  XNOR2_X1  g136(.A(new_n337), .B(KEYINPUT70), .ZN(new_n338));
  XNOR2_X1  g137(.A(G64gat), .B(G92gat), .ZN(new_n339));
  XOR2_X1   g138(.A(new_n338), .B(new_n339), .Z(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n335), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n322), .A2(new_n326), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n336), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT71), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT30), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n336), .A2(new_n343), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(new_n340), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT30), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n344), .A2(KEYINPUT71), .A3(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n346), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n283), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT76), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n351), .B1(new_n281), .B2(new_n282), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(G228gat), .A2(G233gat), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n257), .B1(new_n335), .B2(KEYINPUT29), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n359), .A2(new_n250), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT29), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n342), .B1(new_n258), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n358), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n258), .A2(new_n361), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n358), .B1(new_n364), .B2(new_n335), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n359), .A2(new_n254), .A3(new_n255), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT77), .B1(new_n363), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G22gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(G78gat), .B(G106gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(KEYINPUT31), .B(G50gat), .ZN(new_n372));
  XOR2_X1   g171(.A(new_n371), .B(new_n372), .Z(new_n373));
  NAND3_X1  g172(.A1(new_n369), .A2(new_n370), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n373), .ZN(new_n375));
  OAI21_X1  g174(.A(G22gat), .B1(new_n368), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n363), .A2(KEYINPUT77), .A3(new_n367), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n367), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT77), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n374), .A2(new_n376), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n354), .A2(new_n357), .A3(new_n384), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n281), .A2(new_n282), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT38), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n341), .B1(new_n347), .B2(KEYINPUT37), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT37), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n336), .A2(new_n389), .A3(new_n343), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n387), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  OR2_X1    g190(.A1(new_n391), .A2(KEYINPUT80), .ZN(new_n392));
  INV_X1    g191(.A(new_n343), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n342), .B1(new_n322), .B2(new_n326), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT37), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n395), .A2(new_n390), .A3(new_n387), .A4(new_n340), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n344), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n397), .B1(KEYINPUT80), .B2(new_n391), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n386), .A2(new_n392), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT78), .ZN(new_n400));
  AOI211_X1 g199(.A(KEYINPUT39), .B(new_n207), .C1(new_n269), .C2(new_n270), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n400), .B1(new_n401), .B2(new_n278), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n269), .A2(new_n270), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n265), .ZN(new_n404));
  OAI211_X1 g203(.A(KEYINPUT78), .B(new_n206), .C1(new_n404), .C2(KEYINPUT39), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n265), .B1(new_n264), .B2(new_n266), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT79), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT39), .ZN(new_n409));
  OR3_X1    g208(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n408), .B1(new_n407), .B2(new_n409), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(new_n411), .A3(new_n404), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT40), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n406), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n413), .B1(new_n406), .B2(new_n412), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n280), .B(new_n351), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n374), .A2(new_n376), .A3(new_n382), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n382), .B1(new_n374), .B2(new_n376), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n399), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT34), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n421), .A2(KEYINPUT69), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n245), .B1(new_n323), .B2(new_n325), .ZN(new_n424));
  NAND2_X1  g223(.A1(G227gat), .A2(G233gat), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n297), .A2(new_n302), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n313), .A2(new_n320), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(new_n249), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n424), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT32), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT33), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  XOR2_X1   g232(.A(G15gat), .B(G43gat), .Z(new_n434));
  XNOR2_X1  g233(.A(G71gat), .B(G99gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n434), .B(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n431), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n436), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n430), .B(KEYINPUT32), .C1(new_n432), .C2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n429), .ZN(new_n440));
  AOI22_X1  g239(.A1(new_n440), .A2(new_n425), .B1(KEYINPUT69), .B2(new_n421), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n437), .A2(new_n439), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n442), .B1(new_n437), .B2(new_n439), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n423), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n437), .A2(new_n439), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n441), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n437), .A2(new_n439), .A3(new_n442), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(new_n422), .A3(new_n448), .ZN(new_n449));
  AND2_X1   g248(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT36), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n445), .A2(new_n449), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT36), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n385), .A2(new_n420), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT35), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n354), .A2(new_n357), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n450), .A2(new_n384), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT81), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n459), .A2(new_n461), .A3(new_n457), .A4(new_n355), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n419), .A2(new_n457), .A3(new_n452), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT81), .B1(new_n463), .B2(new_n353), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n202), .B(new_n456), .C1(new_n460), .C2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n419), .A2(new_n452), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n468), .B1(new_n354), .B2(new_n357), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n464), .B(new_n462), .C1(new_n469), .C2(new_n457), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n202), .B1(new_n470), .B2(new_n456), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(G113gat), .B(G141gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(G169gat), .B(G197gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n473), .B(new_n474), .ZN(new_n475));
  XOR2_X1   g274(.A(KEYINPUT83), .B(KEYINPUT11), .Z(new_n476));
  XNOR2_X1  g275(.A(new_n475), .B(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n477), .B(KEYINPUT12), .ZN(new_n478));
  NAND2_X1  g277(.A1(G229gat), .A2(G233gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(G15gat), .B(G22gat), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT90), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n482), .B(G8gat), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT16), .ZN(new_n484));
  AOI21_X1  g283(.A(G1gat), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n483), .B(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(G36gat), .ZN(new_n487));
  INV_X1    g286(.A(G29gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT87), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT87), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(G29gat), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n487), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT85), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI211_X1 g294(.A(KEYINPUT85), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OR3_X1    g296(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n492), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(G43gat), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n500), .A2(G50gat), .ZN(new_n501));
  INV_X1    g300(.A(G50gat), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n502), .A2(G43gat), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT84), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(G43gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n500), .A2(G50gat), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT84), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n504), .A2(KEYINPUT15), .A3(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT15), .ZN(new_n510));
  OR2_X1    g309(.A1(KEYINPUT88), .A2(G50gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(KEYINPUT88), .A2(G50gat), .ZN(new_n512));
  AOI21_X1  g311(.A(G43gat), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n510), .B1(new_n513), .B2(new_n501), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n499), .A2(new_n509), .A3(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT86), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n495), .A2(new_n516), .A3(new_n496), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n516), .B1(new_n495), .B2(new_n496), .ZN(new_n518));
  NOR3_X1   g317(.A1(new_n517), .A2(new_n518), .A3(new_n492), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n504), .A2(KEYINPUT15), .A3(new_n498), .A4(new_n508), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n515), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n486), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT17), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT91), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n509), .A2(new_n514), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n497), .A2(KEYINPUT86), .ZN(new_n526));
  INV_X1    g325(.A(new_n492), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n495), .A2(new_n516), .A3(new_n496), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n520), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n525), .A2(new_n499), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT91), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(new_n532), .A3(KEYINPUT17), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT89), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n529), .A2(new_n530), .ZN(new_n535));
  AOI211_X1 g334(.A(new_n534), .B(KEYINPUT17), .C1(new_n535), .C2(new_n515), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT89), .B1(new_n521), .B2(new_n523), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n524), .B(new_n533), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n479), .B(new_n522), .C1(new_n538), .C2(new_n486), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT94), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n478), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n534), .B1(new_n531), .B2(KEYINPUT17), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n521), .A2(KEYINPUT89), .A3(new_n523), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n486), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n546), .A2(new_n547), .A3(new_n524), .A4(new_n533), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n548), .A2(KEYINPUT18), .A3(new_n479), .A4(new_n522), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n486), .B(new_n521), .ZN(new_n550));
  XOR2_X1   g349(.A(KEYINPUT93), .B(KEYINPUT13), .Z(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(new_n479), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n541), .A2(new_n549), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n543), .A2(new_n554), .ZN(new_n555));
  AOI22_X1  g354(.A1(new_n539), .A2(new_n540), .B1(new_n550), .B2(new_n552), .ZN(new_n556));
  AOI21_X1  g355(.A(KEYINPUT94), .B1(new_n539), .B2(new_n540), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n556), .B(new_n549), .C1(new_n557), .C2(new_n478), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(G57gat), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n561), .A2(G64gat), .ZN(new_n562));
  INV_X1    g361(.A(G64gat), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n563), .A2(G57gat), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT95), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(G57gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n561), .A2(G64gat), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT95), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n565), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G71gat), .B(G78gat), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT96), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT96), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n572), .A2(new_n577), .A3(new_n574), .ZN(new_n578));
  XNOR2_X1  g377(.A(KEYINPUT97), .B(G57gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(G64gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(new_n566), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n574), .A2(new_n570), .ZN(new_n582));
  AOI22_X1  g381(.A1(new_n576), .A2(new_n578), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n583), .A2(KEYINPUT21), .ZN(new_n584));
  AND2_X1   g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT99), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n486), .B1(KEYINPUT21), .B2(new_n583), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n586), .B(KEYINPUT99), .ZN(new_n591));
  INV_X1    g390(.A(new_n589), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(KEYINPUT98), .B(KEYINPUT19), .Z(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT20), .ZN(new_n595));
  XOR2_X1   g394(.A(G127gat), .B(G155gat), .Z(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(G183gat), .B(G211gat), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n590), .A2(new_n593), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n599), .B1(new_n590), .B2(new_n593), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(G85gat), .A2(G92gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT7), .ZN(new_n604));
  XNOR2_X1  g403(.A(G99gat), .B(G106gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(G99gat), .A2(G106gat), .ZN(new_n606));
  INV_X1    g405(.A(G85gat), .ZN(new_n607));
  INV_X1    g406(.A(G92gat), .ZN(new_n608));
  AOI22_X1  g407(.A1(KEYINPUT8), .A2(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AND3_X1   g408(.A1(new_n604), .A2(new_n605), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n605), .B1(new_n604), .B2(new_n609), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n521), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n613), .B(new_n614), .C1(new_n538), .C2(new_n612), .ZN(new_n615));
  XNOR2_X1  g414(.A(G190gat), .B(G218gat), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(KEYINPUT100), .B1(new_n615), .B2(new_n617), .ZN(new_n619));
  XNOR2_X1  g418(.A(G134gat), .B(G162gat), .ZN(new_n620));
  AOI21_X1  g419(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n620), .B(new_n621), .Z(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  OR3_X1    g422(.A1(new_n618), .A2(new_n619), .A3(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n623), .B1(new_n618), .B2(new_n619), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n581), .A2(new_n582), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n572), .A2(new_n577), .A3(new_n574), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n577), .B1(new_n572), .B2(new_n574), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n612), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT10), .ZN(new_n634));
  OAI211_X1 g433(.A(new_n628), .B(new_n612), .C1(new_n629), .C2(new_n630), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT101), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n583), .A2(new_n637), .A3(KEYINPUT10), .A4(new_n612), .ZN(new_n638));
  OAI21_X1  g437(.A(KEYINPUT101), .B1(new_n635), .B2(new_n634), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G230gat), .A2(G233gat), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n633), .A2(new_n635), .ZN(new_n643));
  INV_X1    g442(.A(new_n641), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G120gat), .B(G148gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(G176gat), .B(G204gat), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n647), .B(new_n648), .Z(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n642), .A2(new_n645), .A3(new_n649), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n602), .A2(new_n627), .A3(new_n654), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n472), .A2(new_n560), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n386), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(G1gat), .ZN(G1324gat));
  NOR4_X1   g457(.A1(new_n472), .A2(new_n560), .A3(new_n352), .A4(new_n655), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT102), .B(KEYINPUT16), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(G8gat), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT42), .ZN(new_n663));
  OR3_X1    g462(.A1(new_n662), .A2(KEYINPUT103), .A3(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(KEYINPUT103), .B1(new_n662), .B2(new_n663), .ZN(new_n665));
  INV_X1    g464(.A(new_n662), .ZN(new_n666));
  INV_X1    g465(.A(new_n659), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n663), .B1(new_n667), .B2(G8gat), .ZN(new_n668));
  OAI211_X1 g467(.A(new_n664), .B(new_n665), .C1(new_n666), .C2(new_n668), .ZN(G1325gat));
  INV_X1    g468(.A(G15gat), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n656), .A2(new_n670), .A3(new_n452), .ZN(new_n671));
  INV_X1    g470(.A(new_n455), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n656), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n671), .B1(new_n673), .B2(new_n670), .ZN(G1326gat));
  NAND2_X1  g473(.A1(new_n656), .A2(new_n384), .ZN(new_n675));
  XNOR2_X1  g474(.A(KEYINPUT43), .B(G22gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1327gat));
  NAND2_X1  g476(.A1(new_n489), .A2(new_n491), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n627), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n680), .B1(new_n467), .B2(new_n471), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n470), .A2(new_n456), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n626), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n679), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n602), .B(KEYINPUT105), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n653), .B(KEYINPUT106), .Z(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n686), .A2(new_n560), .A3(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n681), .A2(new_n684), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n678), .B1(new_n690), .B2(new_n283), .ZN(new_n691));
  INV_X1    g490(.A(new_n471), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n466), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n602), .A2(new_n627), .A3(new_n653), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n693), .A2(new_n559), .A3(new_n694), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n283), .A2(new_n678), .ZN(new_n696));
  OR3_X1    g495(.A1(new_n695), .A2(KEYINPUT104), .A3(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT45), .ZN(new_n698));
  OAI21_X1  g497(.A(KEYINPUT104), .B1(new_n695), .B2(new_n696), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n698), .B1(new_n697), .B2(new_n699), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n691), .B1(new_n700), .B2(new_n701), .ZN(G1328gat));
  NOR3_X1   g501(.A1(new_n695), .A2(G36gat), .A3(new_n352), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT46), .ZN(new_n704));
  OAI21_X1  g503(.A(G36gat), .B1(new_n690), .B2(new_n352), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(G1329gat));
  OAI21_X1  g505(.A(new_n500), .B1(new_n695), .B2(new_n450), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n672), .A2(G43gat), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n707), .B1(new_n690), .B2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g509(.A(new_n695), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n511), .A2(new_n512), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n419), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT107), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n681), .A2(new_n684), .A3(new_n384), .A4(new_n689), .ZN(new_n715));
  AOI22_X1  g514(.A1(new_n711), .A2(new_n714), .B1(new_n715), .B2(new_n712), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT48), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n716), .A2(KEYINPUT108), .A3(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(KEYINPUT108), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n717), .A2(KEYINPUT108), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n716), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n718), .A2(new_n721), .ZN(G1331gat));
  INV_X1    g521(.A(new_n601), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n590), .A2(new_n593), .A3(new_n599), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR4_X1   g524(.A1(new_n725), .A2(new_n687), .A3(new_n559), .A4(new_n626), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n682), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(new_n283), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(new_n579), .ZN(G1332gat));
  NOR2_X1   g528(.A1(new_n727), .A2(new_n352), .ZN(new_n730));
  NOR2_X1   g529(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n731));
  AND2_X1   g530(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n733), .B1(new_n730), .B2(new_n731), .ZN(G1333gat));
  NOR3_X1   g533(.A1(new_n727), .A2(G71gat), .A3(new_n450), .ZN(new_n735));
  INV_X1    g534(.A(new_n727), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n672), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n735), .B1(G71gat), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g538(.A1(new_n736), .A2(new_n384), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g540(.A1(new_n602), .A2(new_n559), .A3(new_n654), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n681), .A2(new_n684), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(KEYINPUT109), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT109), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n681), .A2(new_n684), .A3(new_n745), .A4(new_n742), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n744), .A2(new_n386), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT110), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT110), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n744), .A2(new_n749), .A3(new_n386), .A4(new_n746), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n748), .A2(G85gat), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n627), .B1(new_n470), .B2(new_n456), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n602), .A2(new_n559), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n756), .A2(new_n607), .A3(new_n386), .A4(new_n653), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n751), .A2(new_n757), .ZN(G1336gat));
  NOR3_X1   g557(.A1(new_n687), .A2(G92gat), .A3(new_n352), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(G92gat), .B1(new_n743), .B2(new_n352), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n744), .A2(new_n351), .A3(new_n746), .ZN(new_n764));
  NOR2_X1   g563(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n754), .B(new_n765), .ZN(new_n766));
  AOI22_X1  g565(.A1(new_n764), .A2(G92gat), .B1(new_n766), .B2(new_n759), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n763), .B1(new_n767), .B2(new_n762), .ZN(G1337gat));
  NAND3_X1  g567(.A1(new_n744), .A2(new_n672), .A3(new_n746), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G99gat), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n450), .A2(G99gat), .A3(new_n654), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(G1338gat));
  NOR3_X1   g572(.A1(new_n687), .A2(G106gat), .A3(new_n419), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT53), .B1(new_n756), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(KEYINPUT112), .B1(new_n743), .B2(new_n419), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(G106gat), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n743), .A2(KEYINPUT112), .A3(new_n419), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n775), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n744), .A2(new_n384), .A3(new_n746), .ZN(new_n780));
  AOI22_X1  g579(.A1(new_n780), .A2(G106gat), .B1(new_n766), .B2(new_n774), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n779), .B1(new_n781), .B2(new_n782), .ZN(G1339gat));
  AND2_X1   g582(.A1(new_n636), .A2(new_n639), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n784), .A2(KEYINPUT113), .A3(new_n644), .A4(new_n638), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n786), .B1(new_n640), .B2(new_n641), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n788), .B1(new_n640), .B2(new_n641), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n785), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n640), .A2(new_n788), .A3(new_n641), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n791), .A2(new_n650), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(KEYINPUT55), .A3(new_n792), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n793), .A2(new_n652), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT55), .B1(new_n790), .B2(new_n792), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n794), .A2(new_n559), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n556), .A2(new_n478), .A3(new_n549), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n479), .B1(new_n548), .B2(new_n522), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n550), .A2(new_n552), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n477), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n653), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n626), .B1(new_n797), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n793), .A2(new_n652), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n805), .A2(new_n795), .ZN(new_n806));
  AND3_X1   g605(.A1(new_n806), .A2(new_n626), .A3(new_n802), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT114), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT114), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n806), .A2(new_n626), .A3(new_n802), .ZN(new_n810));
  AOI22_X1  g609(.A1(new_n806), .A2(new_n559), .B1(new_n653), .B2(new_n802), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n809), .B(new_n810), .C1(new_n811), .C2(new_n626), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n808), .A2(new_n685), .A3(new_n812), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n725), .A2(new_n626), .A3(new_n653), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n560), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n468), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n283), .A2(new_n351), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n818), .A2(new_n560), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(new_n231), .ZN(G1340gat));
  NOR3_X1   g619(.A1(new_n818), .A2(new_n229), .A3(new_n687), .ZN(new_n821));
  INV_X1    g620(.A(new_n818), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n653), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n821), .B1(new_n229), .B2(new_n823), .ZN(G1341gat));
  OAI21_X1  g623(.A(G127gat), .B1(new_n818), .B2(new_n685), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n725), .A2(G127gat), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n825), .B1(new_n818), .B2(new_n826), .ZN(G1342gat));
  NAND3_X1  g626(.A1(new_n822), .A2(new_n242), .A3(new_n626), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n828), .A2(KEYINPUT56), .ZN(new_n829));
  OAI21_X1  g628(.A(G134gat), .B1(new_n818), .B2(new_n627), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(KEYINPUT56), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(G1343gat));
  XOR2_X1   g631(.A(KEYINPUT73), .B(G141gat), .Z(new_n833));
  NAND2_X1  g632(.A1(new_n455), .A2(new_n817), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n419), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n790), .A2(new_n792), .ZN(new_n837));
  XOR2_X1   g636(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n794), .A2(new_n559), .A3(new_n839), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n840), .A2(new_n803), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n841), .A2(new_n626), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT116), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n807), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n841), .A2(new_n626), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(KEYINPUT116), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n602), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n815), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n836), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n419), .B1(new_n813), .B2(new_n815), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(KEYINPUT57), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n834), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n833), .B1(new_n853), .B2(new_n559), .ZN(new_n854));
  INV_X1    g653(.A(new_n834), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n559), .A2(new_n218), .ZN(new_n858));
  XOR2_X1   g657(.A(new_n858), .B(KEYINPUT117), .Z(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT58), .B1(new_n854), .B2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n836), .ZN(new_n863));
  INV_X1    g662(.A(new_n846), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n810), .B1(new_n845), .B2(KEYINPUT116), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n725), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n863), .B1(new_n866), .B2(new_n815), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n855), .B1(new_n867), .B2(new_n851), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n224), .B1(new_n868), .B2(new_n560), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT58), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n869), .A2(new_n870), .A3(new_n860), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n862), .A2(new_n871), .ZN(G1344gat));
  NAND3_X1  g671(.A1(new_n857), .A2(new_n216), .A3(new_n653), .ZN(new_n873));
  AOI211_X1 g672(.A(KEYINPUT59), .B(new_n216), .C1(new_n853), .C2(new_n653), .ZN(new_n874));
  XNOR2_X1  g673(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n814), .A2(KEYINPUT119), .A3(new_n560), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n877), .B1(new_n655), .B2(new_n559), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n810), .B1(new_n841), .B2(new_n626), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n602), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI211_X1 g681(.A(KEYINPUT120), .B(new_n810), .C1(new_n841), .C2(new_n626), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n879), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n835), .B1(new_n884), .B2(new_n419), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n813), .A2(new_n815), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n836), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(new_n653), .A3(new_n855), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n875), .B1(new_n889), .B2(G148gat), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n873), .B1(new_n874), .B2(new_n890), .ZN(G1345gat));
  NOR3_X1   g690(.A1(new_n868), .A2(new_n208), .A3(new_n685), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n857), .A2(KEYINPUT121), .A3(new_n602), .ZN(new_n893));
  AOI21_X1  g692(.A(KEYINPUT121), .B1(new_n857), .B2(new_n602), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n894), .A2(G155gat), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n892), .B1(new_n893), .B2(new_n895), .ZN(G1346gat));
  AOI21_X1  g695(.A(G162gat), .B1(new_n857), .B2(new_n626), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n627), .A2(new_n209), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n897), .B1(new_n853), .B2(new_n898), .ZN(G1347gat));
  NOR2_X1   g698(.A1(new_n386), .A2(new_n352), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n816), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n901), .A2(new_n560), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(new_n314), .ZN(G1348gat));
  OAI21_X1  g702(.A(G176gat), .B1(new_n901), .B2(new_n687), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n653), .A2(new_n315), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n901), .B2(new_n905), .ZN(G1349gat));
  NAND4_X1  g705(.A1(new_n886), .A2(new_n459), .A3(new_n686), .A4(new_n900), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(G183gat), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n816), .A2(new_n311), .A3(new_n602), .A4(new_n900), .ZN(new_n909));
  OR2_X1    g708(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n910));
  NAND2_X1  g709(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n908), .A2(new_n909), .A3(new_n910), .A4(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n908), .A2(new_n909), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT122), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n908), .A2(KEYINPUT122), .A3(new_n909), .ZN(new_n916));
  AND4_X1   g715(.A1(KEYINPUT123), .A2(new_n915), .A3(KEYINPUT60), .A4(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT60), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n918), .B1(new_n913), .B2(new_n914), .ZN(new_n919));
  AOI21_X1  g718(.A(KEYINPUT123), .B1(new_n919), .B2(new_n916), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n912), .B1(new_n917), .B2(new_n920), .ZN(G1350gat));
  OAI22_X1  g720(.A1(new_n901), .A2(new_n627), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n922));
  NAND2_X1  g721(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n922), .B(new_n923), .ZN(G1351gat));
  AND2_X1   g723(.A1(new_n455), .A2(new_n900), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT126), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n888), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(G197gat), .B1(new_n927), .B2(new_n560), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n850), .A2(new_n925), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT125), .ZN(new_n930));
  INV_X1    g729(.A(G197gat), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n930), .A2(new_n931), .A3(new_n559), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n928), .A2(new_n932), .ZN(G1352gat));
  OAI21_X1  g732(.A(G204gat), .B1(new_n927), .B2(new_n687), .ZN(new_n934));
  INV_X1    g733(.A(G204gat), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n850), .A2(new_n935), .A3(new_n653), .A4(new_n925), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT62), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n934), .A2(new_n938), .A3(KEYINPUT127), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n940));
  INV_X1    g739(.A(new_n926), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n941), .B1(new_n885), .B2(new_n887), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n935), .B1(new_n942), .B2(new_n688), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n940), .B1(new_n943), .B2(new_n937), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n939), .A2(new_n944), .ZN(G1353gat));
  NAND3_X1  g744(.A1(new_n930), .A2(new_n330), .A3(new_n602), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n888), .A2(new_n602), .A3(new_n925), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n947), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n948));
  AOI21_X1  g747(.A(KEYINPUT63), .B1(new_n947), .B2(G211gat), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n946), .B1(new_n948), .B2(new_n949), .ZN(G1354gat));
  OAI21_X1  g749(.A(G218gat), .B1(new_n927), .B2(new_n627), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n930), .A2(new_n331), .A3(new_n626), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1355gat));
endmodule


