//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 1 0 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n434, new_n437, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n569, new_n570, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n632, new_n633, new_n634, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT66), .B(G44), .Z(new_n434));
  INV_X1    g009(.A(new_n434), .ZN(G218));
  INV_X1    g010(.A(G132), .ZN(G219));
  XOR2_X1   g011(.A(KEYINPUT0), .B(G82), .Z(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT67), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n434), .A2(new_n437), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n454), .ZN(new_n458));
  INV_X1    g033(.A(new_n455), .ZN(new_n459));
  AOI22_X1  g034(.A1(new_n458), .A2(G2106), .B1(G567), .B2(new_n459), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT68), .Z(G319));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(G137), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G101), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g041(.A(G125), .B1(new_n462), .B2(new_n463), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT69), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n469));
  OAI211_X1 g044(.A(new_n469), .B(G125), .C1(new_n462), .C2(new_n463), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n468), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n466), .B1(new_n472), .B2(G2105), .ZN(G160));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  OAI21_X1  g049(.A(G2104), .B1(new_n474), .B2(G112), .ZN(new_n475));
  INV_X1    g050(.A(G100), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n475), .B1(new_n476), .B2(new_n474), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT70), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n462), .A2(new_n463), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(new_n474), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n481));
  INV_X1    g056(.A(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  AOI21_X1  g059(.A(G2105), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI22_X1  g060(.A1(new_n480), .A2(G124), .B1(G136), .B2(new_n485), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n478), .A2(new_n486), .ZN(G162));
  NAND2_X1  g062(.A1(G126), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT72), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n474), .A2(G138), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n483), .A2(new_n484), .ZN(new_n493));
  OR2_X1    g068(.A1(KEYINPUT71), .A2(G114), .ZN(new_n494));
  NAND2_X1  g069(.A1(KEYINPUT71), .A2(G114), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n494), .A2(G2105), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n492), .A2(new_n493), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  OAI211_X1 g074(.A(G138), .B(new_n474), .C1(new_n462), .C2(new_n463), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT72), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n500), .A2(new_n490), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  NAND2_X1  g080(.A1(G50), .A2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT5), .B1(new_n507), .B2(KEYINPUT74), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT74), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n509), .A2(new_n510), .A3(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n506), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT73), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT73), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT6), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n515), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n516), .A2(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n514), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(G75), .A2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G62), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n524), .B1(new_n512), .B2(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n523), .A2(KEYINPUT75), .B1(G651), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT75), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n514), .A2(new_n522), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n527), .A2(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  AND2_X1   g106(.A1(new_n508), .A2(new_n511), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n532), .A2(G63), .A3(G651), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT76), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n534), .B1(new_n520), .B2(new_n521), .ZN(new_n535));
  INV_X1    g110(.A(new_n521), .ZN(new_n536));
  XNOR2_X1  g111(.A(KEYINPUT73), .B(KEYINPUT6), .ZN(new_n537));
  OAI211_X1 g112(.A(KEYINPUT76), .B(new_n536), .C1(new_n537), .C2(new_n515), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n535), .A2(G543), .A3(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G51), .ZN(new_n540));
  OAI211_X1 g115(.A(KEYINPUT77), .B(new_n533), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n522), .A2(G89), .A3(new_n532), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT78), .ZN(new_n543));
  NAND3_X1  g118(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT7), .ZN(new_n545));
  AND3_X1   g120(.A1(new_n542), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n543), .B1(new_n542), .B2(new_n545), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n541), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n536), .B1(new_n537), .B2(new_n515), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n507), .B1(new_n549), .B2(new_n534), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n550), .A2(G51), .A3(new_n538), .ZN(new_n551));
  AOI21_X1  g126(.A(KEYINPUT77), .B1(new_n551), .B2(new_n533), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n548), .A2(new_n552), .ZN(G168));
  AOI22_X1  g128(.A1(new_n532), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n554));
  OR2_X1    g129(.A1(new_n554), .A2(new_n515), .ZN(new_n555));
  XOR2_X1   g130(.A(KEYINPUT79), .B(G52), .Z(new_n556));
  NAND3_X1  g131(.A1(new_n550), .A2(new_n538), .A3(new_n556), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n549), .A2(new_n512), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G90), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n555), .A2(new_n557), .A3(new_n559), .ZN(G301));
  INV_X1    g135(.A(G301), .ZN(G171));
  NAND2_X1  g136(.A1(G68), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G56), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n512), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n558), .A2(G81), .B1(G651), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(G43), .ZN(new_n566));
  OAI211_X1 g141(.A(new_n565), .B(G860), .C1(new_n566), .C2(new_n539), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(G188));
  NAND4_X1  g146(.A1(new_n535), .A2(G53), .A3(G543), .A4(new_n538), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(KEYINPUT9), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n550), .A2(new_n574), .A3(G53), .A4(new_n538), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(G78), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G65), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n512), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n558), .A2(G91), .B1(G651), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n576), .A2(new_n580), .ZN(G299));
  INV_X1    g156(.A(G168), .ZN(G286));
  INV_X1    g157(.A(G74), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n515), .B1(new_n512), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n584), .B1(new_n558), .B2(G87), .ZN(new_n585));
  INV_X1    g160(.A(G49), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n586), .B2(new_n539), .ZN(G288));
  NAND3_X1  g162(.A1(new_n508), .A2(new_n511), .A3(G61), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(KEYINPUT80), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT80), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n508), .A2(new_n511), .A3(new_n590), .A4(G61), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT81), .ZN(new_n592));
  INV_X1    g167(.A(G73), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n593), .B2(new_n507), .ZN(new_n594));
  NAND3_X1  g169(.A1(KEYINPUT81), .A2(G73), .A3(G543), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n589), .A2(new_n591), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G651), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT82), .ZN(new_n600));
  NAND2_X1  g175(.A1(G48), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G86), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n512), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n599), .A2(new_n600), .B1(new_n522), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n596), .B1(new_n588), .B2(KEYINPUT80), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n515), .B1(new_n605), .B2(new_n591), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(KEYINPUT82), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n604), .A2(new_n607), .ZN(G305));
  AND3_X1   g183(.A1(new_n535), .A2(G543), .A3(new_n538), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G47), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n532), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n611), .A2(new_n515), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n558), .A2(G85), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(G290));
  NAND2_X1  g189(.A1(G301), .A2(G868), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT83), .ZN(new_n616));
  INV_X1    g191(.A(new_n520), .ZN(new_n617));
  NAND4_X1  g192(.A1(new_n617), .A2(new_n532), .A3(G92), .A4(new_n536), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT10), .ZN(new_n619));
  NAND4_X1  g194(.A1(new_n535), .A2(G54), .A3(G543), .A4(new_n538), .ZN(new_n620));
  NAND2_X1  g195(.A1(G79), .A2(G543), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT84), .B(G66), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n512), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G651), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT85), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n620), .A2(KEYINPUT85), .A3(new_n624), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n619), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n616), .B1(G868), .B2(new_n629), .ZN(G284));
  OAI21_X1  g205(.A(new_n616), .B1(G868), .B2(new_n629), .ZN(G321));
  INV_X1    g206(.A(G868), .ZN(new_n632));
  NOR2_X1   g207(.A1(G286), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G299), .B(KEYINPUT86), .Z(new_n634));
  AOI21_X1  g209(.A(new_n633), .B1(new_n634), .B2(new_n632), .ZN(G297));
  AOI21_X1  g210(.A(new_n633), .B1(new_n634), .B2(new_n632), .ZN(G280));
  INV_X1    g211(.A(G559), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n629), .B1(new_n637), .B2(G860), .ZN(G148));
  NAND2_X1  g213(.A1(new_n629), .A2(new_n637), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(G868), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n565), .B1(new_n566), .B2(new_n539), .ZN(new_n641));
  AOI22_X1  g216(.A1(new_n640), .A2(KEYINPUT87), .B1(new_n632), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(KEYINPUT87), .B2(new_n640), .ZN(G323));
  XNOR2_X1  g218(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g219(.A1(new_n485), .A2(G2104), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT12), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT88), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT13), .Z(new_n648));
  INV_X1    g223(.A(G2100), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n480), .A2(G123), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n485), .A2(G135), .ZN(new_n653));
  NOR2_X1   g228(.A1(G99), .A2(G2105), .ZN(new_n654));
  OAI21_X1  g229(.A(G2104), .B1(new_n474), .B2(G111), .ZN(new_n655));
  OAI211_X1 g230(.A(new_n652), .B(new_n653), .C1(new_n654), .C2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(G2096), .Z(new_n657));
  NAND3_X1  g232(.A1(new_n650), .A2(new_n651), .A3(new_n657), .ZN(G156));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1341), .B(G1348), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2443), .B(G2446), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2427), .B(G2438), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2430), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT15), .B(G2435), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  AND3_X1   g244(.A1(new_n668), .A2(new_n669), .A3(KEYINPUT14), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n664), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n664), .A2(new_n670), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n671), .A2(G14), .A3(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT89), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(G401));
  XOR2_X1   g251(.A(G2084), .B(G2090), .Z(new_n677));
  XNOR2_X1  g252(.A(G2067), .B(G2678), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n677), .ZN(new_n680));
  XOR2_X1   g255(.A(G2072), .B(G2078), .Z(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(KEYINPUT17), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n677), .A2(new_n678), .ZN(new_n684));
  OAI221_X1 g259(.A(new_n679), .B1(new_n678), .B2(new_n682), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n679), .A2(new_n681), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT18), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G2096), .B(G2100), .Z(new_n689));
  XOR2_X1   g264(.A(new_n688), .B(new_n689), .Z(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT90), .B(KEYINPUT91), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(G227));
  XNOR2_X1  g268(.A(G1971), .B(G1976), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT19), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(G1956), .B(G2474), .Z(new_n697));
  XOR2_X1   g272(.A(G1961), .B(G1966), .Z(new_n698));
  AND2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT20), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n697), .A2(new_n698), .ZN(new_n702));
  NOR3_X1   g277(.A1(new_n696), .A2(new_n699), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n696), .B2(new_n702), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G1986), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(G1991), .B(G1996), .ZN(new_n712));
  INV_X1    g287(.A(G1981), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n709), .A2(new_n714), .A3(new_n710), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(G229));
  INV_X1    g294(.A(KEYINPUT93), .ZN(new_n720));
  NOR2_X1   g295(.A1(G288), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n609), .A2(G49), .ZN(new_n722));
  AOI21_X1  g297(.A(KEYINPUT93), .B1(new_n722), .B2(new_n585), .ZN(new_n723));
  OAI21_X1  g298(.A(G16), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G16), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G23), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT33), .B(G1976), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n725), .A2(G22), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G166), .B2(new_n725), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G1971), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n599), .A2(new_n600), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n603), .A2(new_n522), .ZN(new_n736));
  AND3_X1   g311(.A1(new_n735), .A2(new_n607), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G16), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G6), .B2(G16), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT32), .B(G1981), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n727), .A2(new_n729), .B1(new_n739), .B2(new_n741), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n734), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(KEYINPUT34), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT34), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n734), .A2(new_n746), .A3(new_n742), .A4(new_n743), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n480), .A2(G119), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n485), .A2(G131), .ZN(new_n749));
  OR2_X1    g324(.A1(G95), .A2(G2105), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n750), .B(G2104), .C1(G107), .C2(new_n474), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n748), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT92), .Z(new_n753));
  MUX2_X1   g328(.A(G25), .B(new_n753), .S(G29), .Z(new_n754));
  XOR2_X1   g329(.A(KEYINPUT35), .B(G1991), .Z(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n754), .B(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(G290), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(G16), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G16), .B2(G24), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n760), .A2(new_n706), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n760), .A2(new_n706), .ZN(new_n762));
  NOR3_X1   g337(.A1(new_n757), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n745), .A2(new_n747), .A3(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT36), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(G29), .ZN(new_n767));
  NOR2_X1   g342(.A1(G162), .A2(new_n767), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n767), .A2(G35), .ZN(new_n769));
  OR3_X1    g344(.A1(new_n768), .A2(KEYINPUT101), .A3(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(KEYINPUT101), .B1(new_n768), .B2(new_n769), .ZN(new_n771));
  AND3_X1   g346(.A1(new_n770), .A2(KEYINPUT29), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(KEYINPUT29), .B1(new_n770), .B2(new_n771), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(G2090), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n480), .A2(G129), .ZN(new_n776));
  NAND3_X1  g351(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT26), .Z(new_n778));
  NAND3_X1  g353(.A1(new_n474), .A2(G105), .A3(G2104), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n485), .A2(G141), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n776), .A2(new_n778), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  AND3_X1   g357(.A1(new_n782), .A2(KEYINPUT99), .A3(G29), .ZN(new_n783));
  AOI21_X1  g358(.A(KEYINPUT99), .B1(new_n782), .B2(G29), .ZN(new_n784));
  OAI22_X1  g359(.A1(new_n783), .A2(new_n784), .B1(G29), .B2(G32), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT27), .B(G1996), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(KEYINPUT100), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(KEYINPUT100), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n774), .A2(new_n775), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(G29), .A2(G33), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT98), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n485), .A2(G139), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT25), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n493), .A2(G127), .ZN(new_n796));
  NAND2_X1  g371(.A1(G115), .A2(G2104), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n793), .B(new_n795), .C1(new_n798), .C2(new_n474), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n792), .B1(new_n799), .B2(new_n767), .ZN(new_n800));
  INV_X1    g375(.A(G2072), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n767), .A2(G27), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G164), .B2(new_n767), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n805), .A2(G2078), .ZN(new_n806));
  NOR3_X1   g381(.A1(new_n802), .A2(new_n803), .A3(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(G28), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n808), .A2(KEYINPUT30), .ZN(new_n809));
  AOI21_X1  g384(.A(G29), .B1(new_n808), .B2(KEYINPUT30), .ZN(new_n810));
  OR2_X1    g385(.A1(KEYINPUT31), .A2(G11), .ZN(new_n811));
  NAND2_X1  g386(.A1(KEYINPUT31), .A2(G11), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n809), .A2(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n656), .B2(new_n767), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n805), .B2(G2078), .ZN(new_n815));
  NAND2_X1  g390(.A1(G301), .A2(G16), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n725), .A2(G5), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n807), .B(new_n815), .C1(G1961), .C2(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(G1961), .B2(new_n819), .ZN(new_n821));
  AND2_X1   g396(.A1(KEYINPUT24), .A2(G34), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n767), .B1(KEYINPUT24), .B2(G34), .ZN(new_n823));
  OAI22_X1  g398(.A1(G160), .A2(new_n767), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n824), .A2(G2084), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(G2084), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n825), .B(new_n826), .C1(new_n785), .C2(new_n786), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n772), .A2(new_n773), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n827), .B1(new_n828), .B2(G2090), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n790), .A2(new_n821), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n725), .A2(G21), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(G168), .B2(new_n725), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n832), .A2(G1966), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(G1966), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n725), .A2(G20), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT23), .Z(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(G299), .B2(G16), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(G1956), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n833), .A2(new_n834), .A3(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n830), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n725), .A2(G4), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(new_n629), .B2(new_n725), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT94), .ZN(new_n843));
  INV_X1    g418(.A(G1348), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n725), .A2(G19), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(new_n641), .B2(G16), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n848), .A2(G1341), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n848), .A2(G1341), .ZN(new_n850));
  AOI22_X1  g425(.A1(new_n480), .A2(G128), .B1(G140), .B2(new_n485), .ZN(new_n851));
  OAI21_X1  g426(.A(KEYINPUT95), .B1(G104), .B2(G2105), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  NOR3_X1   g428(.A1(KEYINPUT95), .A2(G104), .A3(G2105), .ZN(new_n854));
  OAI221_X1 g429(.A(G2104), .B1(G116), .B2(new_n474), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(G29), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n767), .A2(G26), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT28), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(KEYINPUT96), .B(G2067), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  NOR3_X1   g437(.A1(new_n849), .A2(new_n850), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n845), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT97), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n845), .A2(KEYINPUT97), .A3(new_n863), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n840), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n766), .A2(new_n868), .ZN(G311));
  OR2_X1    g444(.A1(new_n766), .A2(new_n868), .ZN(G150));
  NAND2_X1  g445(.A1(G80), .A2(G543), .ZN(new_n871));
  INV_X1    g446(.A(G67), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n871), .B1(new_n512), .B2(new_n872), .ZN(new_n873));
  AOI22_X1  g448(.A1(new_n558), .A2(G93), .B1(G651), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n550), .A2(G55), .A3(new_n538), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n641), .B(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT38), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n629), .A2(G559), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT39), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n882), .B(KEYINPUT102), .Z(new_n883));
  AOI21_X1  g458(.A(G860), .B1(new_n880), .B2(new_n881), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n876), .A2(G860), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n886), .B(KEYINPUT37), .Z(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(G145));
  XNOR2_X1  g463(.A(new_n856), .B(new_n504), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(new_n781), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n890), .A2(new_n799), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n799), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT105), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n485), .A2(G142), .ZN(new_n897));
  NOR2_X1   g472(.A1(G106), .A2(G2105), .ZN(new_n898));
  OAI21_X1  g473(.A(G2104), .B1(new_n474), .B2(G118), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n480), .A2(G130), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n900), .A2(KEYINPUT103), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n900), .A2(KEYINPUT103), .ZN(new_n902));
  OAI221_X1 g477(.A(new_n897), .B1(new_n898), .B2(new_n899), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT104), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n646), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(KEYINPUT104), .ZN(new_n906));
  INV_X1    g481(.A(new_n646), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n903), .A2(KEYINPUT104), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n752), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n905), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n910), .B1(new_n905), .B2(new_n909), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n895), .B1(new_n891), .B2(new_n892), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n896), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  XOR2_X1   g492(.A(G160), .B(new_n656), .Z(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(G162), .ZN(new_n919));
  INV_X1    g494(.A(new_n913), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n911), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n919), .B1(new_n921), .B2(new_n915), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n917), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n894), .B1(new_n921), .B2(KEYINPUT106), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n914), .A2(new_n925), .A3(new_n893), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n924), .A2(new_n926), .A3(new_n919), .ZN(new_n927));
  INV_X1    g502(.A(G37), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n923), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g505(.A1(new_n876), .A2(new_n632), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n758), .B1(new_n721), .B2(new_n723), .ZN(new_n932));
  NAND2_X1  g507(.A1(G288), .A2(new_n720), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n722), .A2(KEYINPUT93), .A3(new_n585), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n933), .A2(G290), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(G305), .A2(G166), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n737), .A2(G303), .ZN(new_n937));
  AND4_X1   g512(.A1(new_n932), .A2(new_n935), .A3(new_n936), .A4(new_n937), .ZN(new_n938));
  AOI22_X1  g513(.A1(new_n932), .A2(new_n935), .B1(new_n937), .B2(new_n936), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n941));
  OR2_X1    g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n641), .A2(new_n876), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n641), .A2(new_n876), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(new_n639), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT41), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT10), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n618), .B(new_n950), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n620), .A2(KEYINPUT85), .A3(new_n624), .ZN(new_n952));
  AOI21_X1  g527(.A(KEYINPUT85), .B1(new_n620), .B2(new_n624), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n954), .B1(new_n576), .B2(new_n580), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n629), .A2(G299), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n949), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n954), .B(G299), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT41), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n948), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n958), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n960), .B1(new_n961), .B2(new_n948), .ZN(new_n962));
  OR3_X1    g537(.A1(new_n944), .A2(new_n962), .A3(KEYINPUT108), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT108), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n942), .A2(new_n964), .A3(new_n943), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n964), .B1(new_n942), .B2(new_n943), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n965), .B1(new_n966), .B2(new_n962), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n963), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n931), .B1(new_n968), .B2(new_n632), .ZN(G295));
  OAI21_X1  g544(.A(new_n931), .B1(new_n968), .B2(new_n632), .ZN(G331));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT110), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n959), .A2(new_n972), .A3(new_n957), .ZN(new_n973));
  OR2_X1    g548(.A1(new_n546), .A2(new_n547), .ZN(new_n974));
  INV_X1    g549(.A(new_n552), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n974), .A2(new_n975), .A3(G171), .A4(new_n541), .ZN(new_n976));
  OAI21_X1  g551(.A(G301), .B1(new_n548), .B2(new_n552), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n978), .A2(new_n877), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n947), .B1(new_n977), .B2(new_n976), .ZN(new_n980));
  OAI22_X1  g555(.A1(new_n979), .A2(new_n980), .B1(new_n957), .B2(new_n972), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n973), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n978), .A2(new_n877), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT109), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n947), .A2(new_n976), .A3(new_n977), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n947), .A2(KEYINPUT109), .A3(new_n976), .A4(new_n977), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n958), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n940), .B1(new_n982), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT43), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n979), .A2(new_n980), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n940), .B1(new_n991), .B2(new_n961), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n959), .A2(new_n957), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n993), .A2(new_n986), .A3(new_n987), .ZN(new_n994));
  AOI21_X1  g569(.A(G37), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  AND3_X1   g570(.A1(new_n989), .A2(new_n990), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n991), .A2(new_n961), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n940), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n990), .B1(new_n999), .B2(new_n995), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n971), .B1(new_n996), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n999), .A2(new_n995), .A3(new_n990), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n990), .B1(new_n989), .B2(new_n995), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT111), .ZN(new_n1004));
  OAI211_X1 g579(.A(KEYINPUT44), .B(new_n1002), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  AND2_X1   g580(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1001), .B1(new_n1005), .B2(new_n1006), .ZN(G397));
  NAND3_X1  g582(.A1(new_n933), .A2(G1976), .A3(new_n934), .ZN(new_n1008));
  NAND2_X1  g583(.A1(G160), .A2(G40), .ZN(new_n1009));
  INV_X1    g584(.A(G1384), .ZN(new_n1010));
  OR2_X1    g585(.A1(G102), .A2(G2105), .ZN(new_n1011));
  OAI21_X1  g586(.A(G2105), .B1(KEYINPUT71), .B2(G114), .ZN(new_n1012));
  AND2_X1   g587(.A1(KEYINPUT71), .A2(G114), .ZN(new_n1013));
  OAI211_X1 g588(.A(G2104), .B(new_n1011), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n488), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n501), .A2(KEYINPUT72), .ZN(new_n1016));
  INV_X1    g591(.A(G138), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1017), .A2(G2105), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1015), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1014), .B1(new_n1019), .B2(new_n479), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n490), .A2(new_n502), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1021), .B1(new_n485), .B2(G138), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1010), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1009), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G8), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G1976), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT52), .B1(G288), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1008), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n1008), .A2(new_n1026), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1029), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT49), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n713), .B1(new_n604), .B2(new_n607), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n735), .A2(new_n607), .A3(new_n713), .A4(new_n736), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT118), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n604), .A2(new_n1037), .A3(new_n713), .A4(new_n607), .ZN(new_n1038));
  AOI211_X1 g613(.A(new_n1033), .B(new_n1034), .C1(new_n1036), .C2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1034), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT49), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1032), .B1(new_n1043), .B2(new_n1026), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1045), .B1(G303), .B2(G8), .ZN(new_n1046));
  AOI211_X1 g621(.A(KEYINPUT55), .B(new_n1025), .C1(new_n527), .C2(new_n529), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(G1384), .B1(new_n499), .B2(new_n503), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n1050));
  OR2_X1    g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G40), .ZN(new_n1052));
  AOI211_X1 g627(.A(new_n1052), .B(new_n466), .C1(new_n472), .C2(G2105), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT50), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1049), .A2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1051), .A2(new_n775), .A3(new_n1053), .A4(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT45), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1023), .A2(new_n1057), .ZN(new_n1058));
  OAI211_X1 g633(.A(KEYINPUT45), .B(new_n1010), .C1(new_n1020), .C2(new_n1022), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1058), .A2(KEYINPUT115), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1023), .A2(new_n1061), .A3(new_n1057), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1009), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1056), .B1(new_n1063), .B2(G1971), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1048), .B1(new_n1064), .B2(G8), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1066));
  AOI21_X1  g641(.A(G1971), .B1(new_n1066), .B2(new_n1053), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1010), .B(new_n1050), .C1(new_n1020), .C2(new_n1022), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1053), .B(new_n1068), .C1(new_n1054), .C2(new_n1049), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1069), .A2(G2090), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1048), .B(G8), .C1(new_n1067), .C2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT117), .ZN(new_n1072));
  OAI22_X1  g647(.A1(new_n1063), .A2(G1971), .B1(G2090), .B2(new_n1069), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1073), .A2(new_n1074), .A3(G8), .A4(new_n1048), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1065), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G1966), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1059), .A2(KEYINPUT119), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n504), .A2(new_n1079), .A3(KEYINPUT45), .A4(new_n1010), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1053), .A2(new_n1058), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1077), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1068), .B1(new_n1049), .B2(new_n1054), .ZN(new_n1084));
  OR3_X1    g659(.A1(new_n1084), .A2(new_n1009), .A3(G2084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1086), .A2(G8), .A3(G168), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1044), .A2(new_n1076), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT63), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1072), .A2(new_n1075), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1059), .A2(KEYINPUT115), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT45), .B1(new_n504), .B2(new_n1010), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1062), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1053), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(G1971), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1084), .A2(new_n1009), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1097), .A2(new_n1098), .B1(new_n775), .B2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT120), .B1(new_n1100), .B2(new_n1025), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1048), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT120), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1073), .A2(new_n1103), .A3(G8), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1101), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1087), .A2(KEYINPUT63), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1092), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n1033), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1040), .A2(KEYINPUT49), .A3(new_n1041), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1109), .A2(new_n1026), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1032), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1091), .B1(new_n1107), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1087), .A2(KEYINPUT63), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1115), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1116), .A2(KEYINPUT121), .A3(new_n1044), .A4(new_n1105), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1090), .A2(new_n1114), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT54), .ZN(new_n1119));
  INV_X1    g694(.A(G2078), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1120), .B(new_n1053), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1082), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1122), .A2(G2078), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1059), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(G1961), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1124), .A2(new_n1126), .B1(new_n1069), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1123), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1119), .B1(new_n1129), .B2(G171), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1131), .A2(new_n1125), .B1(new_n1069), .B2(new_n1127), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1123), .A2(new_n1132), .A3(G301), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT126), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1123), .A2(new_n1132), .A3(KEYINPUT126), .A4(G301), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1130), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT51), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1083), .A2(G168), .A3(new_n1085), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1138), .B1(new_n1139), .B2(G8), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1139), .A2(G8), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1138), .B1(new_n1086), .B2(G286), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1141), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AND4_X1   g719(.A1(new_n1044), .A2(new_n1137), .A3(new_n1076), .A4(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n844), .B1(new_n1084), .B2(new_n1009), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT122), .ZN(new_n1147));
  INV_X1    g722(.A(G2067), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1053), .A2(new_n1147), .A3(new_n1148), .A4(new_n1049), .ZN(new_n1149));
  NAND4_X1  g724(.A1(G160), .A2(new_n1049), .A3(G40), .A4(new_n1148), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(KEYINPUT122), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1146), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT123), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1152), .A2(new_n1153), .A3(new_n629), .ZN(new_n1154));
  XNOR2_X1  g729(.A(KEYINPUT56), .B(G2072), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1053), .B(new_n1155), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1051), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1157));
  INV_X1    g732(.A(G1956), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT57), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n576), .A2(new_n1161), .A3(new_n580), .ZN(new_n1162));
  AOI22_X1  g737(.A1(new_n1156), .A2(new_n1159), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1153), .B1(new_n1152), .B2(new_n629), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1154), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1156), .A2(new_n1159), .A3(new_n1160), .A4(new_n1162), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(KEYINPUT124), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT124), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1164), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1170), .A2(new_n1173), .ZN(new_n1174));
  OAI211_X1 g749(.A(new_n1169), .B(new_n1166), .C1(new_n1174), .C2(new_n1154), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1176), .B1(new_n1167), .B2(new_n1163), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1173), .A2(KEYINPUT61), .A3(new_n1166), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT60), .ZN(new_n1179));
  OR2_X1    g754(.A1(new_n1152), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1152), .A2(new_n1179), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1180), .A2(new_n629), .A3(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1177), .A2(new_n1178), .A3(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g758(.A(KEYINPUT58), .B(G1341), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1024), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(G1996), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1185), .B1(new_n1186), .B2(new_n1063), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT59), .ZN(new_n1188));
  OR3_X1    g763(.A1(new_n1187), .A2(new_n1188), .A3(new_n641), .ZN(new_n1189));
  OR3_X1    g764(.A1(new_n1152), .A2(new_n1179), .A3(new_n629), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1188), .B1(new_n1187), .B2(new_n641), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  OAI211_X1 g767(.A(new_n1168), .B(new_n1175), .C1(new_n1183), .C2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1123), .A2(new_n1132), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1194), .A2(G171), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1195), .A2(KEYINPUT125), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT125), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1194), .A2(new_n1197), .A3(G171), .ZN(new_n1198));
  OAI211_X1 g773(.A(new_n1196), .B(new_n1198), .C1(G171), .C2(new_n1129), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(new_n1119), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1145), .A2(new_n1193), .A3(new_n1200), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n722), .A2(new_n1027), .A3(new_n585), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1202), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1203));
  INV_X1    g778(.A(new_n1040), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1026), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND4_X1  g780(.A1(new_n1111), .A2(new_n1112), .A3(new_n1072), .A4(new_n1075), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT62), .ZN(new_n1208));
  NOR2_X1   g783(.A1(new_n1143), .A2(new_n1142), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1208), .B1(new_n1209), .B2(new_n1140), .ZN(new_n1210));
  OAI211_X1 g785(.A(new_n1141), .B(KEYINPUT62), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1211));
  AOI22_X1  g786(.A1(new_n1210), .A2(new_n1211), .B1(new_n1198), .B2(new_n1196), .ZN(new_n1212));
  AND2_X1   g787(.A1(new_n1044), .A2(new_n1076), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1207), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g789(.A1(new_n1118), .A2(new_n1201), .A3(new_n1214), .ZN(new_n1215));
  NOR2_X1   g790(.A1(new_n1009), .A2(new_n1058), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n758), .A2(new_n706), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n1216), .B1(new_n1217), .B2(KEYINPUT112), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1218), .B1(KEYINPUT112), .B2(new_n1217), .ZN(new_n1219));
  INV_X1    g794(.A(new_n1216), .ZN(new_n1220));
  NOR3_X1   g795(.A1(new_n1220), .A2(new_n758), .A3(new_n706), .ZN(new_n1221));
  NOR2_X1   g796(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1222));
  XNOR2_X1  g797(.A(new_n1222), .B(KEYINPUT113), .ZN(new_n1223));
  NAND3_X1  g798(.A1(new_n1216), .A2(new_n1186), .A3(new_n782), .ZN(new_n1224));
  XNOR2_X1  g799(.A(new_n1224), .B(KEYINPUT114), .ZN(new_n1225));
  XNOR2_X1  g800(.A(new_n856), .B(new_n1148), .ZN(new_n1226));
  OAI21_X1  g801(.A(new_n1226), .B1(new_n1186), .B2(new_n782), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1227), .A2(new_n1216), .ZN(new_n1228));
  XNOR2_X1  g803(.A(new_n752), .B(new_n755), .ZN(new_n1229));
  OAI211_X1 g804(.A(new_n1225), .B(new_n1228), .C1(new_n1220), .C2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g805(.A1(new_n1223), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n1215), .A2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g807(.A(new_n1220), .B1(new_n1226), .B2(new_n782), .ZN(new_n1233));
  INV_X1    g808(.A(KEYINPUT46), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1216), .A2(new_n1186), .ZN(new_n1235));
  AOI21_X1  g810(.A(new_n1233), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g811(.A(new_n1236), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1237));
  XNOR2_X1  g812(.A(new_n1237), .B(KEYINPUT47), .ZN(new_n1238));
  XNOR2_X1  g813(.A(new_n1219), .B(KEYINPUT48), .ZN(new_n1239));
  OAI21_X1  g814(.A(new_n1238), .B1(new_n1230), .B2(new_n1239), .ZN(new_n1240));
  NOR2_X1   g815(.A1(new_n753), .A2(new_n756), .ZN(new_n1241));
  NAND3_X1  g816(.A1(new_n1225), .A2(new_n1228), .A3(new_n1241), .ZN(new_n1242));
  NAND3_X1  g817(.A1(new_n851), .A2(new_n1148), .A3(new_n855), .ZN(new_n1243));
  AOI21_X1  g818(.A(new_n1220), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NOR2_X1   g819(.A1(new_n1240), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g820(.A1(new_n1232), .A2(new_n1245), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g821(.A1(new_n673), .A2(new_n674), .ZN(new_n1248));
  NOR2_X1   g822(.A1(new_n673), .A2(new_n674), .ZN(new_n1249));
  OAI211_X1 g823(.A(G319), .B(new_n692), .C1(new_n1248), .C2(new_n1249), .ZN(new_n1250));
  INV_X1    g824(.A(KEYINPUT127), .ZN(new_n1251));
  NAND2_X1  g825(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g826(.A1(new_n1252), .A2(new_n718), .ZN(new_n1253));
  NOR2_X1   g827(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1254));
  NOR2_X1   g828(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  OAI211_X1 g829(.A(new_n1255), .B(new_n929), .C1(new_n1000), .C2(new_n996), .ZN(G225));
  INV_X1    g830(.A(G225), .ZN(G308));
endmodule


