//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n541, new_n542, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n596, new_n597, new_n600, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1145, new_n1146, new_n1147, new_n1148;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT67), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT68), .Z(new_n460));
  AOI21_X1  g035(.A(new_n460), .B1(new_n453), .B2(G2106), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(KEYINPUT69), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(G125), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n462), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT70), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(new_n465), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT70), .A2(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n476), .A2(KEYINPUT3), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT71), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g055(.A1(new_n476), .A2(KEYINPUT71), .A3(KEYINPUT3), .A4(new_n477), .ZN(new_n481));
  NAND4_X1  g056(.A1(new_n480), .A2(G137), .A3(new_n464), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n476), .A2(new_n477), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G101), .ZN(new_n484));
  AOI21_X1  g059(.A(G2105), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n474), .A2(new_n485), .ZN(G160));
  NAND3_X1  g061(.A1(new_n480), .A2(new_n464), .A3(new_n481), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(new_n462), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  XOR2_X1   g064(.A(new_n489), .B(KEYINPUT72), .Z(new_n490));
  OR2_X1    g065(.A1(G100), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n487), .A2(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G136), .ZN(new_n494));
  AND3_X1   g069(.A1(new_n490), .A2(new_n492), .A3(new_n494), .ZN(G162));
  AND2_X1   g070(.A1(KEYINPUT4), .A2(G138), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n480), .A2(new_n464), .A3(new_n481), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(G102), .A2(G2104), .ZN(new_n498));
  AOI21_X1  g073(.A(G2105), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n480), .A2(G126), .A3(new_n464), .A4(new_n481), .ZN(new_n500));
  NAND2_X1  g075(.A1(G114), .A2(G2104), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n462), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n467), .A2(KEYINPUT69), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n469), .A2(new_n470), .ZN(new_n504));
  AOI21_X1  g079(.A(G2105), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g080(.A(KEYINPUT4), .B1(new_n505), .B2(G138), .ZN(new_n506));
  NOR3_X1   g081(.A1(new_n499), .A2(new_n502), .A3(new_n506), .ZN(G164));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n508), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n514), .A2(new_n517), .ZN(G166));
  NAND3_X1  g093(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n519));
  INV_X1    g094(.A(G89), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n519), .B1(new_n510), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  INV_X1    g098(.A(G51), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n512), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n521), .A2(new_n525), .ZN(G168));
  INV_X1    g101(.A(G90), .ZN(new_n527));
  INV_X1    g102(.A(G52), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n510), .A2(new_n527), .B1(new_n512), .B2(new_n528), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n516), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n529), .A2(new_n531), .ZN(G171));
  INV_X1    g107(.A(G81), .ZN(new_n533));
  INV_X1    g108(.A(G43), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n510), .A2(new_n533), .B1(new_n512), .B2(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n516), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G860), .ZN(G153));
  NAND4_X1  g114(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g115(.A1(G1), .A2(G3), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT8), .ZN(new_n542));
  NAND4_X1  g117(.A1(G319), .A2(G483), .A3(G661), .A4(new_n542), .ZN(G188));
  AND2_X1   g118(.A1(new_n509), .A2(G65), .ZN(new_n544));
  AND2_X1   g119(.A1(G78), .A2(G543), .ZN(new_n545));
  OAI21_X1  g120(.A(G651), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(G91), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT73), .ZN(new_n548));
  INV_X1    g123(.A(G53), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n512), .B2(new_n549), .ZN(new_n550));
  OAI221_X1 g125(.A(new_n546), .B1(new_n547), .B2(new_n510), .C1(KEYINPUT9), .C2(new_n550), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n508), .A2(KEYINPUT73), .A3(G53), .A4(G543), .ZN(new_n552));
  AND3_X1   g127(.A1(new_n550), .A2(KEYINPUT9), .A3(new_n552), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n551), .A2(new_n553), .ZN(G299));
  INV_X1    g129(.A(G171), .ZN(G301));
  INV_X1    g130(.A(G168), .ZN(G286));
  INV_X1    g131(.A(G166), .ZN(G303));
  OAI21_X1  g132(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(KEYINPUT74), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n560));
  OAI211_X1 g135(.A(new_n560), .B(G651), .C1(new_n509), .C2(G74), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n508), .A2(G49), .A3(G543), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n509), .A2(new_n508), .A3(G87), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n559), .A2(new_n561), .A3(new_n562), .A4(new_n563), .ZN(G288));
  INV_X1    g139(.A(G86), .ZN(new_n565));
  INV_X1    g140(.A(G48), .ZN(new_n566));
  OAI22_X1  g141(.A1(new_n510), .A2(new_n565), .B1(new_n512), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n509), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n568), .A2(new_n516), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT75), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(G305));
  INV_X1    g147(.A(G85), .ZN(new_n573));
  INV_X1    g148(.A(G47), .ZN(new_n574));
  OAI22_X1  g149(.A1(new_n510), .A2(new_n573), .B1(new_n512), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n576), .A2(new_n516), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G290));
  INV_X1    g154(.A(G868), .ZN(new_n580));
  NOR2_X1   g155(.A1(G301), .A2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n509), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G54), .ZN(new_n583));
  OAI22_X1  g158(.A1(new_n582), .A2(new_n516), .B1(new_n512), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT76), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n584), .B(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n509), .A2(new_n508), .A3(G92), .ZN(new_n587));
  XOR2_X1   g162(.A(new_n587), .B(KEYINPUT10), .Z(new_n588));
  AND2_X1   g163(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n589), .A2(KEYINPUT77), .ZN(new_n590));
  AND3_X1   g165(.A1(new_n586), .A2(KEYINPUT77), .A3(new_n588), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n581), .B1(new_n592), .B2(new_n580), .ZN(G284));
  AOI21_X1  g168(.A(new_n581), .B1(new_n592), .B2(new_n580), .ZN(G321));
  NAND2_X1  g169(.A1(G286), .A2(G868), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT78), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n551), .A2(new_n553), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(G868), .B2(new_n597), .ZN(G297));
  OAI21_X1  g173(.A(new_n596), .B1(G868), .B2(new_n597), .ZN(G280));
  XNOR2_X1  g174(.A(KEYINPUT79), .B(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n592), .B1(G860), .B2(new_n600), .ZN(G148));
  NAND2_X1  g176(.A1(new_n592), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n538), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g180(.A1(new_n505), .A2(new_n483), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT12), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT13), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(G2100), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n493), .A2(G135), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n488), .A2(G123), .ZN(new_n611));
  NOR2_X1   g186(.A1(G99), .A2(G2105), .ZN(new_n612));
  OAI21_X1  g187(.A(G2104), .B1(new_n462), .B2(G111), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n610), .B(new_n611), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(G2096), .Z(new_n615));
  NAND2_X1  g190(.A1(new_n609), .A2(new_n615), .ZN(G156));
  XOR2_X1   g191(.A(G2451), .B(G2454), .Z(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT16), .ZN(new_n618));
  XNOR2_X1  g193(.A(G1341), .B(G1348), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(G2443), .B(G2446), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(G2427), .B(G2438), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2430), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT15), .B(G2435), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n626), .A2(new_n627), .A3(KEYINPUT14), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n622), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n622), .A2(new_n629), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n630), .A2(new_n631), .A3(G14), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(G401));
  XNOR2_X1  g208(.A(G2067), .B(G2678), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT80), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT81), .ZN(new_n636));
  XOR2_X1   g211(.A(G2072), .B(G2078), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2084), .B(G2090), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n637), .B(KEYINPUT17), .ZN(new_n640));
  OAI211_X1 g215(.A(new_n638), .B(new_n639), .C1(new_n636), .C2(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT82), .Z(new_n642));
  NOR3_X1   g217(.A1(new_n635), .A2(new_n637), .A3(new_n639), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT18), .Z(new_n644));
  INV_X1    g219(.A(new_n640), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n645), .A2(new_n639), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n644), .B1(new_n636), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2096), .B(G2100), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT83), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n648), .B(new_n650), .ZN(G227));
  XNOR2_X1  g226(.A(G1971), .B(G1976), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT19), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1956), .B(G2474), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1961), .B(G1966), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT20), .Z(new_n659));
  NAND2_X1  g234(.A1(new_n654), .A2(new_n655), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT84), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(new_n653), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n659), .B(new_n663), .C1(new_n653), .C2(new_n660), .ZN(new_n664));
  INV_X1    g239(.A(G1986), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1991), .B(G1996), .ZN(new_n669));
  INV_X1    g244(.A(G1981), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n668), .B(new_n671), .Z(G229));
  INV_X1    g247(.A(G16), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(G22), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n674), .B1(G166), .B2(new_n673), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n675), .A2(G1971), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(G1971), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n673), .A2(G23), .ZN(new_n678));
  INV_X1    g253(.A(G288), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n678), .B1(new_n679), .B2(new_n673), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT33), .B(G1976), .Z(new_n681));
  OAI211_X1 g256(.A(new_n676), .B(new_n677), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(G6), .A2(G16), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(new_n571), .B2(G16), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT32), .B(G1981), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  AOI211_X1 g261(.A(new_n682), .B(new_n686), .C1(new_n680), .C2(new_n681), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT34), .ZN(new_n688));
  NOR2_X1   g263(.A1(G25), .A2(G29), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n493), .A2(G131), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n488), .A2(G119), .ZN(new_n691));
  OR2_X1    g266(.A1(G95), .A2(G2105), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n692), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n690), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n689), .B1(new_n695), .B2(G29), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT35), .B(G1991), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT85), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n696), .A2(new_n698), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n673), .A2(G24), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(new_n578), .B2(new_n673), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(new_n665), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT36), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n703), .B1(KEYINPUT86), .B2(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n700), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n688), .A2(new_n699), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n704), .A2(KEYINPUT86), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n707), .B(new_n708), .Z(new_n709));
  NAND2_X1  g284(.A1(new_n493), .A2(G141), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT91), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n488), .A2(G129), .ZN(new_n712));
  NAND3_X1  g287(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT26), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n483), .A2(G105), .A3(new_n462), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT92), .ZN(new_n716));
  NOR4_X1   g291(.A1(new_n711), .A2(new_n712), .A3(new_n714), .A4(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G29), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT93), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G29), .B2(G32), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT94), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT27), .B(G1996), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(G4), .A2(G16), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT87), .Z(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n592), .B2(G16), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G1348), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G35), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G162), .B2(new_n728), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT29), .B(G2090), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n727), .A2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G28), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n734), .A2(KEYINPUT30), .ZN(new_n735));
  AOI21_X1  g310(.A(G29), .B1(new_n734), .B2(KEYINPUT30), .ZN(new_n736));
  OR2_X1    g311(.A1(KEYINPUT31), .A2(G11), .ZN(new_n737));
  NAND2_X1  g312(.A1(KEYINPUT31), .A2(G11), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n735), .A2(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n614), .B2(new_n728), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT95), .Z(new_n741));
  NAND2_X1  g316(.A1(new_n728), .A2(G26), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT28), .Z(new_n743));
  NAND2_X1  g318(.A1(new_n493), .A2(G140), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n488), .A2(G128), .ZN(new_n745));
  NOR2_X1   g320(.A1(G104), .A2(G2105), .ZN(new_n746));
  OAI21_X1  g321(.A(G2104), .B1(new_n462), .B2(G116), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n744), .B(new_n745), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n743), .B1(new_n748), .B2(G29), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT89), .B(G2067), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(G164), .A2(G29), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G27), .B2(G29), .ZN(new_n753));
  INV_X1    g328(.A(G2078), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR3_X1   g330(.A1(new_n741), .A2(new_n751), .A3(new_n755), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n728), .A2(G33), .ZN(new_n757));
  INV_X1    g332(.A(G127), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n503), .B2(new_n504), .ZN(new_n759));
  AND2_X1   g334(.A1(G115), .A2(G2104), .ZN(new_n760));
  OAI21_X1  g335(.A(G2105), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT90), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n493), .A2(G139), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT25), .Z(new_n765));
  NAND3_X1  g340(.A1(new_n762), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n757), .B1(new_n766), .B2(G29), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G2084), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT24), .ZN(new_n770));
  INV_X1    g345(.A(G34), .ZN(new_n771));
  AOI21_X1  g346(.A(G29), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n770), .B2(new_n771), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G160), .B2(new_n728), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  OAI22_X1  g350(.A1(new_n768), .A2(G2072), .B1(new_n769), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G2072), .B2(new_n768), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n673), .A2(G20), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT23), .Z(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G299), .B2(G16), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1956), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n673), .A2(G5), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G171), .B2(new_n673), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1961), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n673), .A2(G19), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT88), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n538), .B2(new_n673), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G1341), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n673), .A2(G21), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G168), .B2(new_n673), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G1966), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n784), .A2(new_n788), .A3(new_n791), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n781), .B(new_n792), .C1(G2084), .C2(new_n774), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n754), .B2(new_n753), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n733), .A2(new_n756), .A3(new_n777), .A4(new_n794), .ZN(new_n795));
  NOR3_X1   g370(.A1(new_n709), .A2(new_n723), .A3(new_n795), .ZN(G311));
  OR3_X1    g371(.A1(new_n709), .A2(new_n723), .A3(new_n795), .ZN(G150));
  INV_X1    g372(.A(G93), .ZN(new_n798));
  INV_X1    g373(.A(G55), .ZN(new_n799));
  OAI22_X1  g374(.A1(new_n510), .A2(new_n798), .B1(new_n512), .B2(new_n799), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n801), .A2(new_n516), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(G860), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT97), .B(KEYINPUT37), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n592), .A2(G559), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n538), .B(new_n803), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n813), .A2(KEYINPUT39), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n804), .B1(new_n813), .B2(KEYINPUT39), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n807), .B1(new_n814), .B2(new_n815), .ZN(G145));
  NAND2_X1  g391(.A1(new_n497), .A2(new_n498), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(new_n462), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n500), .A2(new_n501), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(G2105), .ZN(new_n820));
  OAI211_X1 g395(.A(G138), .B(new_n462), .C1(new_n468), .C2(new_n471), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT4), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n818), .A2(new_n820), .A3(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n748), .B(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n717), .B(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(new_n766), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n493), .A2(G142), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n488), .A2(G130), .ZN(new_n829));
  NOR2_X1   g404(.A1(G106), .A2(G2105), .ZN(new_n830));
  OAI21_X1  g405(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n828), .B(new_n829), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(new_n607), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(new_n694), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(KEYINPUT98), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n827), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n827), .A2(new_n835), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n614), .B(G160), .ZN(new_n838));
  XNOR2_X1  g413(.A(G162), .B(new_n838), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT99), .Z(new_n840));
  NAND3_X1  g415(.A1(new_n836), .A2(new_n837), .A3(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(G37), .ZN(new_n842));
  INV_X1    g417(.A(new_n839), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n827), .B(new_n834), .ZN(new_n844));
  OAI211_X1 g419(.A(new_n841), .B(new_n842), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g421(.A(new_n571), .B(new_n679), .ZN(new_n847));
  XOR2_X1   g422(.A(G166), .B(new_n578), .Z(new_n848));
  OR2_X1    g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n848), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT102), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT42), .Z(new_n853));
  INV_X1    g428(.A(new_n811), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n602), .B(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT41), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n589), .A2(G299), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n586), .A2(new_n588), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n858), .A2(new_n597), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n856), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n857), .A2(new_n859), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(KEYINPUT41), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n855), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT101), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n855), .A2(new_n862), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT100), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n853), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n852), .B(KEYINPUT42), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n871), .A2(new_n868), .A3(new_n866), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n870), .A2(G868), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT103), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n870), .A2(new_n875), .A3(new_n872), .A4(G868), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n580), .B1(new_n800), .B2(new_n802), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n874), .A2(new_n876), .A3(new_n877), .ZN(G295));
  NAND3_X1  g453(.A1(new_n874), .A2(new_n876), .A3(new_n877), .ZN(G331));
  INV_X1    g454(.A(KEYINPUT44), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n849), .A2(new_n850), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT105), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n849), .A2(KEYINPUT105), .A3(new_n850), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n863), .A2(KEYINPUT106), .A3(new_n860), .ZN(new_n886));
  XNOR2_X1  g461(.A(G171), .B(G168), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n811), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT104), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n811), .A2(new_n887), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n889), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n860), .A2(KEYINPUT106), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n886), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT107), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n857), .A2(new_n859), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n888), .A2(new_n891), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  AOI22_X1  g474(.A1(new_n895), .A2(new_n896), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n886), .A2(new_n894), .A3(new_n893), .A4(KEYINPUT107), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n885), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n898), .B1(new_n864), .B2(new_n861), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n890), .A2(new_n897), .A3(new_n891), .A4(new_n892), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n842), .B1(new_n905), .B2(new_n881), .ZN(new_n906));
  OAI21_X1  g481(.A(KEYINPUT43), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT43), .ZN(new_n908));
  INV_X1    g483(.A(new_n885), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n906), .B1(new_n909), .B2(new_n905), .ZN(new_n910));
  AOI22_X1  g485(.A1(new_n907), .A2(KEYINPUT108), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT108), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n912), .B(KEYINPUT43), .C1(new_n902), .C2(new_n906), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n880), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n905), .A2(new_n881), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n915), .A2(G37), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n900), .A2(new_n901), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n908), .B(new_n916), .C1(new_n917), .C2(new_n885), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n918), .B(new_n880), .C1(new_n908), .C2(new_n910), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT109), .B1(new_n914), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n907), .A2(KEYINPUT108), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n910), .A2(new_n908), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n913), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT44), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT109), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n925), .A2(new_n926), .A3(new_n919), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n921), .A2(new_n927), .ZN(G397));
  INV_X1    g503(.A(G1384), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n824), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT45), .ZN(new_n931));
  INV_X1    g506(.A(G40), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n474), .A2(new_n485), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n934), .A2(G1996), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n717), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n936), .B(KEYINPUT110), .ZN(new_n937));
  XOR2_X1   g512(.A(new_n748), .B(G2067), .Z(new_n938));
  INV_X1    g513(.A(G1996), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n938), .B1(new_n717), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n934), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XOR2_X1   g517(.A(new_n694), .B(new_n698), .Z(new_n943));
  OAI211_X1 g518(.A(new_n937), .B(new_n942), .C1(new_n934), .C2(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n578), .B(new_n665), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n944), .B1(new_n941), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT121), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT111), .ZN(new_n948));
  NOR2_X1   g523(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n948), .B1(G164), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n824), .A2(KEYINPUT111), .A3(new_n949), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(G160), .A2(G40), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n954), .B1(new_n930), .B2(KEYINPUT50), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n953), .A2(new_n955), .A3(new_n769), .ZN(new_n956));
  INV_X1    g531(.A(G1966), .ZN(new_n957));
  AOI22_X1  g532(.A1(new_n819), .A2(G2105), .B1(new_n822), .B2(new_n821), .ZN(new_n958));
  AOI21_X1  g533(.A(G1384), .B1(new_n958), .B2(new_n818), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n933), .B1(new_n959), .B2(KEYINPUT45), .ZN(new_n960));
  NOR3_X1   g535(.A1(G164), .A2(new_n931), .A3(G1384), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n956), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(G286), .A2(G8), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT119), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n966), .B(KEYINPUT120), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n963), .A2(G8), .ZN(new_n968));
  INV_X1    g543(.A(new_n965), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(KEYINPUT51), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT51), .ZN(new_n971));
  INV_X1    g546(.A(G8), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n972), .B1(new_n956), .B2(new_n962), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n971), .B1(new_n973), .B2(new_n965), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n970), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n947), .B1(new_n967), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT120), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n966), .B(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n978), .A2(KEYINPUT121), .A3(new_n974), .A4(new_n970), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT62), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT53), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n954), .B1(new_n930), .B2(new_n931), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n959), .A2(KEYINPUT45), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n983), .A2(new_n754), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n953), .A2(new_n955), .ZN(new_n986));
  INV_X1    g561(.A(G1961), .ZN(new_n987));
  AOI22_X1  g562(.A1(new_n982), .A2(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n983), .A2(new_n984), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n754), .A2(KEYINPUT53), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n991), .A2(G171), .ZN(new_n992));
  INV_X1    g567(.A(G2090), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n953), .A2(new_n955), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G1971), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(new_n960), .B2(new_n961), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT112), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(G303), .A2(G8), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n1000), .B(KEYINPUT55), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n994), .A2(new_n996), .A3(KEYINPUT112), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n999), .A2(G8), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n959), .A2(new_n933), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n679), .A2(G1976), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(G8), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT52), .ZN(new_n1008));
  INV_X1    g583(.A(G1976), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT52), .B1(G288), .B2(new_n1009), .ZN(new_n1010));
  XOR2_X1   g585(.A(new_n1010), .B(KEYINPUT113), .Z(new_n1011));
  NAND4_X1  g586(.A1(new_n1011), .A2(G8), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n570), .A2(G1981), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT49), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n567), .A2(new_n569), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1015), .A2(new_n670), .ZN(new_n1016));
  OR3_X1    g591(.A1(new_n1013), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1014), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1017), .A2(new_n1005), .A3(G8), .A4(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1008), .A2(new_n1012), .A3(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(KEYINPUT114), .B1(G164), .B2(new_n950), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n824), .A2(new_n1022), .A3(new_n949), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT50), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n933), .B1(new_n959), .B2(new_n1025), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n1024), .A2(new_n1026), .A3(G2090), .ZN(new_n1027));
  AOI21_X1  g602(.A(G1971), .B1(new_n983), .B2(new_n984), .ZN(new_n1028));
  OAI21_X1  g603(.A(G8), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1020), .B1(new_n1029), .B2(new_n1001), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1004), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT62), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n976), .A2(new_n979), .A3(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n981), .A2(new_n992), .A3(new_n1032), .A4(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT57), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n597), .B(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g612(.A(KEYINPUT56), .B(G2072), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n983), .A2(new_n984), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G1956), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT117), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1044), .A2(new_n1021), .A3(new_n933), .A4(new_n1023), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT117), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1045), .A2(new_n1046), .A3(new_n1041), .ZN(new_n1047));
  AOI211_X1 g622(.A(new_n1037), .B(new_n1040), .C1(new_n1043), .C2(new_n1047), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1045), .A2(new_n1046), .A3(new_n1041), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1046), .B1(new_n1045), .B2(new_n1041), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1039), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n1037), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1005), .A2(G2067), .ZN(new_n1053));
  INV_X1    g628(.A(G1348), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1053), .B1(new_n986), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n592), .ZN(new_n1056));
  OR2_X1    g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1048), .B1(new_n1052), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1055), .A2(KEYINPUT60), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1059), .A2(new_n1056), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n592), .B1(new_n1055), .B2(KEYINPUT60), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1060), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT61), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1037), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1043), .A2(new_n1047), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1064), .B1(new_n1065), .B2(new_n1039), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1063), .B1(new_n1066), .B2(new_n1048), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1065), .A2(new_n1064), .A3(new_n1039), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1052), .A2(KEYINPUT61), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1005), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT58), .B(G1341), .ZN(new_n1071));
  OAI22_X1  g646(.A1(new_n989), .A2(G1996), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(new_n538), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n1073), .B(KEYINPUT59), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1067), .A2(new_n1069), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT118), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1062), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1067), .A2(KEYINPUT118), .A3(new_n1069), .A4(new_n1074), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1058), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n961), .A2(new_n990), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n983), .A2(KEYINPUT122), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n960), .A2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1080), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT123), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1087));
  OAI211_X1 g662(.A(G301), .B(new_n988), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT124), .ZN(new_n1089));
  XNOR2_X1  g664(.A(new_n1084), .B(new_n1085), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT124), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1090), .A2(new_n1091), .A3(G301), .A4(new_n988), .ZN(new_n1092));
  AOI21_X1  g667(.A(KEYINPUT54), .B1(new_n991), .B2(G171), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1089), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1090), .A2(G171), .A3(new_n988), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n991), .A2(G301), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1095), .A2(KEYINPUT54), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1098), .A2(new_n980), .A3(new_n1032), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1035), .B1(new_n1079), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n968), .A2(G286), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1004), .A2(new_n1030), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT63), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1103), .A2(KEYINPUT115), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT115), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1020), .A2(new_n1104), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1004), .A2(new_n1107), .A3(new_n1102), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n972), .B1(new_n997), .B2(new_n998), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1002), .B1(new_n1109), .B2(new_n1003), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  NOR3_X1   g686(.A1(new_n1105), .A2(new_n1106), .A3(new_n1111), .ZN(new_n1112));
  OR2_X1    g687(.A1(new_n1004), .A2(new_n1020), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n1019), .A2(new_n1009), .A3(new_n679), .ZN(new_n1114));
  OAI211_X1 g689(.A(G8), .B(new_n1005), .C1(new_n1114), .C2(new_n1013), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1101), .B1(new_n1112), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1116), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT115), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1111), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  OAI211_X1 g698(.A(KEYINPUT116), .B(new_n1118), .C1(new_n1123), .C2(new_n1105), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1117), .A2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n946), .B1(new_n1100), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n938), .A2(new_n717), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n941), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n935), .A2(KEYINPUT46), .ZN(new_n1129));
  AND2_X1   g704(.A1(new_n1129), .A2(KEYINPUT125), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT125), .B1(new_n935), .B2(KEYINPUT46), .ZN(new_n1131));
  OAI221_X1 g706(.A(new_n1128), .B1(KEYINPUT46), .B2(new_n935), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n1132), .B(KEYINPUT47), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n937), .A2(new_n942), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1134), .A2(new_n698), .A3(new_n694), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n748), .A2(G2067), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n941), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n934), .A2(G1986), .A3(G290), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1138), .B(KEYINPUT48), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1133), .B(new_n1137), .C1(new_n944), .C2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT126), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n1140), .B(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1126), .A2(new_n1142), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g718(.A1(new_n632), .A2(G319), .ZN(new_n1145));
  NOR3_X1   g719(.A1(G229), .A2(G227), .A3(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g720(.A(new_n1146), .B(KEYINPUT127), .ZN(new_n1147));
  OAI21_X1  g721(.A(new_n918), .B1(new_n908), .B2(new_n910), .ZN(new_n1148));
  NAND3_X1  g722(.A1(new_n1147), .A2(new_n845), .A3(new_n1148), .ZN(G225));
  INV_X1    g723(.A(G225), .ZN(G308));
endmodule


