//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 0 1 0 1 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 1 0 1 0 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965;
  XNOR2_X1  g000(.A(G143), .B(G146), .ZN(new_n187));
  NAND3_X1  g001(.A1(new_n187), .A2(KEYINPUT0), .A3(G128), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT0), .B(G128), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n187), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  AND2_X1   g005(.A1(KEYINPUT64), .A2(G134), .ZN(new_n192));
  NOR2_X1   g006(.A1(KEYINPUT64), .A2(G134), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n191), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT11), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n192), .A2(new_n193), .ZN(new_n197));
  AOI21_X1  g011(.A(KEYINPUT67), .B1(new_n197), .B2(G137), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n199));
  INV_X1    g013(.A(G134), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(KEYINPUT64), .A2(G134), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n201), .A2(KEYINPUT67), .A3(G137), .A4(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n196), .B1(new_n198), .B2(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT65), .B(G137), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT11), .A2(G134), .ZN(new_n207));
  AOI21_X1  g021(.A(KEYINPUT66), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n191), .A2(KEYINPUT65), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G137), .ZN(new_n211));
  AND4_X1   g025(.A1(KEYINPUT66), .A2(new_n209), .A3(new_n211), .A4(new_n207), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n208), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(G131), .B1(new_n205), .B2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n209), .A2(new_n211), .A3(new_n207), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n206), .A2(KEYINPUT66), .A3(new_n207), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n201), .A2(G137), .A3(new_n202), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n203), .ZN(new_n223));
  INV_X1    g037(.A(G131), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n219), .A2(new_n223), .A3(new_n224), .A4(new_n196), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n190), .B1(new_n214), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G128), .ZN(new_n227));
  INV_X1    g041(.A(G146), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G143), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n227), .B1(new_n229), .B2(KEYINPUT1), .ZN(new_n230));
  INV_X1    g044(.A(G143), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G146), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n229), .B(new_n232), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n237), .B1(new_n206), .B2(G134), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n210), .A2(G137), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n191), .A2(KEYINPUT65), .ZN(new_n240));
  OAI211_X1 g054(.A(KEYINPUT68), .B(new_n200), .C1(new_n239), .C2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n238), .A2(new_n194), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n236), .B1(new_n242), .B2(G131), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n243), .A2(new_n225), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n226), .A2(new_n244), .ZN(new_n245));
  XOR2_X1   g059(.A(KEYINPUT2), .B(G113), .Z(new_n246));
  INV_X1    g060(.A(G119), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT70), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G119), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n248), .A2(new_n250), .A3(G116), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n247), .A2(G116), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n246), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT71), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT70), .B(G119), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n252), .B1(new_n256), .B2(G116), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT71), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n258), .A3(new_n246), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n246), .B1(new_n251), .B2(new_n253), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(KEYINPUT72), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT72), .ZN(new_n264));
  AOI211_X1 g078(.A(new_n264), .B(new_n261), .C1(new_n255), .C2(new_n259), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n245), .A2(new_n266), .ZN(new_n267));
  OAI22_X1  g081(.A1(new_n226), .A2(new_n244), .B1(new_n263), .B2(new_n265), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(KEYINPUT78), .A3(new_n268), .ZN(new_n269));
  OR3_X1    g083(.A1(new_n245), .A2(KEYINPUT78), .A3(new_n266), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(new_n270), .A3(KEYINPUT28), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT79), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT28), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n271), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n269), .A2(new_n270), .A3(KEYINPUT79), .A4(KEYINPUT28), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  XOR2_X1   g091(.A(KEYINPUT26), .B(G101), .Z(new_n278));
  XNOR2_X1  g092(.A(new_n278), .B(KEYINPUT74), .ZN(new_n279));
  INV_X1    g093(.A(G210), .ZN(new_n280));
  NOR3_X1   g094(.A1(new_n280), .A2(G237), .A3(G953), .ZN(new_n281));
  XOR2_X1   g095(.A(new_n279), .B(new_n281), .Z(new_n282));
  XNOR2_X1  g096(.A(KEYINPUT73), .B(KEYINPUT27), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n282), .B(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT29), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(G902), .B1(new_n277), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n274), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n268), .A2(KEYINPUT75), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT75), .ZN(new_n291));
  INV_X1    g105(.A(new_n190), .ZN(new_n292));
  AND4_X1   g106(.A1(new_n224), .A2(new_n219), .A3(new_n223), .A4(new_n196), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n222), .A2(new_n203), .B1(new_n195), .B2(new_n194), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n224), .B1(new_n294), .B2(new_n219), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n292), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n243), .A2(new_n225), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n258), .B1(new_n257), .B2(new_n246), .ZN(new_n299));
  AND4_X1   g113(.A1(new_n258), .A2(new_n246), .A3(new_n251), .A4(new_n253), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n262), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n264), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n260), .A2(KEYINPUT72), .A3(new_n262), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n291), .B1(new_n298), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n267), .B1(new_n290), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n289), .B1(new_n306), .B2(KEYINPUT28), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n284), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT77), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n298), .A2(new_n304), .ZN(new_n310));
  NAND2_X1  g124(.A1(KEYINPUT69), .A2(KEYINPUT30), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT69), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT30), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n311), .B(new_n314), .C1(new_n226), .C2(new_n244), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n296), .A2(new_n312), .A3(new_n313), .A4(new_n297), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n310), .B1(new_n317), .B2(new_n304), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n309), .B1(new_n318), .B2(new_n284), .ZN(new_n319));
  INV_X1    g133(.A(new_n318), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(KEYINPUT77), .A3(new_n285), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n308), .A2(new_n319), .A3(new_n286), .A4(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n288), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G472), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT76), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n325), .B1(new_n307), .B2(new_n284), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n317), .A2(new_n304), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n327), .A2(new_n284), .A3(new_n267), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT31), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n318), .A2(KEYINPUT31), .A3(new_n284), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n268), .A2(KEYINPUT75), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n298), .A2(new_n291), .A3(new_n304), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n310), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n274), .B1(new_n335), .B2(new_n273), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(KEYINPUT76), .A3(new_n285), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n326), .A2(new_n332), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT32), .ZN(new_n339));
  NOR2_X1   g153(.A1(G472), .A2(G902), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n339), .B1(new_n338), .B2(new_n340), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n324), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT25), .ZN(new_n344));
  XNOR2_X1  g158(.A(G125), .B(G140), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT16), .ZN(new_n346));
  INV_X1    g160(.A(G125), .ZN(new_n347));
  OR3_X1    g161(.A1(new_n347), .A2(KEYINPUT16), .A3(G140), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(G146), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n345), .A2(new_n228), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G110), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n227), .A2(KEYINPUT23), .A3(G119), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n256), .A2(G128), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT81), .B(KEYINPUT23), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(KEYINPUT82), .A3(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n356), .B1(G128), .B2(new_n256), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT82), .B1(new_n354), .B2(new_n355), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n352), .B(new_n353), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n354), .B1(new_n247), .B2(G128), .ZN(new_n360));
  XNOR2_X1  g174(.A(KEYINPUT24), .B(G110), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n351), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n349), .ZN(new_n364));
  AOI21_X1  g178(.A(G146), .B1(new_n346), .B2(new_n348), .ZN(new_n365));
  OAI22_X1  g179(.A1(new_n364), .A2(new_n365), .B1(new_n360), .B2(new_n361), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n353), .B1(new_n357), .B2(new_n358), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n366), .B1(new_n367), .B2(G110), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(KEYINPUT22), .B(G137), .ZN(new_n370));
  INV_X1    g184(.A(G953), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n371), .A2(G221), .A3(G234), .ZN(new_n372));
  XOR2_X1   g186(.A(new_n370), .B(new_n372), .Z(new_n373));
  NAND2_X1  g187(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n373), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n375), .B1(new_n363), .B2(new_n368), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n344), .B1(new_n377), .B2(G902), .ZN(new_n378));
  INV_X1    g192(.A(G902), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n374), .A2(new_n376), .A3(KEYINPUT25), .A4(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  XOR2_X1   g195(.A(KEYINPUT80), .B(G217), .Z(new_n382));
  AOI21_X1  g196(.A(new_n382), .B1(G234), .B2(new_n379), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n383), .A2(G902), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n374), .A2(new_n376), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(KEYINPUT9), .B(G234), .ZN(new_n389));
  OAI21_X1  g203(.A(G221), .B1(new_n389), .B2(G902), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G469), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n214), .A2(new_n225), .ZN(new_n393));
  INV_X1    g207(.A(G104), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT3), .B1(new_n394), .B2(G107), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT3), .ZN(new_n396));
  INV_X1    g210(.A(G107), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(G104), .ZN(new_n398));
  INV_X1    g212(.A(G101), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n394), .A2(G107), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n395), .A2(new_n398), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n394), .A2(G107), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n397), .A2(G104), .ZN(new_n403));
  OAI21_X1  g217(.A(G101), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n234), .A2(new_n401), .A3(new_n404), .A4(new_n235), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT84), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT10), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n405), .B1(new_n406), .B2(KEYINPUT10), .ZN(new_n409));
  OAI22_X1  g223(.A1(new_n408), .A2(new_n409), .B1(new_n406), .B2(KEYINPUT10), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n395), .A2(new_n398), .A3(new_n400), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G101), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(KEYINPUT4), .A3(new_n401), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT83), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n413), .B(new_n414), .C1(KEYINPUT4), .C2(new_n412), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n412), .A2(KEYINPUT83), .A3(KEYINPUT4), .A4(new_n401), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n190), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n393), .B1(new_n410), .B2(new_n417), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n234), .A2(new_n235), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n401), .A2(new_n404), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT10), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n419), .B(new_n421), .C1(KEYINPUT84), .C2(new_n422), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n423), .A2(new_n407), .B1(KEYINPUT84), .B2(new_n422), .ZN(new_n424));
  INV_X1    g238(.A(new_n413), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n414), .B1(new_n412), .B2(KEYINPUT4), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n416), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n292), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n424), .A2(new_n428), .A3(new_n214), .A4(new_n225), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n418), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(G110), .B(G140), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n371), .A2(G227), .ZN(new_n432));
  XOR2_X1   g246(.A(new_n431), .B(new_n432), .Z(new_n433));
  NAND3_X1  g247(.A1(new_n430), .A2(KEYINPUT85), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n433), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n236), .A2(new_n420), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n405), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n393), .A2(KEYINPUT12), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(KEYINPUT12), .B1(new_n393), .B2(new_n437), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n429), .B(new_n435), .C1(new_n438), .C2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n434), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(KEYINPUT85), .B1(new_n430), .B2(new_n433), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n392), .B(new_n379), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n429), .A2(new_n435), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n429), .B1(new_n438), .B2(new_n439), .ZN(new_n445));
  AOI22_X1  g259(.A1(new_n418), .A2(new_n444), .B1(new_n445), .B2(new_n433), .ZN(new_n446));
  OAI21_X1  g260(.A(G469), .B1(new_n446), .B2(G902), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n391), .B1(new_n443), .B2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(G110), .B(G122), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n302), .A2(new_n303), .B1(new_n415), .B2(new_n416), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n257), .A2(KEYINPUT5), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n452), .B(G113), .C1(KEYINPUT5), .C2(new_n251), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(new_n260), .A3(new_n421), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n450), .B1(new_n451), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n427), .B1(new_n263), .B2(new_n265), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(new_n454), .A3(new_n449), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n456), .A2(KEYINPUT6), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n419), .A2(new_n347), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n460), .B1(new_n347), .B2(new_n190), .ZN(new_n461));
  INV_X1    g275(.A(G224), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n462), .A2(G953), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(KEYINPUT86), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n461), .B(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT6), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n466), .B(new_n450), .C1(new_n451), .C2(new_n455), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n459), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT7), .ZN(new_n469));
  OR3_X1    g283(.A1(new_n461), .A2(new_n469), .A3(new_n463), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n461), .B1(new_n469), .B2(new_n463), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n453), .A2(new_n260), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n420), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n454), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n449), .B(KEYINPUT8), .ZN(new_n475));
  AOI22_X1  g289(.A1(new_n470), .A2(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(G902), .B1(new_n476), .B2(new_n458), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n468), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(G210), .B1(G237), .B2(G902), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n468), .A2(new_n477), .A3(new_n479), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(G214), .B1(G237), .B2(G902), .ZN(new_n484));
  INV_X1    g298(.A(G952), .ZN(new_n485));
  AOI211_X1 g299(.A(G953), .B(new_n485), .C1(G234), .C2(G237), .ZN(new_n486));
  XNOR2_X1  g300(.A(KEYINPUT21), .B(G898), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(KEYINPUT94), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  AOI211_X1 g303(.A(new_n379), .B(new_n371), .C1(G234), .C2(G237), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n486), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n448), .A2(new_n483), .A3(new_n484), .A4(new_n492), .ZN(new_n493));
  NOR3_X1   g307(.A1(new_n382), .A2(G953), .A3(new_n389), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT91), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n496), .B1(new_n227), .B2(G143), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n231), .A2(KEYINPUT91), .A3(G128), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n499), .B1(G128), .B2(new_n231), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n500), .A2(new_n193), .A3(new_n192), .ZN(new_n501));
  XOR2_X1   g315(.A(G116), .B(G122), .Z(new_n502));
  XNOR2_X1  g316(.A(new_n502), .B(new_n397), .ZN(new_n503));
  OR2_X1    g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT13), .ZN(new_n505));
  AOI22_X1  g319(.A1(new_n499), .A2(new_n505), .B1(new_n227), .B2(G143), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n506), .B1(new_n505), .B2(new_n499), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT92), .B1(new_n507), .B2(G134), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n507), .A2(KEYINPUT92), .A3(G134), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n504), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n500), .B(new_n197), .ZN(new_n512));
  INV_X1    g326(.A(G122), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(G116), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n397), .B1(new_n514), .B2(KEYINPUT14), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n502), .B(new_n515), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n495), .B1(new_n511), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n517), .ZN(new_n519));
  INV_X1    g333(.A(new_n510), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n520), .A2(new_n508), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n519), .B(new_n494), .C1(new_n521), .C2(new_n504), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n518), .A2(KEYINPUT93), .A3(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT93), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n524), .B(new_n495), .C1(new_n511), .C2(new_n517), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(new_n379), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(G478), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n527), .A2(KEYINPUT15), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n528), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n523), .A2(new_n379), .A3(new_n525), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(G475), .A2(G902), .ZN(new_n534));
  XOR2_X1   g348(.A(KEYINPUT87), .B(G143), .Z(new_n535));
  INV_X1    g349(.A(G237), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n536), .A2(new_n371), .A3(G214), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT87), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n537), .B1(new_n540), .B2(new_n231), .ZN(new_n541));
  OAI21_X1  g355(.A(G131), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT17), .ZN(new_n543));
  OR2_X1    g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT90), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(new_n364), .B2(new_n365), .ZN(new_n546));
  INV_X1    g360(.A(new_n365), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n547), .A2(KEYINPUT90), .A3(new_n349), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n538), .B1(KEYINPUT87), .B2(G143), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n549), .B(new_n224), .C1(new_n538), .C2(new_n535), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n542), .A2(new_n550), .A3(new_n543), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n544), .A2(new_n546), .A3(new_n548), .A4(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(G113), .B(G122), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(new_n394), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT18), .ZN(new_n555));
  OAI221_X1 g369(.A(new_n549), .B1(new_n555), .B2(new_n224), .C1(new_n538), .C2(new_n535), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n345), .B(new_n228), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n556), .B(new_n557), .C1(new_n555), .C2(new_n542), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n552), .A2(new_n554), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n345), .A2(new_n560), .ZN(new_n561));
  XOR2_X1   g375(.A(KEYINPUT88), .B(KEYINPUT19), .Z(new_n562));
  OAI21_X1  g376(.A(new_n561), .B1(new_n345), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n349), .B1(new_n563), .B2(G146), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT89), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n542), .A2(new_n550), .ZN(new_n567));
  OAI211_X1 g381(.A(KEYINPUT89), .B(new_n349), .C1(new_n563), .C2(G146), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n554), .B1(new_n569), .B2(new_n558), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n534), .B1(new_n559), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT20), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT20), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n573), .B(new_n534), .C1(new_n559), .C2(new_n570), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n554), .B1(new_n552), .B2(new_n558), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n379), .B1(new_n559), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g390(.A1(new_n572), .A2(new_n574), .B1(G475), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n533), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n493), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n343), .A2(new_n388), .A3(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(G101), .ZN(G3));
  NAND2_X1  g395(.A1(new_n338), .A2(new_n379), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(G472), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n583), .A2(KEYINPUT95), .B1(new_n340), .B2(new_n338), .ZN(new_n584));
  INV_X1    g398(.A(G472), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n585), .B1(new_n338), .B2(new_n379), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT95), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n443), .A2(new_n447), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n390), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n589), .A2(new_n387), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(KEYINPUT96), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT98), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n481), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n478), .A2(KEYINPUT98), .A3(new_n480), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT97), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n482), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n482), .A2(new_n597), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n595), .B(new_n596), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n484), .ZN(new_n601));
  INV_X1    g415(.A(new_n577), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n523), .A2(new_n603), .A3(new_n525), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n518), .A2(KEYINPUT33), .A3(new_n522), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n604), .A2(G478), .A3(new_n379), .A4(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT99), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n526), .A2(new_n527), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n607), .B1(new_n606), .B2(new_n608), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n602), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n601), .A2(new_n491), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n593), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(G104), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G6));
  NOR2_X1   g430(.A1(new_n533), .A2(new_n602), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n601), .A2(new_n491), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n593), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT102), .B(G107), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT101), .B(KEYINPUT35), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G9));
  INV_X1    g438(.A(new_n579), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n375), .A2(KEYINPUT36), .ZN(new_n626));
  XOR2_X1   g440(.A(new_n369), .B(new_n626), .Z(new_n627));
  AOI22_X1  g441(.A1(new_n381), .A2(new_n383), .B1(new_n385), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n584), .A2(new_n588), .A3(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT103), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n625), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n584), .A2(KEYINPUT103), .A3(new_n588), .A4(new_n629), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT37), .B(G110), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G12));
  INV_X1    g450(.A(new_n486), .ZN(new_n637));
  INV_X1    g451(.A(new_n490), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n637), .B1(new_n638), .B2(G900), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n617), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n591), .A2(new_n628), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n640), .A2(new_n484), .A3(new_n641), .A4(new_n600), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n585), .B1(new_n288), .B2(new_n322), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n332), .A2(new_n337), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT76), .B1(new_n336), .B2(new_n285), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n340), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT32), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n643), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n642), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(new_n227), .ZN(G30));
  XNOR2_X1  g465(.A(new_n639), .B(KEYINPUT39), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n591), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(KEYINPUT40), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(KEYINPUT40), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n483), .B(KEYINPUT38), .ZN(new_n658));
  INV_X1    g472(.A(new_n484), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n533), .A2(new_n577), .A3(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n657), .A2(new_n628), .A3(new_n658), .A4(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n647), .A2(new_n648), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n320), .A2(new_n284), .ZN(new_n663));
  AND2_X1   g477(.A1(new_n269), .A2(new_n270), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n663), .B(new_n379), .C1(new_n284), .C2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(G472), .ZN(new_n666));
  AOI21_X1  g480(.A(KEYINPUT104), .B1(new_n662), .B2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n662), .A2(KEYINPUT104), .A3(new_n666), .ZN(new_n669));
  AOI211_X1 g483(.A(new_n656), .B(new_n661), .C1(new_n668), .C2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(new_n231), .ZN(G45));
  NOR3_X1   g485(.A1(new_n601), .A2(new_n591), .A3(new_n628), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n602), .B(new_n639), .C1(new_n609), .C2(new_n610), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n672), .A2(new_n343), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G146), .ZN(G48));
  AOI21_X1  g490(.A(new_n387), .B1(new_n662), .B2(new_n324), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n379), .B1(new_n441), .B2(new_n442), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(G469), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n680), .A2(new_n390), .A3(new_n443), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n683), .A2(new_n612), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT41), .B(G113), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G15));
  AND2_X1   g500(.A1(new_n683), .A2(new_n619), .ZN(new_n687));
  XOR2_X1   g501(.A(new_n687), .B(G116), .Z(G18));
  INV_X1    g502(.A(KEYINPUT105), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n577), .A2(new_n529), .A3(new_n531), .A4(new_n492), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n628), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n600), .A2(new_n681), .A3(new_n691), .A4(new_n484), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n689), .B1(new_n649), .B2(new_n692), .ZN(new_n693));
  AND4_X1   g507(.A1(new_n484), .A2(new_n600), .A3(new_n681), .A4(new_n691), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n343), .A3(KEYINPUT105), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  NAND2_X1  g511(.A1(new_n600), .A2(new_n660), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n600), .A2(new_n660), .A3(KEYINPUT107), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n682), .A2(new_n491), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n704));
  INV_X1    g518(.A(new_n340), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n275), .A2(new_n285), .A3(new_n276), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n705), .B1(new_n706), .B2(new_n332), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n707), .B1(new_n582), .B2(G472), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n704), .B1(new_n708), .B2(new_n388), .ZN(new_n709));
  NOR4_X1   g523(.A1(new_n586), .A2(KEYINPUT106), .A3(new_n387), .A4(new_n707), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n702), .B(new_n703), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G122), .ZN(G24));
  NOR3_X1   g526(.A1(new_n601), .A2(new_n682), .A3(new_n673), .ZN(new_n713));
  AOI21_X1  g527(.A(KEYINPUT108), .B1(new_n708), .B2(new_n629), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n715));
  NOR4_X1   g529(.A1(new_n586), .A2(new_n715), .A3(new_n628), .A4(new_n707), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n713), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G125), .ZN(G27));
  NOR2_X1   g532(.A1(new_n483), .A2(new_n659), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n448), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n720), .A2(new_n673), .ZN(new_n721));
  AOI21_X1  g535(.A(KEYINPUT42), .B1(new_n677), .B2(new_n721), .ZN(new_n722));
  AND4_X1   g536(.A1(KEYINPUT42), .A2(new_n343), .A3(new_n388), .A4(new_n721), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(new_n224), .ZN(G33));
  AND3_X1   g539(.A1(new_n640), .A2(new_n448), .A3(new_n719), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n677), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G134), .ZN(G36));
  OAI21_X1  g542(.A(new_n577), .B1(new_n609), .B2(new_n610), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT109), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(KEYINPUT43), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(new_n589), .A3(new_n629), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT111), .ZN(new_n734));
  OR3_X1    g548(.A1(new_n733), .A2(new_n734), .A3(KEYINPUT44), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n734), .B1(new_n733), .B2(KEYINPUT44), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n446), .A2(KEYINPUT45), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n446), .A2(KEYINPUT45), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(G469), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(G469), .A2(G902), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT46), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n739), .A2(KEYINPUT46), .A3(new_n740), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(new_n443), .A3(new_n744), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n745), .A2(new_n390), .ZN(new_n746));
  XOR2_X1   g560(.A(new_n719), .B(KEYINPUT110), .Z(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(new_n652), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n748), .B1(new_n733), .B2(KEYINPUT44), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n735), .A2(new_n736), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G137), .ZN(G39));
  OR2_X1    g565(.A1(new_n746), .A2(KEYINPUT47), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n746), .A2(KEYINPUT47), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n719), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n673), .A2(new_n755), .A3(new_n388), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n754), .A2(new_n649), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G140), .ZN(G42));
  INV_X1    g572(.A(new_n669), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n759), .A2(new_n667), .A3(new_n387), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n680), .A2(new_n443), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT49), .ZN(new_n762));
  AOI211_X1 g576(.A(new_n391), .B(new_n659), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n763), .B1(new_n762), .B2(new_n761), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n764), .A2(new_n658), .A3(new_n729), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n760), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n721), .B1(new_n714), .B2(new_n716), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n533), .A2(new_n577), .A3(new_n639), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n720), .A2(new_n628), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n343), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n768), .A2(new_n727), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n724), .A2(new_n772), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n677), .B(new_n681), .C1(new_n612), .C2(new_n619), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(new_n696), .A3(new_n711), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT112), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n774), .A2(new_n696), .A3(new_n711), .A4(KEYINPUT112), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n532), .A2(KEYINPUT113), .A3(new_n577), .ZN(new_n779));
  AOI21_X1  g593(.A(KEYINPUT113), .B1(new_n532), .B2(new_n577), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n493), .B1(new_n781), .B2(new_n611), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n584), .A2(new_n782), .A3(new_n388), .A4(new_n588), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n580), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n784), .B1(new_n632), .B2(new_n633), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n773), .A2(new_n777), .A3(new_n778), .A4(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n672), .A2(new_n343), .A3(new_n640), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n717), .A2(new_n787), .A3(new_n675), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT114), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n628), .A2(new_n639), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n789), .B1(new_n790), .B2(new_n591), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n448), .A2(KEYINPUT114), .A3(new_n628), .A4(new_n639), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n701), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT107), .B1(new_n600), .B2(new_n660), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n796), .B1(new_n668), .B2(new_n669), .ZN(new_n797));
  OAI21_X1  g611(.A(KEYINPUT52), .B1(new_n788), .B2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n707), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n583), .A2(new_n629), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n715), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n708), .A2(KEYINPUT108), .A3(new_n629), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n650), .B1(new_n803), .B2(new_n713), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n702), .B(new_n793), .C1(new_n759), .C2(new_n667), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n804), .A2(new_n805), .A3(new_n806), .A4(new_n675), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n798), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n767), .B1(new_n786), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(KEYINPUT115), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT115), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n811), .B(new_n767), .C1(new_n786), .C2(new_n808), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n768), .A2(new_n727), .A3(new_n771), .A4(KEYINPUT53), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n806), .B1(new_n717), .B2(new_n787), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n817), .A2(new_n798), .A3(new_n807), .A4(new_n785), .ZN(new_n818));
  OR3_X1    g632(.A1(new_n775), .A2(new_n724), .A3(KEYINPUT116), .ZN(new_n819));
  OAI21_X1  g633(.A(KEYINPUT116), .B1(new_n775), .B2(new_n724), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n818), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n813), .A2(new_n814), .A3(new_n822), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n798), .A2(new_n807), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n773), .A2(new_n785), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n777), .A2(new_n778), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n767), .B1(new_n804), .B2(new_n806), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n824), .A2(new_n825), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n814), .B1(new_n828), .B2(new_n809), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n823), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT119), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n682), .A2(new_n832), .A3(new_n755), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT119), .B1(new_n681), .B2(new_n719), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n833), .A2(new_n637), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n760), .A2(new_n835), .ZN(new_n836));
  OR4_X1    g650(.A1(new_n602), .A2(new_n836), .A3(new_n609), .A4(new_n610), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n835), .A2(new_n803), .A3(new_n731), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n709), .A2(new_n710), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n840), .A2(new_n486), .A3(new_n731), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n747), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  AOI22_X1  g657(.A1(new_n754), .A2(KEYINPUT117), .B1(new_n391), .B2(new_n761), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n844), .B1(KEYINPUT117), .B2(new_n754), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n839), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n658), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n682), .A2(new_n484), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT118), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n848), .A2(KEYINPUT118), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n841), .A2(new_n847), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT50), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT51), .B1(new_n846), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n601), .A2(new_n682), .ZN(new_n855));
  AOI211_X1 g669(.A(new_n485), .B(G953), .C1(new_n841), .C2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n835), .A2(new_n677), .A3(new_n731), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT48), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n761), .A2(new_n391), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n752), .A2(new_n753), .A3(new_n860), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n861), .A2(KEYINPUT120), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(KEYINPUT120), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n843), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n837), .A2(new_n864), .A3(KEYINPUT51), .A4(new_n838), .ZN(new_n865));
  OAI221_X1 g679(.A(new_n859), .B1(new_n611), .B2(new_n836), .C1(new_n865), .C2(new_n852), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n831), .A2(new_n854), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(G952), .A2(G953), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n766), .B1(new_n867), .B2(new_n868), .ZN(G75));
  NAND2_X1  g683(.A1(new_n459), .A2(new_n467), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(new_n465), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT55), .Z(new_n872));
  AOI21_X1  g686(.A(new_n821), .B1(new_n810), .B2(new_n812), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n873), .A2(new_n280), .A3(new_n379), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n872), .B1(new_n874), .B2(KEYINPUT56), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n371), .A2(G952), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT123), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g692(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n872), .A2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(KEYINPUT122), .B1(new_n874), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n813), .A2(new_n822), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n883), .A2(G210), .A3(G902), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT122), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n884), .A2(new_n885), .A3(new_n880), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n878), .B1(new_n882), .B2(new_n886), .ZN(G51));
  AOI21_X1  g701(.A(new_n814), .B1(new_n813), .B2(new_n822), .ZN(new_n888));
  AOI211_X1 g702(.A(KEYINPUT54), .B(new_n821), .C1(new_n810), .C2(new_n812), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n740), .B(KEYINPUT57), .ZN(new_n891));
  OAI22_X1  g705(.A1(new_n890), .A2(new_n891), .B1(new_n442), .B2(new_n441), .ZN(new_n892));
  OR3_X1    g706(.A1(new_n873), .A2(new_n379), .A3(new_n739), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n876), .B1(new_n892), .B2(new_n893), .ZN(G54));
  NOR2_X1   g708(.A1(new_n873), .A2(new_n379), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n559), .A2(new_n570), .ZN(new_n896));
  AND2_X1   g710(.A1(KEYINPUT58), .A2(G475), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n896), .B1(new_n895), .B2(new_n897), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n898), .A2(new_n899), .A3(new_n876), .ZN(G60));
  NAND2_X1  g714(.A1(new_n604), .A2(new_n605), .ZN(new_n901));
  NAND2_X1  g715(.A1(G478), .A2(G902), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT59), .Z(new_n903));
  NOR2_X1   g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n904), .B1(new_n888), .B2(new_n889), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n877), .ZN(new_n906));
  INV_X1    g720(.A(new_n901), .ZN(new_n907));
  INV_X1    g721(.A(new_n903), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n907), .B1(new_n831), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT124), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n829), .B1(new_n873), .B2(new_n814), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n901), .B1(new_n911), .B2(new_n903), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT124), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n912), .A2(new_n913), .A3(new_n877), .A4(new_n905), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n910), .A2(new_n914), .ZN(G63));
  NAND2_X1  g729(.A1(G217), .A2(G902), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT60), .Z(new_n917));
  NAND2_X1  g731(.A1(new_n883), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n377), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n627), .B(KEYINPUT125), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n883), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n919), .A2(new_n877), .A3(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT61), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n919), .A2(KEYINPUT61), .A3(new_n877), .A4(new_n921), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(G66));
  OAI21_X1  g740(.A(G953), .B1(new_n489), .B2(new_n462), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n826), .A2(new_n785), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n927), .B1(new_n929), .B2(G953), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n870), .B1(G898), .B2(new_n371), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT126), .Z(new_n932));
  XNOR2_X1  g746(.A(new_n930), .B(new_n932), .ZN(G69));
  OR2_X1    g747(.A1(new_n670), .A2(new_n788), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n934), .A2(KEYINPUT62), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n654), .A2(new_n719), .ZN(new_n936));
  AOI211_X1 g750(.A(new_n936), .B(new_n678), .C1(new_n611), .C2(new_n781), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n934), .A2(KEYINPUT62), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n938), .A2(new_n750), .A3(new_n757), .A4(new_n939), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n940), .A2(new_n371), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n317), .B(new_n563), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n371), .A2(G900), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n746), .A2(new_n652), .A3(new_n702), .ZN(new_n945));
  INV_X1    g759(.A(new_n726), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n678), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n947), .A2(new_n724), .A3(new_n788), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n750), .A2(new_n757), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n944), .B1(new_n949), .B2(new_n371), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT127), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n943), .B1(new_n950), .B2(new_n951), .ZN(new_n953));
  OAI22_X1  g767(.A1(new_n941), .A2(new_n943), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n371), .B1(G227), .B2(G900), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n954), .B(new_n955), .ZN(G72));
  OR2_X1    g770(.A1(new_n940), .A2(new_n928), .ZN(new_n957));
  NAND2_X1  g771(.A1(G472), .A2(G902), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT63), .Z(new_n959));
  AOI21_X1  g773(.A(new_n663), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n321), .A2(new_n328), .A3(new_n319), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n959), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n962), .B1(new_n828), .B2(new_n809), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n959), .B1(new_n949), .B2(new_n928), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n964), .A2(new_n285), .A3(new_n318), .ZN(new_n965));
  NOR4_X1   g779(.A1(new_n960), .A2(new_n876), .A3(new_n963), .A4(new_n965), .ZN(G57));
endmodule


