//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 0 0 0 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 1 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 1 0 1 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1263, new_n1264, new_n1265, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n204), .C2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT65), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n204), .A2(new_n205), .ZN(new_n214));
  INV_X1    g0014(.A(G50), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  INV_X1    g0017(.A(G20), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  XOR2_X1   g0020(.A(KEYINPUT66), .B(G244), .Z(new_n221));
  INV_X1    g0021(.A(G77), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G107), .A2(G264), .ZN(new_n227));
  NAND4_X1  g0027(.A1(new_n224), .A2(new_n225), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n210), .B1(new_n223), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n213), .B(new_n220), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n215), .A2(G68), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n203), .A2(G50), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n243), .B(new_n248), .ZN(G351));
  AND2_X1   g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  OAI21_X1  g0050(.A(KEYINPUT67), .B1(new_n250), .B2(new_n217), .ZN(new_n251));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n252), .B1(G41), .B2(G45), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT67), .ZN(new_n256));
  NAND4_X1  g0056(.A1(new_n255), .A2(new_n256), .A3(G1), .A4(G13), .ZN(new_n257));
  NAND4_X1  g0057(.A1(new_n251), .A2(new_n254), .A3(G274), .A4(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n251), .A2(new_n257), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(new_n254), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT68), .B(G226), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G1698), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n263), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(new_n264), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n267), .A2(G223), .B1(new_n269), .B2(G77), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT3), .B(G33), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(G222), .A3(new_n263), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n250), .A2(new_n217), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n258), .B(new_n262), .C1(new_n273), .C2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G190), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n278), .B1(G200), .B2(new_n276), .ZN(new_n279));
  AOI21_X1  g0079(.A(KEYINPUT10), .B1(new_n279), .B2(KEYINPUT70), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n217), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT69), .ZN(new_n283));
  INV_X1    g0083(.A(G33), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n283), .B1(new_n284), .B2(G20), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n218), .A2(KEYINPUT69), .A3(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT8), .B(G58), .ZN(new_n289));
  INV_X1    g0089(.A(G150), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G20), .A2(G33), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  OAI22_X1  g0092(.A1(new_n288), .A2(new_n289), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n218), .B1(new_n214), .B2(new_n215), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n282), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n252), .A2(G13), .A3(G20), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(new_n282), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n252), .A2(G20), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n298), .A2(G50), .A3(new_n299), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n295), .B(new_n300), .C1(G50), .C2(new_n296), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n301), .B(KEYINPUT9), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n279), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n280), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n279), .B(new_n302), .C1(KEYINPUT70), .C2(KEYINPUT10), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n276), .A2(G179), .ZN(new_n306));
  INV_X1    g0106(.A(G169), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n276), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n306), .A2(new_n301), .A3(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n304), .A2(new_n305), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n282), .ZN(new_n311));
  INV_X1    g0111(.A(new_n289), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n312), .A2(new_n291), .B1(G20), .B2(G77), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT15), .B(G87), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n287), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n311), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n298), .A2(G77), .A3(new_n299), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n318), .B1(G77), .B2(new_n296), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n259), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n253), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n323), .A2(new_n221), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n267), .A2(G238), .B1(new_n269), .B2(G107), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n271), .A2(G232), .A3(new_n263), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n274), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n324), .A2(new_n258), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n321), .B1(new_n330), .B2(G190), .ZN(new_n331));
  INV_X1    g0131(.A(G200), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n331), .B1(new_n332), .B2(new_n330), .ZN(new_n333));
  INV_X1    g0133(.A(G179), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n329), .A2(new_n307), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(new_n321), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n310), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT71), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n267), .A2(new_n340), .A3(G232), .ZN(new_n341));
  OAI211_X1 g0141(.A(G232), .B(G1698), .C1(new_n268), .C2(new_n264), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT71), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  OAI211_X1 g0144(.A(G226), .B(new_n263), .C1(new_n268), .C2(new_n264), .ZN(new_n345));
  NAND2_X1  g0145(.A1(G33), .A2(G97), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n349), .A2(KEYINPUT72), .A3(new_n274), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT72), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n347), .B1(new_n341), .B2(new_n343), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n351), .B1(new_n352), .B2(new_n275), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT13), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT73), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n323), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G238), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n358), .B1(new_n260), .B2(KEYINPUT73), .ZN(new_n359));
  INV_X1    g0159(.A(G274), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n259), .A2(new_n360), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n357), .A2(new_n359), .B1(new_n254), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n354), .A2(new_n355), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n355), .B1(new_n354), .B2(new_n362), .ZN(new_n365));
  OAI21_X1  g0165(.A(G200), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n288), .A2(new_n222), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n292), .A2(new_n215), .B1(new_n218), .B2(G68), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n282), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT11), .ZN(new_n370));
  OR2_X1    g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n297), .A2(KEYINPUT74), .A3(new_n203), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT12), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT74), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n296), .B2(G68), .ZN(new_n375));
  OR2_X1    g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n373), .A2(new_n375), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n298), .A2(G68), .A3(new_n299), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n369), .A2(new_n370), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n371), .A2(new_n378), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  XNOR2_X1  g0181(.A(new_n381), .B(KEYINPUT75), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT72), .B1(new_n349), .B2(new_n274), .ZN(new_n383));
  NOR3_X1   g0183(.A1(new_n352), .A2(new_n351), .A3(new_n275), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n362), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT13), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n386), .A2(G190), .A3(new_n363), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n366), .A2(new_n382), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n307), .A2(KEYINPUT76), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(new_n364), .B2(new_n365), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT14), .ZN(new_n392));
  INV_X1    g0192(.A(new_n390), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n386), .B2(new_n363), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT14), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n386), .A2(G179), .A3(new_n363), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n392), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n382), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n389), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n298), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n312), .A2(new_n299), .ZN(new_n402));
  OAI22_X1  g0202(.A1(new_n401), .A2(new_n402), .B1(new_n296), .B2(new_n312), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(KEYINPUT7), .B1(new_n269), .B2(new_n218), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT7), .ZN(new_n406));
  NOR4_X1   g0206(.A1(new_n268), .A2(new_n264), .A3(new_n406), .A4(G20), .ZN(new_n407));
  OAI21_X1  g0207(.A(G68), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n204), .B(new_n205), .C1(new_n202), .C2(new_n203), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n409), .A2(G20), .B1(G159), .B2(new_n291), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT16), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n311), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n408), .A2(KEYINPUT16), .A3(new_n410), .ZN(new_n414));
  AOI21_X1  g0214(.A(KEYINPUT77), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n406), .B1(new_n271), .B2(G20), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n269), .A2(KEYINPUT7), .A3(new_n218), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n203), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n202), .A2(new_n203), .ZN(new_n419));
  OAI21_X1  g0219(.A(G20), .B1(new_n214), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n291), .A2(G159), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n412), .B1(new_n418), .B2(new_n422), .ZN(new_n423));
  AND4_X1   g0223(.A1(KEYINPUT77), .A2(new_n423), .A3(new_n282), .A4(new_n414), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n404), .B1(new_n415), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(G223), .A2(G1698), .ZN(new_n426));
  INV_X1    g0226(.A(G226), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n426), .B1(new_n427), .B2(G1698), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n428), .A2(new_n271), .B1(G33), .B2(G87), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n258), .B1(new_n429), .B2(new_n275), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n251), .A2(G232), .A3(new_n253), .A4(new_n257), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT78), .ZN(new_n432));
  OR2_X1    g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n432), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n430), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n435), .A2(G179), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n435), .A2(new_n307), .ZN(new_n437));
  OR2_X1    g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT18), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n425), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n423), .A2(new_n282), .A3(new_n414), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT77), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n413), .A2(KEYINPUT77), .A3(new_n414), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n403), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n436), .A2(new_n437), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT18), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n433), .A2(new_n434), .ZN(new_n448));
  INV_X1    g0248(.A(new_n430), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(new_n449), .A3(new_n277), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(new_n435), .B2(G200), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n404), .B(new_n451), .C1(new_n415), .C2(new_n424), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT17), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n445), .A2(KEYINPUT17), .A3(new_n451), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n440), .A2(new_n447), .A3(new_n454), .A4(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n339), .A2(new_n400), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(G107), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n297), .A2(KEYINPUT25), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT25), .B1(new_n297), .B2(new_n459), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n252), .A2(G33), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n296), .A2(new_n463), .A3(new_n217), .A4(new_n281), .ZN(new_n464));
  OAI22_X1  g0264(.A1(new_n461), .A2(new_n462), .B1(new_n459), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n271), .A2(G257), .A3(G1698), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G33), .A2(G294), .ZN(new_n468));
  OAI211_X1 g0268(.A(G250), .B(new_n263), .C1(new_n268), .C2(new_n264), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n274), .ZN(new_n471));
  INV_X1    g0271(.A(G45), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(G1), .ZN(new_n473));
  NAND2_X1  g0273(.A1(KEYINPUT5), .A2(G41), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(KEYINPUT5), .A2(G41), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n473), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n322), .A2(G264), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n252), .A2(G45), .ZN(new_n479));
  OR2_X1    g0279(.A1(KEYINPUT5), .A2(G41), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n479), .B1(new_n480), .B2(new_n474), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n481), .A2(G274), .A3(new_n251), .A4(new_n257), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n471), .A2(new_n478), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n332), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n484), .B1(G190), .B2(new_n483), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT87), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n218), .B(G87), .C1(new_n268), .C2(new_n264), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT22), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT22), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n271), .A2(new_n489), .A3(new_n218), .A4(G87), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n459), .A2(G20), .ZN(new_n492));
  NAND2_X1  g0292(.A1(G33), .A2(G116), .ZN(new_n493));
  OAI22_X1  g0293(.A1(new_n492), .A2(KEYINPUT23), .B1(G20), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n492), .A2(KEYINPUT23), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT86), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n492), .A2(KEYINPUT86), .A3(KEYINPUT23), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n494), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n491), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT24), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT24), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n491), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n486), .B1(new_n504), .B2(new_n282), .ZN(new_n505));
  AOI211_X1 g0305(.A(KEYINPUT87), .B(new_n311), .C1(new_n501), .C2(new_n503), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n466), .B(new_n485), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n259), .A2(new_n481), .ZN(new_n509));
  AOI22_X1  g0309(.A1(G264), .A2(new_n509), .B1(new_n470), .B2(new_n274), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n510), .A2(KEYINPUT88), .A3(G179), .A4(new_n482), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n307), .B1(new_n510), .B2(new_n482), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n471), .A2(new_n478), .A3(G179), .A4(new_n482), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT88), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n511), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n491), .A2(new_n502), .A3(new_n499), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n502), .B1(new_n491), .B2(new_n499), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n282), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT87), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n504), .A2(new_n486), .A3(new_n282), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n516), .B1(new_n522), .B2(new_n466), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n508), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n477), .A2(new_n251), .A3(G257), .A4(new_n257), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n482), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT80), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n482), .A2(new_n525), .A3(KEYINPUT80), .ZN(new_n529));
  OAI211_X1 g0329(.A(G250), .B(G1698), .C1(new_n268), .C2(new_n264), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G283), .ZN(new_n531));
  OAI211_X1 g0331(.A(G244), .B(new_n263), .C1(new_n268), .C2(new_n264), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT4), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n530), .B(new_n531), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n532), .A2(new_n533), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n274), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n528), .A2(new_n529), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT81), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT81), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n528), .A2(new_n536), .A3(new_n539), .A4(new_n529), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n538), .A2(G190), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n537), .A2(G200), .ZN(new_n542));
  OAI211_X1 g0342(.A(KEYINPUT79), .B(G107), .C1(new_n405), .C2(new_n407), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n459), .A2(KEYINPUT6), .A3(G97), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT6), .ZN(new_n546));
  AND2_X1   g0346(.A1(G97), .A2(G107), .ZN(new_n547));
  NOR2_X1   g0347(.A1(G97), .A2(G107), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n550), .A2(G20), .B1(G77), .B2(new_n291), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n543), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n459), .B1(new_n416), .B2(new_n417), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n553), .A2(KEYINPUT79), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n282), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(G97), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n297), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(new_n464), .B2(new_n556), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n542), .A2(new_n555), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n532), .A2(new_n533), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n271), .A2(KEYINPUT4), .A3(G244), .A4(new_n263), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n561), .A2(new_n562), .A3(new_n530), .A4(new_n531), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n527), .A2(new_n526), .B1(new_n563), .B2(new_n274), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n539), .B1(new_n564), .B2(new_n529), .ZN(new_n565));
  INV_X1    g0365(.A(new_n540), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n307), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n537), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n568), .A2(new_n334), .B1(new_n555), .B2(new_n559), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n541), .A2(new_n560), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT83), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n473), .A2(new_n360), .ZN(new_n572));
  INV_X1    g0372(.A(G250), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n479), .A2(new_n573), .ZN(new_n574));
  AND4_X1   g0374(.A1(new_n251), .A2(new_n572), .A3(new_n257), .A4(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(G244), .B(G1698), .C1(new_n268), .C2(new_n264), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT82), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT82), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n271), .A2(new_n578), .A3(G244), .A4(G1698), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n271), .A2(G238), .A3(new_n263), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n577), .A2(new_n579), .A3(new_n493), .A4(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n575), .B1(new_n581), .B2(new_n274), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n334), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n271), .A2(new_n218), .A3(G68), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT19), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n218), .B1(new_n346), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(G87), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n548), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n556), .B1(new_n285), .B2(new_n286), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n584), .B(new_n589), .C1(new_n590), .C2(KEYINPUT19), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n282), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n315), .A2(new_n296), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n592), .B(new_n594), .C1(new_n314), .C2(new_n464), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n583), .B(new_n595), .C1(G169), .C2(new_n582), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n581), .A2(new_n274), .ZN(new_n597));
  INV_X1    g0397(.A(new_n575), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(G190), .A3(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n464), .A2(new_n587), .ZN(new_n600));
  AOI211_X1 g0400(.A(new_n593), .B(new_n600), .C1(new_n591), .C2(new_n282), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n599), .B(new_n601), .C1(new_n332), .C2(new_n582), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n571), .B1(new_n596), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n596), .A2(new_n571), .A3(new_n602), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(G116), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n297), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n311), .A2(G116), .A3(new_n296), .A4(new_n463), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n281), .A2(new_n217), .B1(G20), .B2(new_n607), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n531), .B(new_n218), .C1(G33), .C2(new_n556), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n610), .A2(KEYINPUT20), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT20), .B1(new_n610), .B2(new_n611), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n608), .B(new_n609), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(G264), .B(G1698), .C1(new_n268), .C2(new_n264), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n265), .A2(G303), .A3(new_n266), .ZN(new_n616));
  OAI211_X1 g0416(.A(G257), .B(new_n263), .C1(new_n268), .C2(new_n264), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n618), .A2(new_n274), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n477), .A2(new_n251), .A3(G270), .A4(new_n257), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n482), .A2(new_n620), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n614), .B(G169), .C1(new_n619), .C2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT84), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(KEYINPUT21), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT21), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n622), .A2(new_n623), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n614), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n618), .A2(new_n274), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n629), .A2(G179), .A3(new_n482), .A4(new_n620), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n625), .A2(new_n627), .A3(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n621), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n629), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n628), .B1(new_n635), .B2(new_n277), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n619), .A2(new_n621), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n637), .A2(new_n332), .ZN(new_n638));
  OAI21_X1  g0438(.A(KEYINPUT85), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n614), .B1(new_n637), .B2(G190), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT85), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n640), .B(new_n641), .C1(new_n332), .C2(new_n637), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n633), .B1(new_n639), .B2(new_n642), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n524), .A2(new_n570), .A3(new_n606), .A4(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n458), .A2(new_n644), .ZN(G372));
  INV_X1    g0445(.A(new_n309), .ZN(new_n646));
  INV_X1    g0446(.A(new_n337), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n647), .B1(new_n398), .B2(new_n399), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n388), .A2(new_n454), .A3(new_n455), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n447), .B(new_n440), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n304), .A2(new_n305), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n646), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n458), .ZN(new_n653));
  AOI21_X1  g0453(.A(G169), .B1(new_n538), .B2(new_n540), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n528), .A2(new_n536), .A3(new_n334), .A4(new_n529), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n291), .A2(G77), .ZN(new_n656));
  XNOR2_X1  g0456(.A(G97), .B(G107), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n544), .B1(new_n657), .B2(new_n546), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n656), .B1(new_n658), .B2(new_n218), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n659), .B1(KEYINPUT79), .B2(new_n553), .ZN(new_n660));
  OAI21_X1  g0460(.A(G107), .B1(new_n405), .B2(new_n407), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT79), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n311), .B1(new_n660), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n655), .B1(new_n664), .B2(new_n558), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n654), .A2(new_n665), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n596), .A2(new_n571), .A3(new_n602), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n666), .B(KEYINPUT26), .C1(new_n667), .C2(new_n603), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT26), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n567), .A2(new_n569), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n596), .A2(new_n602), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n631), .B1(new_n624), .B2(KEYINPUT21), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n465), .B1(new_n520), .B2(new_n521), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n627), .B(new_n674), .C1(new_n675), .C2(new_n516), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n671), .B1(new_n675), .B2(new_n485), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(new_n570), .A3(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n673), .A2(new_n596), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n653), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n652), .A2(new_n680), .ZN(G369));
  NAND3_X1  g0481(.A1(new_n252), .A2(new_n218), .A3(G13), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n683), .A2(G213), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G343), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n524), .B1(new_n675), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n466), .B1(new_n505), .B2(new_n506), .ZN(new_n688));
  INV_X1    g0488(.A(new_n516), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n687), .B1(new_n690), .B2(new_n686), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n628), .A2(new_n686), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n633), .A2(new_n692), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n625), .A2(new_n627), .A3(new_n632), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n642), .A2(new_n639), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n693), .B1(new_n696), .B2(new_n692), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n691), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n633), .A2(new_n686), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n524), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n686), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n702), .B1(new_n690), .B2(new_n703), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n699), .A2(new_n704), .ZN(G399));
  NOR2_X1   g0505(.A1(new_n588), .A2(G116), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT89), .ZN(new_n707));
  INV_X1    g0507(.A(new_n211), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G41), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n707), .A2(new_n252), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n710), .B1(new_n216), .B2(new_n709), .ZN(new_n711));
  XOR2_X1   g0511(.A(new_n711), .B(KEYINPUT28), .Z(new_n712));
  INV_X1    g0512(.A(G330), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n630), .A2(KEYINPUT90), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT90), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n634), .A2(new_n715), .A3(G179), .A4(new_n629), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n714), .A2(new_n716), .A3(new_n582), .A4(new_n510), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n718), .A2(KEYINPUT30), .A3(new_n538), .A4(new_n540), .ZN(new_n719));
  NOR3_X1   g0519(.A1(new_n637), .A2(new_n582), .A3(G179), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n720), .A2(new_n537), .A3(new_n483), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n538), .A2(new_n540), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n722), .B1(new_n723), .B2(new_n717), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n719), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n703), .ZN(new_n726));
  AOI21_X1  g0526(.A(KEYINPUT31), .B1(new_n725), .B2(new_n703), .ZN(new_n727));
  OAI21_X1  g0527(.A(KEYINPUT91), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n725), .A2(new_n703), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT31), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT91), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n703), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n728), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT92), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(new_n644), .B2(new_n703), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n690), .A2(new_n507), .A3(new_n694), .A4(new_n695), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n664), .A2(new_n558), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n541), .A2(new_n739), .A3(new_n542), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n670), .B(new_n740), .C1(new_n667), .C2(new_n603), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n742), .A2(KEYINPUT92), .A3(new_n686), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n737), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n713), .B1(new_n735), .B2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n679), .A2(new_n686), .ZN(new_n747));
  AOI21_X1  g0547(.A(KEYINPUT29), .B1(new_n747), .B2(KEYINPUT93), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n666), .B(new_n669), .C1(new_n667), .C2(new_n603), .ZN(new_n749));
  OAI21_X1  g0549(.A(KEYINPUT26), .B1(new_n670), .B2(new_n671), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n749), .A2(new_n750), .A3(new_n596), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n751), .A2(KEYINPUT94), .ZN(new_n752));
  AND2_X1   g0552(.A1(new_n596), .A2(new_n602), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n670), .A2(new_n507), .A3(new_n740), .A4(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n633), .B1(new_n688), .B2(new_n689), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n756), .B1(new_n751), .B2(KEYINPUT94), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n703), .B1(new_n752), .B2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT29), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT93), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n760), .B1(new_n747), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n748), .B1(new_n759), .B2(new_n762), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n746), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n712), .B1(new_n764), .B2(G1), .ZN(G364));
  INV_X1    g0565(.A(G13), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n252), .B1(new_n767), .B2(G45), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n709), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n698), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(G330), .B2(new_n697), .ZN(new_n772));
  INV_X1    g0572(.A(new_n770), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n218), .A2(G179), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n774), .A2(G190), .A3(G200), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n587), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n218), .A2(new_n334), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G200), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n277), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT32), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G190), .A2(G200), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n774), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G159), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n780), .A2(new_n215), .B1(new_n781), .B2(new_n785), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n776), .B(new_n786), .C1(new_n781), .C2(new_n785), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n777), .A2(G190), .A3(new_n332), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n271), .B1(new_n788), .B2(new_n202), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n778), .A2(G190), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n774), .A2(new_n277), .A3(G200), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n791), .A2(new_n203), .B1(new_n792), .B2(new_n459), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n277), .A2(G179), .A3(G200), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n218), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n789), .B(new_n793), .C1(G97), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n777), .A2(new_n782), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n798), .A2(KEYINPUT98), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(KEYINPUT98), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n787), .B(new_n797), .C1(new_n222), .C2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G303), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n269), .B1(new_n775), .B2(new_n803), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT99), .Z(new_n805));
  INV_X1    g0605(.A(G311), .ZN(new_n806));
  INV_X1    g0606(.A(G329), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n798), .A2(new_n806), .B1(new_n783), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n788), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n808), .B1(G322), .B2(new_n809), .ZN(new_n810));
  AOI22_X1  g0610(.A1(G294), .A2(new_n796), .B1(new_n779), .B2(G326), .ZN(new_n811));
  XNOR2_X1  g0611(.A(KEYINPUT33), .B(G317), .ZN(new_n812));
  INV_X1    g0612(.A(new_n792), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n790), .A2(new_n812), .B1(new_n813), .B2(G283), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n805), .A2(new_n810), .A3(new_n811), .A4(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT100), .ZN(new_n816));
  OR2_X1    g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n815), .A2(new_n816), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n802), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n217), .B1(G20), .B2(new_n307), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n773), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n766), .A2(new_n284), .A3(KEYINPUT97), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT97), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(G13), .B2(G33), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n826), .A2(G20), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(new_n820), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n208), .A2(KEYINPUT95), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n830), .A2(new_n211), .A3(new_n271), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n208), .A2(KEYINPUT95), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n831), .A2(new_n832), .B1(G116), .B2(new_n211), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT96), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n708), .A2(new_n271), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(new_n216), .B2(new_n472), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n472), .B2(new_n248), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n833), .A2(new_n834), .ZN(new_n840));
  AND3_X1   g0640(.A1(new_n835), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n827), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n821), .B1(new_n829), .B2(new_n841), .C1(new_n697), .C2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n772), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT101), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(G396));
  AOI22_X1  g0646(.A1(G137), .A2(new_n779), .B1(new_n809), .B2(G143), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n847), .B1(new_n290), .B2(new_n791), .C1(new_n801), .C2(new_n784), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT34), .Z(new_n849));
  OAI22_X1  g0649(.A1(new_n215), .A2(new_n775), .B1(new_n792), .B2(new_n203), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT103), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n850), .A2(new_n851), .ZN(new_n853));
  INV_X1    g0653(.A(G132), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n271), .B1(new_n783), .B2(new_n854), .C1(new_n795), .C2(new_n202), .ZN(new_n855));
  NOR4_X1   g0655(.A1(new_n849), .A2(new_n852), .A3(new_n853), .A4(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(G283), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n801), .A2(new_n607), .B1(new_n857), .B2(new_n791), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT102), .ZN(new_n859));
  INV_X1    g0659(.A(G294), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n269), .B1(new_n783), .B2(new_n806), .C1(new_n788), .C2(new_n860), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n780), .A2(new_n803), .B1(new_n556), .B2(new_n795), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n587), .A2(new_n792), .B1(new_n775), .B2(new_n459), .ZN(new_n863));
  NOR4_X1   g0663(.A1(new_n859), .A2(new_n861), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n820), .B1(new_n856), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n825), .A2(new_n820), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n773), .B1(new_n222), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n337), .A2(new_n703), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n321), .A2(new_n703), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n869), .B(KEYINPUT104), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n333), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n868), .B1(new_n871), .B2(new_n337), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n865), .B(new_n867), .C1(new_n872), .C2(new_n826), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n871), .A2(new_n647), .A3(new_n703), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n668), .A2(new_n672), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n596), .B1(new_n754), .B2(new_n755), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(KEYINPUT105), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT105), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n679), .A2(new_n879), .A3(new_n874), .ZN(new_n880));
  INV_X1    g0680(.A(new_n872), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n878), .A2(new_n880), .B1(new_n747), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n770), .B1(new_n746), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n746), .A2(new_n883), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n873), .B1(new_n885), .B2(new_n886), .ZN(G384));
  OR2_X1    g0687(.A1(new_n550), .A2(KEYINPUT35), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n550), .A2(KEYINPUT35), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n888), .A2(new_n889), .A3(G116), .A4(new_n219), .ZN(new_n890));
  XOR2_X1   g0690(.A(new_n890), .B(KEYINPUT36), .Z(new_n891));
  OAI211_X1 g0691(.A(new_n216), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n892));
  AOI211_X1 g0692(.A(new_n252), .B(G13), .C1(new_n892), .C2(new_n244), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n868), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n679), .A2(new_n879), .A3(new_n874), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n879), .B1(new_n679), .B2(new_n874), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(KEYINPUT106), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n878), .A2(new_n880), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT106), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n900), .A2(new_n901), .A3(new_n895), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n452), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n403), .B1(new_n413), .B2(new_n414), .ZN(new_n905));
  INV_X1    g0705(.A(new_n685), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n905), .B1(new_n446), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(KEYINPUT37), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n425), .A2(new_n438), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n425), .A2(new_n685), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT37), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n909), .A2(new_n910), .A3(new_n911), .A4(new_n452), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT107), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n905), .A2(new_n906), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n456), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n914), .B1(new_n456), .B2(new_n915), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT38), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI211_X1 g0720(.A(KEYINPUT38), .B(new_n913), .C1(new_n916), .C2(new_n917), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n397), .B1(new_n394), .B2(new_n395), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n391), .A2(KEYINPUT14), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n399), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n399), .A2(new_n703), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n925), .A2(new_n388), .A3(new_n926), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n399), .B(new_n703), .C1(new_n398), .C2(new_n389), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n903), .A2(new_n922), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n440), .A2(new_n447), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n906), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n909), .A2(new_n910), .A3(new_n452), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT37), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n912), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n456), .A2(new_n425), .A3(new_n685), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT38), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n921), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT39), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n398), .A2(new_n399), .A3(new_n686), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n941), .B(new_n943), .C1(new_n922), .C2(new_n940), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n930), .A2(new_n932), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n652), .B1(new_n763), .B2(new_n458), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n945), .B(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n733), .A2(KEYINPUT108), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT108), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n725), .A2(new_n949), .A3(KEYINPUT31), .A4(new_n703), .ZN(new_n950));
  AND3_X1   g0750(.A1(new_n948), .A2(new_n731), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n744), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n939), .A2(new_n952), .A3(new_n872), .A4(new_n929), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT40), .B1(new_n920), .B2(new_n921), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n929), .A2(new_n872), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n948), .A2(new_n731), .A3(new_n950), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(new_n737), .B2(new_n743), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n953), .A2(KEYINPUT40), .B1(new_n954), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n458), .B2(new_n957), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n954), .A2(new_n958), .ZN(new_n961));
  AOI21_X1  g0761(.A(KEYINPUT92), .B1(new_n742), .B2(new_n686), .ZN(new_n962));
  NOR4_X1   g0762(.A1(new_n738), .A2(new_n741), .A3(new_n736), .A4(new_n703), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n872), .B(new_n929), .C1(new_n964), .C2(new_n956), .ZN(new_n965));
  INV_X1    g0765(.A(new_n913), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n456), .A2(new_n915), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(KEYINPUT107), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n456), .A2(new_n914), .A3(new_n915), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n966), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n937), .B1(new_n970), .B2(KEYINPUT38), .ZN(new_n971));
  OAI21_X1  g0771(.A(KEYINPUT40), .B1(new_n965), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n961), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n973), .A2(new_n653), .A3(new_n952), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n960), .A2(new_n974), .A3(G330), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n947), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n252), .B2(new_n767), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n947), .A2(new_n975), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n894), .B1(new_n977), .B2(new_n978), .ZN(G367));
  OAI21_X1  g0779(.A(new_n828), .B1(new_n211), .B2(new_n314), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n239), .A2(new_n837), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n770), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n801), .A2(new_n215), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n791), .A2(new_n784), .B1(new_n792), .B2(new_n222), .ZN(new_n984));
  INV_X1    g0784(.A(G137), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n271), .B1(new_n783), .B2(new_n985), .C1(new_n788), .C2(new_n290), .ZN(new_n986));
  NOR3_X1   g0786(.A1(new_n983), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n775), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n779), .A2(G143), .B1(new_n988), .B2(G58), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n987), .B(new_n989), .C1(new_n203), .C2(new_n795), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(G116), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT46), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n269), .B1(new_n788), .B2(new_n803), .ZN(new_n993));
  INV_X1    g0793(.A(new_n783), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n993), .B1(G317), .B2(new_n994), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n992), .B(new_n995), .C1(new_n857), .C2(new_n801), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n790), .A2(G294), .B1(new_n813), .B2(G97), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(new_n459), .B2(new_n795), .C1(new_n806), .C2(new_n780), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n990), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT47), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n982), .B1(new_n1000), .B2(new_n820), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n601), .A2(new_n686), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT109), .Z(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n596), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n753), .B2(new_n1003), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n827), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1001), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n570), .B1(new_n739), .B2(new_n686), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n666), .A2(new_n703), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n704), .A2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT44), .Z(new_n1013));
  NOR2_X1   g0813(.A1(new_n704), .A2(new_n1011), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT45), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n699), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n699), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1013), .A2(new_n1018), .A3(new_n1015), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n702), .B1(new_n691), .B2(new_n701), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(new_n698), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n764), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n764), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n709), .B(KEYINPUT41), .Z(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n769), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(KEYINPUT114), .B1(new_n1018), .B2(new_n1011), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT110), .ZN(new_n1029));
  AOI21_X1  g0829(.A(KEYINPUT43), .B1(new_n1005), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n1029), .B2(new_n1005), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT113), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT114), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n699), .A2(new_n1035), .A3(new_n1010), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1028), .A2(new_n1034), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1034), .B1(new_n1028), .B2(new_n1036), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1004), .B(KEYINPUT43), .C1(new_n753), .C2(new_n1003), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT112), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1010), .A2(new_n524), .A3(new_n701), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1043), .A2(KEYINPUT42), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT111), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n670), .B1(new_n1008), .B2(new_n690), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n1043), .A2(KEYINPUT42), .B1(new_n1046), .B2(new_n686), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1042), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1040), .B(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1007), .B1(new_n1027), .B2(new_n1051), .ZN(G387));
  OR2_X1    g0852(.A1(new_n691), .A2(new_n842), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n707), .A2(new_n211), .A3(new_n271), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(G107), .B2(new_n211), .ZN(new_n1055));
  AOI211_X1 g0855(.A(G45), .B(new_n707), .C1(G68), .C2(G77), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1056), .A2(KEYINPUT115), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(KEYINPUT115), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n289), .A2(G50), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1059), .B(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1057), .A2(new_n1058), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n837), .B1(new_n236), .B2(G45), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1055), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n770), .B1(new_n1064), .B2(new_n829), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n798), .A2(new_n203), .B1(new_n783), .B2(new_n290), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n269), .B(new_n1066), .C1(G50), .C2(new_n809), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n988), .A2(G77), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n315), .A2(new_n796), .B1(new_n790), .B2(new_n312), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n779), .A2(G159), .B1(new_n813), .B2(G97), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n271), .B1(new_n994), .B2(G326), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n795), .A2(new_n857), .B1(new_n775), .B2(new_n860), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G311), .A2(new_n790), .B1(new_n809), .B2(G317), .ZN(new_n1074));
  INV_X1    g0874(.A(G322), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1074), .B1(new_n1075), .B2(new_n780), .C1(new_n801), .C2(new_n803), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT48), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1073), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n1077), .B2(new_n1076), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT49), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1072), .B1(new_n607), .B2(new_n792), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1071), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1065), .B1(new_n1083), .B2(new_n820), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n1022), .A2(new_n769), .B1(new_n1053), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1023), .A2(new_n709), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n764), .A2(new_n1022), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(G393));
  NAND3_X1  g0888(.A1(new_n1017), .A2(new_n769), .A3(new_n1019), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n828), .B1(new_n556), .B2(new_n211), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n243), .A2(new_n837), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n770), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n780), .A2(new_n290), .B1(new_n784), .B2(new_n788), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT51), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n792), .A2(new_n587), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n269), .B(new_n1095), .C1(G143), .C2(new_n994), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n796), .A2(G77), .B1(new_n988), .B2(G68), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1094), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n801), .A2(new_n289), .B1(new_n215), .B2(new_n791), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT117), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(G317), .A2(new_n779), .B1(new_n809), .B2(G311), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT52), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n791), .A2(new_n803), .B1(new_n792), .B2(new_n459), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n269), .B1(new_n783), .B2(new_n1075), .C1(new_n860), .C2(new_n798), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n795), .A2(new_n607), .B1(new_n775), .B2(new_n857), .ZN(new_n1105));
  OR3_X1    g0905(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n1098), .A2(new_n1100), .B1(new_n1102), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1092), .B1(new_n1107), .B2(new_n820), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n1010), .B2(new_n842), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1089), .A2(new_n1109), .ZN(new_n1110));
  OR2_X1    g0910(.A1(new_n1110), .A2(KEYINPUT118), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(KEYINPUT118), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n709), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1111), .A2(new_n1112), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(G390));
  AOI21_X1  g0918(.A(new_n868), .B1(new_n758), .B2(new_n872), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n929), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n939), .A2(new_n942), .ZN(new_n1122));
  OR2_X1    g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n728), .B(new_n734), .C1(new_n962), .C2(new_n963), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1124), .A2(G330), .A3(new_n872), .A4(new_n929), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n943), .B1(new_n903), .B2(new_n929), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n941), .B1(new_n922), .B2(new_n940), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1123), .B(new_n1125), .C1(new_n1126), .C2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n901), .B1(new_n900), .B2(new_n895), .ZN(new_n1131));
  AOI211_X1 g0931(.A(KEYINPUT106), .B(new_n868), .C1(new_n878), .C2(new_n880), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n929), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n942), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1130), .B1(new_n1134), .B2(new_n1127), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n955), .A2(new_n957), .A3(new_n713), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1129), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n952), .A2(new_n653), .A3(G330), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n652), .B(new_n1139), .C1(new_n763), .C2(new_n458), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT119), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n713), .B(new_n881), .C1(new_n744), .C2(new_n951), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1141), .B1(new_n1142), .B2(new_n929), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n1125), .A2(new_n1119), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n952), .A2(G330), .A3(new_n872), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1145), .A2(KEYINPUT119), .A3(new_n1120), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1143), .A2(new_n1144), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n929), .B1(new_n745), .B2(new_n872), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n903), .B1(new_n1148), .B2(new_n1136), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1140), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1138), .A2(new_n1151), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1129), .B(new_n1150), .C1(new_n1135), .C2(new_n1137), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1152), .A2(new_n709), .A3(new_n1153), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1129), .B(new_n769), .C1(new_n1135), .C2(new_n1137), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n866), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n770), .B1(new_n1156), .B2(new_n312), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n795), .A2(new_n222), .B1(new_n788), .B2(new_n607), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT121), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n271), .B(new_n776), .C1(G294), .C2(new_n994), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n556), .B2(new_n801), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n780), .A2(new_n857), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n791), .A2(new_n459), .B1(new_n792), .B2(new_n203), .ZN(new_n1163));
  NOR4_X1   g0963(.A1(new_n1159), .A2(new_n1161), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  OR2_X1    g0965(.A1(new_n1165), .A2(KEYINPUT122), .ZN(new_n1166));
  INV_X1    g0966(.A(G128), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n780), .A2(new_n1167), .B1(new_n854), .B2(new_n788), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT120), .ZN(new_n1169));
  INV_X1    g0969(.A(G125), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n271), .B1(new_n783), .B2(new_n1170), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n795), .A2(new_n784), .B1(new_n792), .B2(new_n215), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1171), .B(new_n1172), .C1(G137), .C2(new_n790), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(KEYINPUT54), .B(G143), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n801), .A2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n775), .A2(new_n290), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT53), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1169), .A2(new_n1173), .A3(new_n1175), .A4(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1165), .A2(KEYINPUT122), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1166), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1157), .B1(new_n1180), .B2(new_n820), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n1128), .B2(new_n826), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1155), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1154), .A2(new_n1184), .ZN(G378));
  NAND2_X1  g0985(.A1(new_n301), .A2(new_n685), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n651), .A2(new_n309), .A3(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n310), .A2(new_n301), .A3(new_n685), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1189));
  AND3_X1   g0989(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1189), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n973), .B2(G330), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n713), .B(new_n1192), .C1(new_n961), .C2(new_n972), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n945), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1192), .B1(new_n959), .B2(new_n713), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n973), .A2(G330), .A3(new_n1193), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n944), .A2(new_n932), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1197), .A2(new_n1198), .A3(new_n930), .A4(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1196), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n769), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1156), .A2(G50), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n792), .A2(new_n202), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n780), .A2(new_n607), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1204), .B(new_n1205), .C1(G97), .C2(new_n790), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n271), .A2(G41), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G283), .B2(new_n994), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n798), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n809), .A2(G107), .B1(new_n1209), .B2(new_n315), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n796), .A2(G68), .B1(new_n988), .B2(G77), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1206), .A2(new_n1208), .A3(new_n1210), .A4(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT58), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1207), .B(new_n215), .C1(G33), .C2(G41), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n1170), .A2(new_n780), .B1(new_n791), .B2(new_n854), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n809), .A2(G128), .B1(new_n1209), .B2(G137), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n775), .B2(new_n1174), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1217), .B(new_n1219), .C1(G150), .C2(new_n796), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(KEYINPUT59), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n813), .A2(G159), .ZN(new_n1223));
  AOI211_X1 g1023(.A(G33), .B(G41), .C1(new_n994), .C2(G124), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1221), .A2(KEYINPUT59), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1216), .B1(new_n1213), .B2(new_n1212), .C1(new_n1225), .C2(new_n1226), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n773), .B(new_n1203), .C1(new_n1227), .C2(new_n820), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n1193), .B2(new_n826), .ZN(new_n1229));
  AND2_X1   g1029(.A1(new_n1202), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1140), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1153), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT57), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n709), .ZN(new_n1236));
  AOI21_X1  g1036(.A(KEYINPUT57), .B1(new_n1232), .B2(new_n1201), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1230), .B1(new_n1236), .B2(new_n1237), .ZN(G375));
  AOI21_X1  g1038(.A(new_n768), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1239), .A2(KEYINPUT123), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n770), .B1(new_n1156), .B2(G68), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n854), .A2(new_n780), .B1(new_n791), .B2(new_n1174), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1204), .B(new_n1242), .C1(G50), .C2(new_n796), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n775), .A2(new_n784), .B1(new_n783), .B2(new_n1167), .ZN(new_n1244));
  XOR2_X1   g1044(.A(new_n1244), .B(KEYINPUT125), .Z(new_n1245));
  OAI21_X1  g1045(.A(new_n271), .B1(new_n788), .B2(new_n985), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(G150), .B2(new_n1209), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1243), .A2(new_n1245), .A3(new_n1247), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n801), .A2(new_n459), .B1(new_n607), .B2(new_n791), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(KEYINPUT124), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n780), .A2(new_n860), .B1(new_n775), .B2(new_n556), .ZN(new_n1251));
  OAI221_X1 g1051(.A(new_n269), .B1(new_n783), .B2(new_n803), .C1(new_n788), .C2(new_n857), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n795), .A2(new_n314), .B1(new_n792), .B2(new_n222), .ZN(new_n1253));
  OR3_X1    g1053(.A1(new_n1251), .A2(new_n1252), .A3(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1248), .B1(new_n1250), .B2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1241), .B1(new_n1255), .B2(new_n820), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n929), .B2(new_n826), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1257), .B1(new_n1239), .B2(KEYINPUT123), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1240), .A2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1147), .A2(new_n1149), .A3(new_n1140), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1151), .A2(new_n1026), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1259), .A2(new_n1261), .ZN(G381));
  INV_X1    g1062(.A(G384), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1117), .A2(new_n1263), .ZN(new_n1264));
  OR4_X1    g1064(.A1(G396), .A2(new_n1264), .A3(G387), .A4(G393), .ZN(new_n1265));
  OR4_X1    g1065(.A1(G378), .A2(new_n1265), .A3(G375), .A4(G381), .ZN(G407));
  AOI21_X1  g1066(.A(new_n1114), .B1(new_n1138), .B2(new_n1151), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1183), .B1(new_n1267), .B2(new_n1153), .ZN(new_n1268));
  INV_X1    g1068(.A(G343), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(G213), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1268), .A2(new_n1271), .ZN(new_n1272));
  OAI211_X1 g1072(.A(G407), .B(G213), .C1(G375), .C2(new_n1272), .ZN(G409));
  NOR2_X1   g1073(.A1(new_n1117), .A2(G387), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1117), .A2(G387), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(G393), .B(new_n845), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1275), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1277), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1276), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1279), .B1(new_n1280), .B2(new_n1274), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT61), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1278), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  OAI211_X1 g1083(.A(G378), .B(new_n1230), .C1(new_n1236), .C2(new_n1237), .ZN(new_n1284));
  AND3_X1   g1084(.A1(new_n1232), .A2(new_n1026), .A3(new_n1201), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1202), .A2(new_n1229), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1268), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1271), .B1(new_n1284), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT60), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1260), .B1(new_n1150), .B2(new_n1290), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1147), .A2(new_n1149), .A3(KEYINPUT60), .A4(new_n1140), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1291), .A2(new_n709), .A3(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1259), .A2(new_n1293), .A3(G384), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(G384), .B1(new_n1259), .B2(new_n1293), .ZN(new_n1296));
  OAI211_X1 g1096(.A(G2897), .B(new_n1271), .C1(new_n1295), .C2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1296), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1271), .A2(G2897), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1298), .A2(new_n1294), .A3(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1297), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1283), .B1(new_n1289), .B2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1284), .A2(new_n1287), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1304), .A2(KEYINPUT63), .A3(new_n1270), .A4(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT126), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1288), .A2(KEYINPUT126), .A3(KEYINPUT63), .A4(new_n1305), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1304), .A2(new_n1270), .A3(new_n1305), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT63), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1303), .A2(new_n1308), .A3(new_n1309), .A4(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT62), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1288), .A2(new_n1314), .A3(new_n1305), .ZN(new_n1315));
  XNOR2_X1  g1115(.A(KEYINPUT127), .B(KEYINPUT61), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1316), .B1(new_n1288), .B2(new_n1301), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1314), .B1(new_n1288), .B2(new_n1305), .ZN(new_n1318));
  NOR3_X1   g1118(.A1(new_n1315), .A2(new_n1317), .A3(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1278), .A2(new_n1281), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1320), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1313), .B1(new_n1319), .B2(new_n1321), .ZN(G405));
  NAND2_X1  g1122(.A1(G375), .A2(new_n1268), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1305), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1323), .A2(new_n1284), .A3(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1324), .B1(new_n1323), .B2(new_n1284), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  XNOR2_X1  g1128(.A(new_n1328), .B(new_n1321), .ZN(G402));
endmodule


