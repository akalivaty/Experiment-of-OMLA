//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 1 0 1 0 1 0 0 0 0 1 1 1 0 0 0 1 1 0 0 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n640, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n806,
    new_n807, new_n809, new_n810, new_n811, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  INV_X1    g004(.A(G8gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G29gat), .A2(G36gat), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT87), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT14), .ZN(new_n211));
  INV_X1    g010(.A(G29gat), .ZN(new_n212));
  INV_X1    g011(.A(G36gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n209), .A2(KEYINPUT87), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n208), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT15), .ZN(new_n218));
  OR2_X1    g017(.A1(G43gat), .A2(G50gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(G43gat), .A2(G50gat), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT88), .B(G43gat), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n218), .B(new_n220), .C1(new_n223), .C2(G50gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT89), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n214), .A2(new_n225), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n211), .A2(new_n212), .A3(new_n213), .A4(KEYINPUT89), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n226), .A2(new_n227), .A3(new_n209), .ZN(new_n228));
  INV_X1    g027(.A(new_n221), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n224), .A2(new_n228), .A3(new_n229), .A4(new_n208), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT17), .ZN(new_n231));
  AND3_X1   g030(.A1(new_n222), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n231), .B1(new_n222), .B2(new_n230), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n207), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G229gat), .A2(G233gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n205), .B(G8gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n222), .A2(new_n230), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n234), .A2(new_n235), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT18), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n234), .A2(KEYINPUT18), .A3(new_n235), .A4(new_n238), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n236), .B(new_n237), .ZN(new_n243));
  XOR2_X1   g042(.A(new_n235), .B(KEYINPUT13), .Z(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n241), .A2(new_n242), .A3(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G113gat), .B(G141gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(G197gat), .ZN(new_n248));
  XOR2_X1   g047(.A(KEYINPUT11), .B(G169gat), .Z(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n250), .B(KEYINPUT12), .Z(new_n251));
  NAND2_X1  g050(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n251), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n253), .A2(new_n241), .A3(new_n242), .A4(new_n245), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n257));
  XNOR2_X1  g056(.A(G197gat), .B(G204gat), .ZN(new_n258));
  INV_X1    g057(.A(G211gat), .ZN(new_n259));
  INV_X1    g058(.A(G218gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n258), .B1(KEYINPUT22), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G211gat), .B(G218gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n257), .B1(new_n264), .B2(KEYINPUT29), .ZN(new_n265));
  INV_X1    g064(.A(G141gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G148gat), .ZN(new_n267));
  INV_X1    g066(.A(G148gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(G141gat), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT2), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G155gat), .B(G162gat), .ZN(new_n271));
  OR3_X1    g070(.A1(new_n270), .A2(KEYINPUT74), .A3(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT74), .B1(new_n270), .B2(new_n271), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n271), .ZN(new_n275));
  INV_X1    g074(.A(G155gat), .ZN(new_n276));
  INV_X1    g075(.A(G162gat), .ZN(new_n277));
  OAI21_X1  g076(.A(KEYINPUT2), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT77), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI211_X1 g079(.A(KEYINPUT77), .B(KEYINPUT2), .C1(new_n276), .C2(new_n277), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n275), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT75), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT76), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n266), .A2(KEYINPUT75), .A3(G148gat), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n268), .A2(KEYINPUT76), .A3(G141gat), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n284), .A2(new_n286), .A3(new_n287), .A4(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n282), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n265), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n274), .A2(new_n257), .A3(new_n290), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT79), .ZN(new_n294));
  AOI22_X1  g093(.A1(new_n272), .A2(new_n273), .B1(new_n282), .B2(new_n289), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT79), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(new_n296), .A3(new_n257), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT29), .B1(new_n294), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n264), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n292), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT81), .ZN(new_n301));
  NAND2_X1  g100(.A1(G228gat), .A2(G233gat), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT81), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n303), .B(new_n292), .C1(new_n298), .C2(new_n299), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n301), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n300), .A2(KEYINPUT81), .A3(G228gat), .A4(G233gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G22gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n305), .A2(G22gat), .A3(new_n306), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G78gat), .B(G106gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(KEYINPUT31), .B(G50gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n312), .B(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(G22gat), .B1(new_n305), .B2(new_n306), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT82), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n311), .A2(new_n317), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n309), .A2(new_n316), .A3(new_n310), .A4(new_n314), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT83), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G1gat), .B(G29gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n323), .B(KEYINPUT0), .ZN(new_n324));
  XNOR2_X1  g123(.A(G57gat), .B(G85gat), .ZN(new_n325));
  XOR2_X1   g124(.A(new_n324), .B(new_n325), .Z(new_n326));
  XNOR2_X1  g125(.A(G113gat), .B(G120gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n327), .A2(KEYINPUT1), .ZN(new_n328));
  XNOR2_X1  g127(.A(G127gat), .B(G134gat), .ZN(new_n329));
  OR2_X1    g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT69), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT1), .ZN(new_n333));
  INV_X1    g132(.A(G120gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n334), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n332), .A2(new_n333), .A3(new_n329), .A4(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n330), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n295), .B(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(G225gat), .A2(G233gat), .ZN(new_n339));
  XOR2_X1   g138(.A(new_n339), .B(KEYINPUT80), .Z(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT5), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n337), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n345), .B1(new_n294), .B2(new_n297), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n291), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT78), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n348), .B1(new_n295), .B2(new_n257), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  OR3_X1    g149(.A1(new_n291), .A2(KEYINPUT4), .A3(new_n337), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n345), .A2(new_n295), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT4), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n346), .A2(new_n350), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n344), .B1(new_n341), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n354), .A2(KEYINPUT5), .A3(new_n341), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n326), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT6), .ZN(new_n359));
  INV_X1    g158(.A(new_n326), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n346), .A2(new_n350), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n351), .A2(new_n353), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n363), .A2(new_n340), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n360), .B(new_n356), .C1(new_n364), .C2(new_n344), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n358), .A2(new_n359), .A3(new_n365), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n355), .A2(new_n357), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n367), .A2(KEYINPUT6), .A3(new_n360), .ZN(new_n368));
  INV_X1    g167(.A(G226gat), .ZN(new_n369));
  INV_X1    g168(.A(G233gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(G169gat), .ZN(new_n372));
  INV_X1    g171(.A(G176gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n373), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n374), .B1(KEYINPUT26), .B2(new_n375), .ZN(new_n376));
  NOR3_X1   g175(.A1(new_n375), .A2(KEYINPUT68), .A3(KEYINPUT26), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT68), .ZN(new_n378));
  NOR2_X1   g177(.A1(G169gat), .A2(G176gat), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT26), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n376), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  XOR2_X1   g181(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n383));
  XNOR2_X1  g182(.A(KEYINPUT27), .B(G183gat), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n383), .B1(new_n385), .B2(G190gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(G183gat), .A2(G190gat), .ZN(new_n387));
  INV_X1    g186(.A(G190gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n384), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n382), .A2(new_n386), .A3(new_n387), .A4(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n392), .B(KEYINPUT64), .ZN(new_n393));
  INV_X1    g192(.A(G183gat), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n394), .A2(new_n388), .A3(KEYINPUT65), .ZN(new_n395));
  NAND3_X1  g194(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT65), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n397), .B1(G183gat), .B2(G190gat), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n393), .A2(new_n395), .A3(new_n396), .A4(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT66), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT23), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n375), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT66), .B1(new_n379), .B2(KEYINPUT23), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n374), .B1(KEYINPUT23), .B2(new_n379), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT25), .B1(new_n399), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n392), .B1(new_n394), .B2(new_n388), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n396), .ZN(new_n409));
  AND4_X1   g208(.A1(KEYINPUT25), .A2(new_n409), .A3(new_n404), .A4(new_n405), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n391), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT29), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n371), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n371), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n406), .A2(KEYINPUT25), .A3(new_n409), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n404), .A2(new_n405), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n395), .A2(new_n398), .A3(new_n396), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n416), .B1(new_n417), .B2(new_n393), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n415), .B1(new_n418), .B2(KEYINPUT25), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n414), .B1(new_n419), .B2(new_n391), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n264), .B1(new_n413), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n411), .A2(new_n371), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT29), .B1(new_n419), .B2(new_n391), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n422), .B(new_n299), .C1(new_n423), .C2(new_n371), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT73), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n421), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n413), .A2(new_n420), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n427), .A2(KEYINPUT73), .A3(new_n299), .ZN(new_n428));
  XNOR2_X1  g227(.A(G8gat), .B(G36gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(G64gat), .B(G92gat), .ZN(new_n430));
  XOR2_X1   g229(.A(new_n429), .B(new_n430), .Z(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n426), .A2(new_n428), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT30), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n426), .A2(new_n428), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n435), .A3(new_n431), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n431), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n437), .A2(KEYINPUT30), .A3(new_n433), .ZN(new_n438));
  AOI22_X1  g237(.A1(new_n366), .A2(new_n368), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n318), .A2(KEYINPUT83), .A3(new_n319), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n322), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n434), .B(new_n437), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT39), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT84), .B1(new_n363), .B2(new_n340), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT84), .ZN(new_n446));
  NOR3_X1   g245(.A1(new_n354), .A2(new_n446), .A3(new_n341), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n444), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n363), .A2(KEYINPUT84), .A3(new_n340), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n446), .B1(new_n354), .B2(new_n341), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n444), .B1(new_n338), .B2(new_n341), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n448), .A2(new_n326), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT40), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n448), .A2(KEYINPUT40), .A3(new_n326), .A4(new_n452), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n443), .A2(new_n455), .A3(new_n365), .A4(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n426), .A2(KEYINPUT37), .A3(new_n428), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT37), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT86), .B1(new_n435), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT86), .ZN(new_n461));
  AOI211_X1 g260(.A(new_n461), .B(KEYINPUT37), .C1(new_n426), .C2(new_n428), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n458), .B(new_n432), .C1(new_n460), .C2(new_n462), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n463), .A2(KEYINPUT38), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT85), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n424), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n466), .A2(new_n459), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n421), .A2(new_n424), .A3(new_n465), .ZN(new_n468));
  AOI21_X1  g267(.A(KEYINPUT38), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n432), .B(new_n469), .C1(new_n460), .C2(new_n462), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n470), .A2(new_n368), .A3(new_n366), .A4(new_n437), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n457), .B(new_n320), .C1(new_n464), .C2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT72), .ZN(new_n473));
  XOR2_X1   g272(.A(G15gat), .B(G43gat), .Z(new_n474));
  XNOR2_X1  g273(.A(G71gat), .B(G99gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(new_n475), .ZN(new_n476));
  AND2_X1   g275(.A1(G227gat), .A2(G233gat), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n411), .A2(new_n337), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n419), .A2(new_n345), .A3(new_n391), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n476), .B1(new_n481), .B2(KEYINPUT33), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT32), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n479), .A2(new_n480), .A3(new_n478), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT70), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(KEYINPUT34), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n482), .A2(new_n484), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n486), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT34), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n488), .B(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n490), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n493), .B1(new_n494), .B2(new_n485), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n473), .B1(new_n491), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n494), .A2(new_n485), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT72), .B1(new_n497), .B2(new_n489), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(KEYINPUT71), .B(KEYINPUT36), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT36), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n491), .A2(new_n495), .ZN(new_n503));
  OAI22_X1  g302(.A1(new_n499), .A2(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n442), .A2(new_n472), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n320), .A2(new_n439), .A3(new_n499), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT35), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n366), .A2(new_n368), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n436), .A2(new_n438), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n508), .A2(KEYINPUT35), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n503), .B1(new_n318), .B2(new_n319), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n506), .A2(new_n507), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n256), .B1(new_n505), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(new_n276), .ZN(new_n515));
  XNOR2_X1  g314(.A(G183gat), .B(G211gat), .ZN(new_n516));
  XOR2_X1   g315(.A(new_n515), .B(new_n516), .Z(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(G57gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(G64gat), .ZN(new_n520));
  INV_X1    g319(.A(G64gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(G57gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT91), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT91), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n520), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(G71gat), .A2(G78gat), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  OR2_X1    g327(.A1(new_n528), .A2(KEYINPUT9), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n524), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(G71gat), .A2(G78gat), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT90), .B1(new_n532), .B2(new_n527), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT90), .ZN(new_n534));
  NOR3_X1   g333(.A1(new_n528), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n530), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT92), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n520), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n522), .A2(KEYINPUT92), .ZN(new_n540));
  OAI221_X1 g339(.A(new_n529), .B1(new_n528), .B2(new_n531), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n542), .A2(KEYINPUT21), .ZN(new_n543));
  NAND2_X1  g342(.A1(G231gat), .A2(G233gat), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n543), .B(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(G127gat), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n236), .B1(KEYINPUT21), .B2(new_n542), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n546), .A2(new_n547), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n550), .B1(new_n548), .B2(new_n551), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n518), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n554), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n556), .A2(new_n552), .A3(new_n517), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G99gat), .A2(G106gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g359(.A1(G85gat), .A2(G92gat), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT7), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(G85gat), .ZN(new_n564));
  INV_X1    g363(.A(G92gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n560), .A2(new_n563), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G99gat), .B(G106gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT93), .ZN(new_n572));
  AOI22_X1  g371(.A1(KEYINPUT8), .A2(new_n559), .B1(new_n564), .B2(new_n565), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n573), .A2(new_n569), .A3(new_n563), .A4(new_n567), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n571), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n568), .A2(KEYINPUT93), .A3(new_n570), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT94), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT94), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n575), .A2(new_n579), .A3(new_n576), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n578), .B(new_n580), .C1(new_n232), .C2(new_n233), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n575), .A2(new_n579), .A3(new_n576), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n579), .B1(new_n575), .B2(new_n576), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n237), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n581), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(G190gat), .B(G218gat), .Z(new_n587));
  AND2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n586), .A2(new_n587), .ZN(new_n589));
  XNOR2_X1  g388(.A(G134gat), .B(G162gat), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  OR3_X1    g392(.A1(new_n588), .A2(new_n589), .A3(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n593), .B1(new_n588), .B2(new_n589), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n558), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(G230gat), .A2(G233gat), .ZN(new_n598));
  XOR2_X1   g397(.A(KEYINPUT95), .B(KEYINPUT10), .Z(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n537), .A2(new_n541), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(new_n577), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n571), .A2(new_n574), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n537), .A2(new_n541), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n600), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n537), .A2(new_n541), .A3(KEYINPUT10), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n606), .B1(new_n578), .B2(new_n580), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n598), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  AOI22_X1  g408(.A1(new_n537), .A2(new_n541), .B1(new_n575), .B2(new_n576), .ZN(new_n610));
  AND3_X1   g409(.A1(new_n537), .A2(new_n541), .A3(new_n603), .ZN(new_n611));
  NOR3_X1   g410(.A1(new_n610), .A2(new_n611), .A3(new_n598), .ZN(new_n612));
  XOR2_X1   g411(.A(G120gat), .B(G148gat), .Z(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT96), .ZN(new_n614));
  XNOR2_X1  g413(.A(G176gat), .B(G204gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  OR3_X1    g416(.A1(new_n609), .A2(new_n612), .A3(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n617), .B1(new_n609), .B2(new_n612), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n597), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n513), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n622), .A2(new_n508), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n623), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g423(.A1(new_n622), .A2(new_n509), .ZN(new_n625));
  XOR2_X1   g424(.A(KEYINPUT16), .B(G8gat), .Z(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n627), .B1(new_n206), .B2(new_n625), .ZN(new_n628));
  MUX2_X1   g427(.A(new_n627), .B(new_n628), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g428(.A(G15gat), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n622), .A2(new_n630), .A3(new_n504), .ZN(new_n631));
  INV_X1    g430(.A(new_n499), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n630), .B1(new_n622), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT97), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n631), .B1(new_n635), .B2(new_n636), .ZN(G1326gat));
  NAND2_X1  g436(.A1(new_n322), .A2(new_n441), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(KEYINPUT43), .B(G22gat), .Z(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(G1327gat));
  INV_X1    g440(.A(new_n558), .ZN(new_n642));
  INV_X1    g441(.A(new_n620), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n644), .A2(new_n596), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n513), .A2(new_n645), .ZN(new_n646));
  NOR3_X1   g445(.A1(new_n646), .A2(G29gat), .A3(new_n508), .ZN(new_n647));
  XNOR2_X1  g446(.A(KEYINPUT98), .B(KEYINPUT45), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n472), .A2(new_n504), .ZN(new_n650));
  AND3_X1   g449(.A1(new_n318), .A2(KEYINPUT83), .A3(new_n319), .ZN(new_n651));
  AOI21_X1  g450(.A(KEYINPUT83), .B1(new_n318), .B2(new_n319), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n651), .A2(new_n652), .A3(new_n439), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n512), .B1(new_n650), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n596), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(KEYINPUT44), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT99), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT44), .B1(new_n654), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT100), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n596), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n594), .A2(KEYINPUT100), .A3(new_n595), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n664), .B1(new_n658), .B2(KEYINPUT44), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n657), .B1(new_n659), .B2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n644), .A2(new_n256), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(G29gat), .B1(new_n669), .B2(new_n508), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n649), .A2(new_n670), .ZN(G1328gat));
  NOR3_X1   g470(.A1(new_n646), .A2(G36gat), .A3(new_n509), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT46), .ZN(new_n673));
  OAI21_X1  g472(.A(G36gat), .B1(new_n669), .B2(new_n509), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(G1329gat));
  OAI21_X1  g474(.A(new_n223), .B1(new_n669), .B2(new_n504), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT47), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n677), .A2(KEYINPUT101), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n646), .A2(new_n223), .A3(new_n632), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n679), .B1(KEYINPUT101), .B2(new_n677), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n676), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n678), .B1(new_n676), .B2(new_n680), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(G1330gat));
  NOR2_X1   g482(.A1(new_n669), .A2(new_n320), .ZN(new_n684));
  INV_X1    g483(.A(G50gat), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n651), .A2(new_n652), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n513), .A2(new_n685), .A3(new_n687), .A4(new_n645), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT48), .ZN(new_n689));
  INV_X1    g488(.A(new_n688), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n667), .A2(new_n687), .A3(new_n668), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n690), .B1(new_n691), .B2(G50gat), .ZN(new_n692));
  OAI22_X1  g491(.A1(new_n686), .A2(new_n689), .B1(new_n692), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g492(.A1(new_n597), .A2(new_n255), .A3(new_n643), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n654), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(new_n508), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(new_n519), .ZN(G1332gat));
  NOR2_X1   g496(.A1(new_n695), .A2(new_n509), .ZN(new_n698));
  NOR2_X1   g497(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n699));
  AND2_X1   g498(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(new_n698), .B2(new_n699), .ZN(G1333gat));
  OR3_X1    g501(.A1(new_n695), .A2(G71gat), .A3(new_n632), .ZN(new_n703));
  OAI21_X1  g502(.A(G71gat), .B1(new_n695), .B2(new_n504), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g505(.A1(new_n695), .A2(new_n638), .ZN(new_n707));
  XOR2_X1   g506(.A(KEYINPUT102), .B(G78gat), .Z(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(G1335gat));
  NOR2_X1   g508(.A1(new_n558), .A2(new_n255), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(new_n643), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n654), .A2(new_n658), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n666), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n713), .B1(new_n717), .B2(new_n657), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(G85gat), .B1(new_n719), .B2(new_n508), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n596), .B1(new_n505), .B2(new_n512), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n711), .B1(new_n721), .B2(KEYINPUT103), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT103), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n656), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT51), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n722), .A2(new_n724), .A3(KEYINPUT51), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n508), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n731), .A2(new_n564), .A3(new_n620), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n720), .B1(new_n730), .B2(new_n732), .ZN(G1336gat));
  NAND3_X1  g532(.A1(new_n443), .A2(new_n565), .A3(new_n620), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT105), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n722), .A2(new_n724), .A3(KEYINPUT51), .ZN(new_n736));
  AOI21_X1  g535(.A(KEYINPUT51), .B1(new_n722), .B2(new_n724), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT104), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n721), .A2(new_n715), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n443), .B(new_n712), .C1(new_n716), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(G92gat), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n738), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n740), .A2(new_n744), .A3(KEYINPUT52), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT52), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n738), .B(new_n743), .C1(new_n739), .C2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(G1337gat));
  OAI21_X1  g547(.A(G99gat), .B1(new_n719), .B2(new_n504), .ZN(new_n749));
  OR3_X1    g548(.A1(new_n632), .A2(G99gat), .A3(new_n643), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n730), .B2(new_n750), .ZN(G1338gat));
  INV_X1    g550(.A(new_n320), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n667), .A2(new_n752), .A3(new_n712), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT107), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT107), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n667), .A2(new_n755), .A3(new_n752), .A4(new_n712), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n754), .A2(G106gat), .A3(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(G106gat), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n752), .A2(new_n758), .A3(new_n620), .ZN(new_n759));
  XOR2_X1   g558(.A(new_n759), .B(KEYINPUT106), .Z(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT53), .B1(new_n729), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n757), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n758), .B1(new_n718), .B2(new_n687), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n760), .B1(new_n727), .B2(new_n728), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT53), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n763), .A2(new_n766), .ZN(G1339gat));
  NOR2_X1   g566(.A1(new_n243), .A2(new_n244), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n235), .B1(new_n234), .B2(new_n238), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n250), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n254), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT54), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n616), .B1(new_n609), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n599), .B1(new_n610), .B2(new_n611), .ZN(new_n774));
  OAI211_X1 g573(.A(KEYINPUT10), .B(new_n542), .C1(new_n582), .C2(new_n583), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n772), .B1(new_n776), .B2(new_n598), .ZN(new_n777));
  INV_X1    g576(.A(new_n598), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n774), .A2(new_n775), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT108), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  AND4_X1   g579(.A1(KEYINPUT108), .A2(new_n608), .A3(KEYINPUT54), .A4(new_n779), .ZN(new_n781));
  OAI211_X1 g580(.A(KEYINPUT55), .B(new_n773), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n782), .A2(new_n618), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n773), .B1(new_n780), .B2(new_n781), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n663), .A2(new_n771), .A3(new_n783), .A4(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n783), .A2(new_n255), .A3(new_n786), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n620), .A2(new_n771), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n663), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n642), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  AND4_X1   g591(.A1(new_n256), .A2(new_n558), .A3(new_n596), .A4(new_n643), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n687), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n508), .A2(new_n443), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n795), .A2(new_n499), .A3(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(G113gat), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n797), .A2(new_n798), .A3(new_n256), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n508), .B1(new_n792), .B2(new_n794), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n800), .A2(new_n511), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n509), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n255), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n799), .B1(new_n804), .B2(new_n798), .ZN(G1340gat));
  NOR3_X1   g604(.A1(new_n797), .A2(new_n334), .A3(new_n643), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n803), .A2(new_n620), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n806), .B1(new_n807), .B2(new_n334), .ZN(G1341gat));
  OAI21_X1  g607(.A(G127gat), .B1(new_n797), .B2(new_n642), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n558), .A2(new_n547), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n809), .B1(new_n802), .B2(new_n810), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(KEYINPUT109), .ZN(G1342gat));
  NOR3_X1   g611(.A1(new_n443), .A2(G134gat), .A3(new_n596), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n801), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n814), .A2(KEYINPUT56), .ZN(new_n815));
  XOR2_X1   g614(.A(new_n815), .B(KEYINPUT110), .Z(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(KEYINPUT56), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(KEYINPUT111), .ZN(new_n818));
  OAI21_X1  g617(.A(G134gat), .B1(new_n797), .B2(new_n596), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n816), .A2(new_n818), .A3(new_n819), .ZN(G1343gat));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n638), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n823));
  INV_X1    g622(.A(new_n790), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n784), .A2(KEYINPUT112), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT112), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n826), .B(new_n773), .C1(new_n780), .C2(new_n781), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n825), .A2(new_n785), .A3(new_n827), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n782), .A2(new_n255), .A3(new_n618), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n824), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n787), .B1(new_n830), .B2(new_n655), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n831), .A2(new_n642), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n822), .B(new_n823), .C1(new_n832), .C2(new_n793), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n687), .A2(KEYINPUT57), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n793), .B1(new_n831), .B2(new_n642), .ZN(new_n835));
  OAI21_X1  g634(.A(KEYINPUT113), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n320), .B1(new_n792), .B2(new_n794), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n833), .B(new_n836), .C1(KEYINPUT57), .C2(new_n837), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n504), .A2(new_n796), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n838), .A2(new_n255), .A3(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT114), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n840), .A2(new_n841), .A3(G141gat), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n841), .B1(new_n840), .B2(G141gat), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n504), .A2(new_n752), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n800), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n845), .A2(new_n266), .A3(new_n255), .A4(new_n509), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n842), .A2(new_n843), .A3(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT58), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n850), .B1(G141gat), .B2(new_n840), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT115), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI211_X1 g652(.A(KEYINPUT115), .B(new_n850), .C1(new_n840), .C2(G141gat), .ZN(new_n854));
  OAI22_X1  g653(.A1(new_n848), .A2(new_n849), .B1(new_n853), .B2(new_n854), .ZN(G1344gat));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n783), .A2(new_n655), .A3(new_n771), .A4(new_n786), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n857), .B1(new_n830), .B2(new_n655), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n793), .B1(new_n858), .B2(new_n642), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT118), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n687), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AOI211_X1 g660(.A(KEYINPUT118), .B(new_n793), .C1(new_n858), .C2(new_n642), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n821), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(KEYINPUT119), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n865), .B(new_n821), .C1(new_n861), .C2(new_n862), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n789), .A2(new_n790), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n664), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n558), .B1(new_n868), .B2(new_n787), .ZN(new_n869));
  OAI211_X1 g668(.A(KEYINPUT57), .B(new_n752), .C1(new_n869), .C2(new_n793), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT117), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n837), .A2(KEYINPUT117), .A3(KEYINPUT57), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n864), .A2(new_n866), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n839), .A2(new_n620), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n268), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n856), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI22_X1  g679(.A1(new_n863), .A2(KEYINPUT119), .B1(new_n872), .B2(new_n873), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n876), .B1(new_n881), .B2(new_n866), .ZN(new_n882));
  OAI211_X1 g681(.A(KEYINPUT120), .B(KEYINPUT59), .C1(new_n882), .C2(new_n268), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n838), .A2(new_n839), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n879), .B(G148gat), .C1(new_n884), .C2(new_n643), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n880), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n845), .A2(new_n509), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n887), .A2(G148gat), .A3(new_n643), .ZN(new_n888));
  XOR2_X1   g687(.A(new_n888), .B(KEYINPUT116), .Z(new_n889));
  NAND2_X1  g688(.A1(new_n886), .A2(new_n889), .ZN(G1345gat));
  OAI21_X1  g689(.A(G155gat), .B1(new_n884), .B2(new_n642), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n558), .A2(new_n276), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n891), .B1(new_n887), .B2(new_n892), .ZN(G1346gat));
  OAI21_X1  g692(.A(G162gat), .B1(new_n884), .B2(new_n664), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n845), .A2(new_n277), .A3(new_n509), .A4(new_n655), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1347gat));
  AOI21_X1  g695(.A(new_n731), .B1(new_n792), .B2(new_n794), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n511), .A2(new_n443), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(G169gat), .B1(new_n900), .B2(new_n255), .ZN(new_n901));
  AND4_X1   g700(.A1(new_n508), .A2(new_n795), .A3(new_n443), .A4(new_n499), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n256), .A2(new_n372), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(G1348gat));
  NAND3_X1  g703(.A1(new_n900), .A2(new_n373), .A3(new_n620), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n902), .A2(new_n620), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n905), .B1(new_n906), .B2(new_n373), .ZN(G1349gat));
  NAND3_X1  g706(.A1(new_n900), .A2(new_n384), .A3(new_n558), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n902), .A2(new_n558), .ZN(new_n909));
  OAI211_X1 g708(.A(KEYINPUT121), .B(new_n908), .C1(new_n909), .C2(new_n394), .ZN(new_n910));
  XOR2_X1   g709(.A(KEYINPUT122), .B(KEYINPUT60), .Z(new_n911));
  XNOR2_X1  g710(.A(new_n910), .B(new_n911), .ZN(G1350gat));
  AOI21_X1  g711(.A(new_n388), .B1(new_n902), .B2(new_n655), .ZN(new_n913));
  XOR2_X1   g712(.A(new_n913), .B(KEYINPUT61), .Z(new_n914));
  NAND3_X1  g713(.A1(new_n900), .A2(new_n388), .A3(new_n663), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1351gat));
  NAND3_X1  g715(.A1(new_n897), .A2(new_n443), .A3(new_n844), .ZN(new_n917));
  XOR2_X1   g716(.A(new_n917), .B(KEYINPUT123), .Z(new_n918));
  AOI21_X1  g717(.A(G197gat), .B1(new_n918), .B2(new_n255), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n504), .A2(new_n508), .A3(new_n443), .ZN(new_n920));
  XOR2_X1   g719(.A(new_n920), .B(KEYINPUT124), .Z(new_n921));
  AOI21_X1  g720(.A(new_n921), .B1(new_n881), .B2(new_n866), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n255), .A2(G197gat), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(G1352gat));
  NOR3_X1   g723(.A1(new_n917), .A2(G204gat), .A3(new_n643), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT62), .ZN(new_n926));
  AOI211_X1 g725(.A(new_n643), .B(new_n921), .C1(new_n881), .C2(new_n866), .ZN(new_n927));
  INV_X1    g726(.A(G204gat), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT125), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI211_X1 g730(.A(KEYINPUT125), .B(new_n926), .C1(new_n927), .C2(new_n928), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1353gat));
  NAND3_X1  g732(.A1(new_n918), .A2(new_n259), .A3(new_n558), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n922), .A2(new_n558), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n935), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n936));
  AOI21_X1  g735(.A(KEYINPUT63), .B1(new_n935), .B2(G211gat), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(G1354gat));
  NAND3_X1  g737(.A1(new_n918), .A2(new_n260), .A3(new_n663), .ZN(new_n939));
  AOI211_X1 g738(.A(new_n596), .B(new_n921), .C1(new_n881), .C2(new_n866), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n940), .B2(new_n260), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(KEYINPUT126), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n943));
  OAI211_X1 g742(.A(new_n943), .B(new_n939), .C1(new_n940), .C2(new_n260), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n942), .A2(new_n944), .ZN(G1355gat));
endmodule


