

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X1 U325 ( .A(KEYINPUT46), .B(KEYINPUT106), .ZN(n372) );
  XNOR2_X1 U326 ( .A(n373), .B(n372), .ZN(n390) );
  XNOR2_X1 U327 ( .A(n420), .B(KEYINPUT48), .ZN(n421) );
  XNOR2_X1 U328 ( .A(n422), .B(n421), .ZN(n545) );
  NOR2_X1 U329 ( .A1(n529), .A2(n453), .ZN(n564) );
  XNOR2_X1 U330 ( .A(n371), .B(n370), .ZN(n571) );
  XNOR2_X1 U331 ( .A(n454), .B(G190GAT), .ZN(n455) );
  XNOR2_X1 U332 ( .A(n456), .B(n455), .ZN(G1351GAT) );
  XOR2_X1 U333 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n294) );
  XNOR2_X1 U334 ( .A(KEYINPUT19), .B(G183GAT), .ZN(n293) );
  XNOR2_X1 U335 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U336 ( .A(G169GAT), .B(n295), .Z(n334) );
  XOR2_X1 U337 ( .A(KEYINPUT81), .B(KEYINPUT20), .Z(n297) );
  XNOR2_X1 U338 ( .A(KEYINPUT80), .B(KEYINPUT79), .ZN(n296) );
  XNOR2_X1 U339 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U340 ( .A(G99GAT), .B(G190GAT), .Z(n299) );
  XOR2_X1 U341 ( .A(G43GAT), .B(G134GAT), .Z(n402) );
  XOR2_X1 U342 ( .A(G120GAT), .B(G71GAT), .Z(n352) );
  XNOR2_X1 U343 ( .A(n402), .B(n352), .ZN(n298) );
  XNOR2_X1 U344 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U345 ( .A(n301), .B(n300), .Z(n303) );
  NAND2_X1 U346 ( .A1(G227GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U347 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U348 ( .A(n304), .B(G176GAT), .Z(n307) );
  XNOR2_X1 U349 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n305) );
  XNOR2_X1 U350 ( .A(n305), .B(G127GAT), .ZN(n436) );
  XNOR2_X1 U351 ( .A(G15GAT), .B(n436), .ZN(n306) );
  XNOR2_X1 U352 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U353 ( .A(n334), .B(n308), .Z(n519) );
  INV_X1 U354 ( .A(n519), .ZN(n529) );
  XOR2_X1 U355 ( .A(KEYINPUT22), .B(KEYINPUT82), .Z(n314) );
  XOR2_X1 U356 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n310) );
  XNOR2_X1 U357 ( .A(G106GAT), .B(G204GAT), .ZN(n309) );
  XNOR2_X1 U358 ( .A(n310), .B(n309), .ZN(n312) );
  XNOR2_X1 U359 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n311) );
  XNOR2_X1 U360 ( .A(n311), .B(KEYINPUT2), .ZN(n435) );
  XNOR2_X1 U361 ( .A(n312), .B(n435), .ZN(n313) );
  XNOR2_X1 U362 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U363 ( .A(G50GAT), .B(G162GAT), .Z(n408) );
  XOR2_X1 U364 ( .A(G148GAT), .B(G78GAT), .Z(n344) );
  XOR2_X1 U365 ( .A(n408), .B(n344), .Z(n316) );
  NAND2_X1 U366 ( .A1(G228GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U367 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U368 ( .A(n318), .B(n317), .Z(n324) );
  XOR2_X1 U369 ( .A(G141GAT), .B(G22GAT), .Z(n356) );
  XNOR2_X1 U370 ( .A(G211GAT), .B(KEYINPUT83), .ZN(n319) );
  XNOR2_X1 U371 ( .A(n319), .B(KEYINPUT21), .ZN(n320) );
  XOR2_X1 U372 ( .A(n320), .B(KEYINPUT84), .Z(n322) );
  XNOR2_X1 U373 ( .A(G197GAT), .B(G218GAT), .ZN(n321) );
  XNOR2_X1 U374 ( .A(n322), .B(n321), .ZN(n333) );
  XNOR2_X1 U375 ( .A(n356), .B(n333), .ZN(n323) );
  XNOR2_X1 U376 ( .A(n324), .B(n323), .ZN(n462) );
  XNOR2_X1 U377 ( .A(KEYINPUT54), .B(KEYINPUT117), .ZN(n426) );
  XOR2_X1 U378 ( .A(G36GAT), .B(G190GAT), .Z(n405) );
  XOR2_X1 U379 ( .A(G64GAT), .B(G92GAT), .Z(n326) );
  XNOR2_X1 U380 ( .A(G176GAT), .B(G204GAT), .ZN(n325) );
  XNOR2_X1 U381 ( .A(n326), .B(n325), .ZN(n349) );
  XOR2_X1 U382 ( .A(n405), .B(n349), .Z(n328) );
  NAND2_X1 U383 ( .A1(G226GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U384 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U385 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n330) );
  XNOR2_X1 U386 ( .A(G8GAT), .B(KEYINPUT90), .ZN(n329) );
  XNOR2_X1 U387 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U388 ( .A(n332), .B(n331), .Z(n336) );
  XNOR2_X1 U389 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U390 ( .A(n336), .B(n335), .Z(n504) );
  XOR2_X1 U391 ( .A(KEYINPUT116), .B(n504), .Z(n423) );
  INV_X1 U392 ( .A(KEYINPUT33), .ZN(n337) );
  NAND2_X1 U393 ( .A1(n337), .A2(KEYINPUT31), .ZN(n340) );
  INV_X1 U394 ( .A(KEYINPUT31), .ZN(n338) );
  NAND2_X1 U395 ( .A1(n338), .A2(KEYINPUT33), .ZN(n339) );
  NAND2_X1 U396 ( .A1(n340), .A2(n339), .ZN(n342) );
  XNOR2_X1 U397 ( .A(KEYINPUT72), .B(KEYINPUT32), .ZN(n341) );
  XNOR2_X1 U398 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U399 ( .A(n344), .B(n343), .Z(n346) );
  NAND2_X1 U400 ( .A1(G230GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U401 ( .A(n346), .B(n345), .ZN(n351) );
  XOR2_X1 U402 ( .A(KEYINPUT71), .B(G85GAT), .Z(n348) );
  XNOR2_X1 U403 ( .A(G99GAT), .B(G106GAT), .ZN(n347) );
  XNOR2_X1 U404 ( .A(n348), .B(n347), .ZN(n407) );
  XOR2_X1 U405 ( .A(n407), .B(n349), .Z(n350) );
  XNOR2_X1 U406 ( .A(n351), .B(n350), .ZN(n354) );
  XOR2_X1 U407 ( .A(G57GAT), .B(KEYINPUT13), .Z(n375) );
  XNOR2_X1 U408 ( .A(n352), .B(n375), .ZN(n353) );
  XNOR2_X1 U409 ( .A(n354), .B(n353), .ZN(n574) );
  XNOR2_X1 U410 ( .A(KEYINPUT41), .B(n574), .ZN(n498) );
  XNOR2_X1 U411 ( .A(G15GAT), .B(G1GAT), .ZN(n355) );
  XNOR2_X1 U412 ( .A(n355), .B(G8GAT), .ZN(n374) );
  XOR2_X1 U413 ( .A(n374), .B(n356), .Z(n358) );
  XNOR2_X1 U414 ( .A(G36GAT), .B(G50GAT), .ZN(n357) );
  XNOR2_X1 U415 ( .A(n358), .B(n357), .ZN(n363) );
  XNOR2_X1 U416 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n359) );
  XNOR2_X1 U417 ( .A(n359), .B(KEYINPUT8), .ZN(n394) );
  XOR2_X1 U418 ( .A(n394), .B(KEYINPUT69), .Z(n361) );
  NAND2_X1 U419 ( .A1(G229GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U420 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U421 ( .A(n363), .B(n362), .Z(n371) );
  XOR2_X1 U422 ( .A(G113GAT), .B(G197GAT), .Z(n365) );
  XNOR2_X1 U423 ( .A(G169GAT), .B(G43GAT), .ZN(n364) );
  XNOR2_X1 U424 ( .A(n365), .B(n364), .ZN(n369) );
  XOR2_X1 U425 ( .A(KEYINPUT70), .B(KEYINPUT30), .Z(n367) );
  XNOR2_X1 U426 ( .A(KEYINPUT68), .B(KEYINPUT29), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U428 ( .A(n369), .B(n368), .ZN(n370) );
  NAND2_X1 U429 ( .A1(n498), .A2(n571), .ZN(n373) );
  XOR2_X1 U430 ( .A(n375), .B(n374), .Z(n377) );
  NAND2_X1 U431 ( .A1(G231GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U432 ( .A(n377), .B(n376), .ZN(n381) );
  XOR2_X1 U433 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n379) );
  XNOR2_X1 U434 ( .A(KEYINPUT12), .B(KEYINPUT78), .ZN(n378) );
  XNOR2_X1 U435 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U436 ( .A(n381), .B(n380), .Z(n389) );
  XOR2_X1 U437 ( .A(G78GAT), .B(G155GAT), .Z(n383) );
  XNOR2_X1 U438 ( .A(G22GAT), .B(G211GAT), .ZN(n382) );
  XNOR2_X1 U439 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U440 ( .A(G64GAT), .B(G71GAT), .Z(n385) );
  XNOR2_X1 U441 ( .A(G183GAT), .B(G127GAT), .ZN(n384) );
  XNOR2_X1 U442 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U443 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U444 ( .A(n389), .B(n388), .Z(n580) );
  INV_X1 U445 ( .A(n580), .ZN(n483) );
  NAND2_X1 U446 ( .A1(n390), .A2(n483), .ZN(n391) );
  XNOR2_X1 U447 ( .A(n391), .B(KEYINPUT107), .ZN(n413) );
  XOR2_X1 U448 ( .A(KEYINPUT76), .B(KEYINPUT9), .Z(n393) );
  XNOR2_X1 U449 ( .A(KEYINPUT77), .B(KEYINPUT75), .ZN(n392) );
  XNOR2_X1 U450 ( .A(n393), .B(n392), .ZN(n398) );
  XOR2_X1 U451 ( .A(n394), .B(KEYINPUT66), .Z(n396) );
  NAND2_X1 U452 ( .A1(G232GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U453 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U454 ( .A(n398), .B(n397), .Z(n412) );
  XOR2_X1 U455 ( .A(KEYINPUT67), .B(KEYINPUT10), .Z(n400) );
  XNOR2_X1 U456 ( .A(G92GAT), .B(KEYINPUT74), .ZN(n399) );
  XNOR2_X1 U457 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U458 ( .A(n401), .B(KEYINPUT11), .Z(n404) );
  XNOR2_X1 U459 ( .A(n402), .B(G218GAT), .ZN(n403) );
  XNOR2_X1 U460 ( .A(n404), .B(n403), .ZN(n406) );
  XOR2_X1 U461 ( .A(n406), .B(n405), .Z(n410) );
  XNOR2_X1 U462 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U463 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U464 ( .A(n412), .B(n411), .ZN(n554) );
  INV_X1 U465 ( .A(n554), .ZN(n470) );
  NAND2_X1 U466 ( .A1(n413), .A2(n470), .ZN(n414) );
  XNOR2_X1 U467 ( .A(n414), .B(KEYINPUT47), .ZN(n419) );
  XOR2_X1 U468 ( .A(KEYINPUT36), .B(n554), .Z(n583) );
  NOR2_X1 U469 ( .A1(n483), .A2(n583), .ZN(n415) );
  XNOR2_X1 U470 ( .A(n415), .B(KEYINPUT45), .ZN(n416) );
  NAND2_X1 U471 ( .A1(n416), .A2(n574), .ZN(n417) );
  NOR2_X1 U472 ( .A1(n417), .A2(n571), .ZN(n418) );
  NOR2_X1 U473 ( .A1(n419), .A2(n418), .ZN(n422) );
  XOR2_X1 U474 ( .A(KEYINPUT64), .B(KEYINPUT108), .Z(n420) );
  NAND2_X1 U475 ( .A1(n423), .A2(n545), .ZN(n424) );
  XNOR2_X1 U476 ( .A(n424), .B(KEYINPUT118), .ZN(n425) );
  XNOR2_X1 U477 ( .A(n426), .B(n425), .ZN(n449) );
  XOR2_X1 U478 ( .A(G57GAT), .B(KEYINPUT85), .Z(n428) );
  XNOR2_X1 U479 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n427) );
  XNOR2_X1 U480 ( .A(n428), .B(n427), .ZN(n440) );
  XOR2_X1 U481 ( .A(KEYINPUT87), .B(KEYINPUT86), .Z(n430) );
  XNOR2_X1 U482 ( .A(G120GAT), .B(KEYINPUT6), .ZN(n429) );
  XNOR2_X1 U483 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U484 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n432) );
  XNOR2_X1 U485 ( .A(KEYINPUT89), .B(KEYINPUT88), .ZN(n431) );
  XNOR2_X1 U486 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U487 ( .A(n434), .B(n433), .Z(n438) );
  XNOR2_X1 U488 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U489 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U490 ( .A(n440), .B(n439), .ZN(n448) );
  NAND2_X1 U491 ( .A1(G225GAT), .A2(G233GAT), .ZN(n446) );
  XOR2_X1 U492 ( .A(G148GAT), .B(G162GAT), .Z(n442) );
  XNOR2_X1 U493 ( .A(G141GAT), .B(G134GAT), .ZN(n441) );
  XNOR2_X1 U494 ( .A(n442), .B(n441), .ZN(n444) );
  XOR2_X1 U495 ( .A(G29GAT), .B(G85GAT), .Z(n443) );
  XNOR2_X1 U496 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U497 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U498 ( .A(n448), .B(n447), .Z(n546) );
  INV_X1 U499 ( .A(n546), .ZN(n500) );
  NAND2_X1 U500 ( .A1(n449), .A2(n500), .ZN(n450) );
  XNOR2_X1 U501 ( .A(KEYINPUT65), .B(n450), .ZN(n570) );
  NAND2_X1 U502 ( .A1(n462), .A2(n570), .ZN(n452) );
  INV_X1 U503 ( .A(KEYINPUT55), .ZN(n451) );
  XNOR2_X1 U504 ( .A(n452), .B(n451), .ZN(n453) );
  NAND2_X1 U505 ( .A1(n564), .A2(n554), .ZN(n456) );
  XOR2_X1 U506 ( .A(KEYINPUT58), .B(KEYINPUT121), .Z(n454) );
  NAND2_X1 U507 ( .A1(n574), .A2(n571), .ZN(n457) );
  XNOR2_X1 U508 ( .A(n457), .B(KEYINPUT73), .ZN(n488) );
  XOR2_X1 U509 ( .A(n504), .B(KEYINPUT27), .Z(n465) );
  XOR2_X1 U510 ( .A(n462), .B(KEYINPUT28), .Z(n522) );
  INV_X1 U511 ( .A(n522), .ZN(n508) );
  NAND2_X1 U512 ( .A1(n465), .A2(n508), .ZN(n458) );
  NOR2_X1 U513 ( .A1(n500), .A2(n458), .ZN(n527) );
  NAND2_X1 U514 ( .A1(n527), .A2(n529), .ZN(n459) );
  XOR2_X1 U515 ( .A(KEYINPUT93), .B(n459), .Z(n469) );
  INV_X1 U516 ( .A(n504), .ZN(n516) );
  NAND2_X1 U517 ( .A1(n519), .A2(n516), .ZN(n460) );
  NAND2_X1 U518 ( .A1(n462), .A2(n460), .ZN(n461) );
  XOR2_X1 U519 ( .A(KEYINPUT25), .B(n461), .Z(n466) );
  XNOR2_X1 U520 ( .A(KEYINPUT26), .B(KEYINPUT94), .ZN(n464) );
  NOR2_X1 U521 ( .A1(n519), .A2(n462), .ZN(n463) );
  XNOR2_X1 U522 ( .A(n464), .B(n463), .ZN(n569) );
  NAND2_X1 U523 ( .A1(n569), .A2(n465), .ZN(n548) );
  NAND2_X1 U524 ( .A1(n466), .A2(n548), .ZN(n467) );
  NAND2_X1 U525 ( .A1(n500), .A2(n467), .ZN(n468) );
  NAND2_X1 U526 ( .A1(n469), .A2(n468), .ZN(n482) );
  NAND2_X1 U527 ( .A1(n470), .A2(n580), .ZN(n471) );
  XOR2_X1 U528 ( .A(KEYINPUT16), .B(n471), .Z(n472) );
  AND2_X1 U529 ( .A1(n482), .A2(n472), .ZN(n499) );
  NAND2_X1 U530 ( .A1(n488), .A2(n499), .ZN(n479) );
  NOR2_X1 U531 ( .A1(n500), .A2(n479), .ZN(n474) );
  XNOR2_X1 U532 ( .A(KEYINPUT95), .B(KEYINPUT34), .ZN(n473) );
  XNOR2_X1 U533 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U534 ( .A(G1GAT), .B(n475), .ZN(G1324GAT) );
  NOR2_X1 U535 ( .A1(n504), .A2(n479), .ZN(n476) );
  XOR2_X1 U536 ( .A(G8GAT), .B(n476), .Z(G1325GAT) );
  NOR2_X1 U537 ( .A1(n529), .A2(n479), .ZN(n478) );
  XNOR2_X1 U538 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n478), .B(n477), .ZN(G1326GAT) );
  NOR2_X1 U540 ( .A1(n508), .A2(n479), .ZN(n480) );
  XOR2_X1 U541 ( .A(KEYINPUT96), .B(n480), .Z(n481) );
  XNOR2_X1 U542 ( .A(G22GAT), .B(n481), .ZN(G1327GAT) );
  NAND2_X1 U543 ( .A1(n483), .A2(n482), .ZN(n484) );
  NOR2_X1 U544 ( .A1(n583), .A2(n484), .ZN(n486) );
  XNOR2_X1 U545 ( .A(KEYINPUT37), .B(KEYINPUT97), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U547 ( .A(KEYINPUT98), .B(n487), .ZN(n512) );
  NAND2_X1 U548 ( .A1(n488), .A2(n512), .ZN(n489) );
  XNOR2_X1 U549 ( .A(KEYINPUT38), .B(n489), .ZN(n496) );
  NOR2_X1 U550 ( .A1(n496), .A2(n500), .ZN(n491) );
  XNOR2_X1 U551 ( .A(KEYINPUT99), .B(KEYINPUT39), .ZN(n490) );
  XNOR2_X1 U552 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U553 ( .A(G29GAT), .B(n492), .Z(G1328GAT) );
  NOR2_X1 U554 ( .A1(n496), .A2(n504), .ZN(n493) );
  XOR2_X1 U555 ( .A(G36GAT), .B(n493), .Z(G1329GAT) );
  NOR2_X1 U556 ( .A1(n496), .A2(n529), .ZN(n494) );
  XOR2_X1 U557 ( .A(KEYINPUT40), .B(n494), .Z(n495) );
  XNOR2_X1 U558 ( .A(G43GAT), .B(n495), .ZN(G1330GAT) );
  NOR2_X1 U559 ( .A1(n496), .A2(n508), .ZN(n497) );
  XOR2_X1 U560 ( .A(G50GAT), .B(n497), .Z(G1331GAT) );
  INV_X1 U561 ( .A(n498), .ZN(n532) );
  NOR2_X1 U562 ( .A1(n571), .A2(n532), .ZN(n511) );
  NAND2_X1 U563 ( .A1(n511), .A2(n499), .ZN(n507) );
  NOR2_X1 U564 ( .A1(n500), .A2(n507), .ZN(n502) );
  XNOR2_X1 U565 ( .A(KEYINPUT42), .B(KEYINPUT100), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U567 ( .A(G57GAT), .B(n503), .Z(G1332GAT) );
  NOR2_X1 U568 ( .A1(n504), .A2(n507), .ZN(n505) );
  XOR2_X1 U569 ( .A(G64GAT), .B(n505), .Z(G1333GAT) );
  NOR2_X1 U570 ( .A1(n529), .A2(n507), .ZN(n506) );
  XOR2_X1 U571 ( .A(G71GAT), .B(n506), .Z(G1334GAT) );
  NOR2_X1 U572 ( .A1(n508), .A2(n507), .ZN(n510) );
  XNOR2_X1 U573 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n510), .B(n509), .ZN(G1335GAT) );
  NAND2_X1 U575 ( .A1(n512), .A2(n511), .ZN(n513) );
  XNOR2_X1 U576 ( .A(n513), .B(KEYINPUT101), .ZN(n523) );
  NAND2_X1 U577 ( .A1(n546), .A2(n523), .ZN(n514) );
  XNOR2_X1 U578 ( .A(KEYINPUT102), .B(n514), .ZN(n515) );
  XNOR2_X1 U579 ( .A(G85GAT), .B(n515), .ZN(G1336GAT) );
  XOR2_X1 U580 ( .A(G92GAT), .B(KEYINPUT103), .Z(n518) );
  NAND2_X1 U581 ( .A1(n523), .A2(n516), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n518), .B(n517), .ZN(G1337GAT) );
  NAND2_X1 U583 ( .A1(n523), .A2(n519), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n520), .B(KEYINPUT104), .ZN(n521) );
  XNOR2_X1 U585 ( .A(G99GAT), .B(n521), .ZN(G1338GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT44), .B(KEYINPUT105), .Z(n525) );
  NAND2_X1 U587 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  NAND2_X1 U590 ( .A1(n545), .A2(n527), .ZN(n528) );
  NOR2_X1 U591 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U592 ( .A(KEYINPUT109), .B(n530), .Z(n540) );
  NAND2_X1 U593 ( .A1(n571), .A2(n540), .ZN(n531) );
  XNOR2_X1 U594 ( .A(G113GAT), .B(n531), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT111), .B(KEYINPUT49), .Z(n534) );
  NAND2_X1 U596 ( .A1(n540), .A2(n498), .ZN(n533) );
  XNOR2_X1 U597 ( .A(n534), .B(n533), .ZN(n536) );
  XOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT110), .Z(n535) );
  XNOR2_X1 U599 ( .A(n536), .B(n535), .ZN(G1341GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT112), .B(KEYINPUT50), .Z(n538) );
  NAND2_X1 U601 ( .A1(n540), .A2(n580), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U603 ( .A(G127GAT), .B(n539), .Z(G1342GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n542) );
  NAND2_X1 U605 ( .A1(n540), .A2(n554), .ZN(n541) );
  XNOR2_X1 U606 ( .A(n542), .B(n541), .ZN(n544) );
  XOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT113), .Z(n543) );
  XNOR2_X1 U608 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  NAND2_X1 U609 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U610 ( .A1(n548), .A2(n547), .ZN(n555) );
  NAND2_X1 U611 ( .A1(n571), .A2(n555), .ZN(n549) );
  XNOR2_X1 U612 ( .A(G141GAT), .B(n549), .ZN(G1344GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n551) );
  NAND2_X1 U614 ( .A1(n555), .A2(n498), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(n552), .ZN(G1345GAT) );
  NAND2_X1 U617 ( .A1(n580), .A2(n555), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n553), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U619 ( .A(G162GAT), .B(KEYINPUT115), .Z(n557) );
  NAND2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n557), .B(n556), .ZN(G1347GAT) );
  NAND2_X1 U622 ( .A1(n564), .A2(n571), .ZN(n558) );
  XNOR2_X1 U623 ( .A(G169GAT), .B(n558), .ZN(G1348GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT57), .B(KEYINPUT120), .Z(n560) );
  XNOR2_X1 U625 ( .A(G176GAT), .B(KEYINPUT119), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U627 ( .A(KEYINPUT56), .B(n561), .Z(n563) );
  NAND2_X1 U628 ( .A1(n564), .A2(n498), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1349GAT) );
  NAND2_X1 U630 ( .A1(n580), .A2(n564), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT123), .Z(n567) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT122), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(n568) );
  XOR2_X1 U635 ( .A(KEYINPUT59), .B(n568), .Z(n573) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n582) );
  INV_X1 U637 ( .A(n582), .ZN(n579) );
  NAND2_X1 U638 ( .A1(n579), .A2(n571), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  NOR2_X1 U640 ( .A1(n582), .A2(n574), .ZN(n578) );
  XOR2_X1 U641 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n576) );
  XNOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n575) );
  XNOR2_X1 U643 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n585) );
  XNOR2_X1 U648 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(G218GAT), .B(n586), .Z(G1355GAT) );
endmodule

