//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036;
  INV_X1    g000(.A(KEYINPUT31), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT65), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  NAND2_X1  g004(.A1(KEYINPUT65), .A2(G146), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(G143), .A3(new_n191), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n189), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  AND2_X1   g008(.A1(KEYINPUT0), .A2(G128), .ZN(new_n195));
  AND3_X1   g009(.A1(new_n192), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G128), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  AND2_X1   g012(.A1(KEYINPUT65), .A2(G146), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT65), .A2(G146), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n198), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n189), .A2(G143), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n197), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n196), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(G137), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT11), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(G137), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G137), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT67), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT67), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G137), .ZN(new_n213));
  AND2_X1   g027(.A1(KEYINPUT11), .A2(G134), .ZN(new_n214));
  AND3_X1   g028(.A1(new_n211), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NOR3_X1   g029(.A1(new_n209), .A2(G131), .A3(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G131), .ZN(new_n217));
  AND2_X1   g031(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n218));
  NOR2_X1   g032(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n208), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n206), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n211), .A2(new_n213), .A3(new_n214), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n217), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n204), .B1(new_n216), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G128), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n192), .A2(new_n194), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n226), .B1(new_n192), .B2(KEYINPUT1), .ZN(new_n229));
  INV_X1    g043(.A(new_n202), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT65), .B(G146), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(new_n198), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n228), .B1(new_n229), .B2(new_n232), .ZN(new_n233));
  OR2_X1    g047(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n234));
  NAND2_X1  g048(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n235));
  AOI22_X1  g049(.A1(new_n234), .A2(new_n235), .B1(new_n205), .B2(G137), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n217), .B(new_n223), .C1(new_n236), .C2(new_n206), .ZN(new_n237));
  AOI21_X1  g051(.A(G134), .B1(new_n211), .B2(new_n213), .ZN(new_n238));
  OAI21_X1  g052(.A(G131), .B1(new_n238), .B2(new_n206), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n233), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(G116), .B(G119), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT2), .B(G113), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n241), .B(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n225), .A2(new_n240), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT71), .ZN(new_n245));
  AND2_X1   g059(.A1(KEYINPUT69), .A2(G953), .ZN(new_n246));
  NOR2_X1   g060(.A1(KEYINPUT69), .A2(G953), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G237), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(G210), .A3(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT26), .B(G101), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n248), .A2(new_n251), .A3(G210), .A4(new_n249), .ZN(new_n255));
  AND3_X1   g069(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n254), .B1(new_n253), .B2(new_n255), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n244), .A2(new_n245), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n245), .B1(new_n244), .B2(new_n258), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n225), .A2(new_n240), .A3(KEYINPUT30), .ZN(new_n262));
  INV_X1    g076(.A(new_n243), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NOR3_X1   g078(.A1(new_n199), .A2(new_n200), .A3(new_n198), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT1), .ZN(new_n266));
  OAI21_X1  g080(.A(G128), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n201), .A2(new_n202), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n199), .A2(new_n200), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n193), .B1(new_n269), .B2(G143), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n267), .A2(new_n268), .B1(new_n270), .B2(new_n227), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n237), .A2(new_n239), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT68), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT68), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n233), .A2(new_n274), .A3(new_n237), .A4(new_n239), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n273), .A2(new_n275), .A3(new_n225), .ZN(new_n276));
  XOR2_X1   g090(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n264), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n187), .B1(new_n261), .B2(new_n279), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n225), .A2(new_n240), .A3(new_n243), .ZN(new_n281));
  INV_X1    g095(.A(new_n258), .ZN(new_n282));
  OAI21_X1  g096(.A(KEYINPUT71), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n244), .A2(new_n245), .A3(new_n258), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n276), .A2(new_n278), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n237), .A2(new_n239), .ZN(new_n287));
  OAI21_X1  g101(.A(G131), .B1(new_n209), .B2(new_n215), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n237), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n233), .A2(new_n287), .B1(new_n289), .B2(new_n204), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n243), .B1(new_n290), .B2(KEYINPUT30), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n285), .A2(new_n292), .A3(KEYINPUT31), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n271), .A2(new_n272), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n192), .A2(new_n194), .A3(new_n195), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n296), .B1(new_n232), .B2(new_n197), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n297), .B1(new_n237), .B2(new_n288), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n294), .B1(new_n295), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n225), .A2(new_n240), .A3(KEYINPUT72), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(new_n243), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT28), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n281), .B1(new_n276), .B2(new_n263), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n303), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  AOI22_X1  g119(.A1(new_n280), .A2(new_n293), .B1(new_n305), .B2(new_n282), .ZN(new_n306));
  NOR2_X1   g120(.A1(G472), .A2(G902), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT32), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n276), .A2(new_n263), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n302), .B1(new_n310), .B2(new_n244), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n225), .A2(new_n240), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n263), .B1(new_n312), .B2(new_n294), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT28), .B1(new_n313), .B2(new_n300), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n282), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  NOR3_X1   g129(.A1(new_n261), .A2(new_n279), .A3(new_n187), .ZN(new_n316));
  AOI21_X1  g130(.A(KEYINPUT31), .B1(new_n285), .B2(new_n292), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT32), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(new_n319), .A3(new_n307), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n309), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n312), .A2(new_n263), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n302), .B1(new_n323), .B2(new_n244), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n314), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n282), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(G902), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT73), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n281), .B1(new_n286), .B2(new_n291), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n329), .B1(new_n330), .B2(new_n258), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n240), .A2(KEYINPUT68), .B1(new_n289), .B2(new_n204), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n277), .B1(new_n332), .B2(new_n275), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n244), .B1(new_n333), .B2(new_n264), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(KEYINPUT73), .A3(new_n282), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n303), .B(new_n258), .C1(new_n302), .C2(new_n304), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n326), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n328), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G472), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n321), .A2(new_n322), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n322), .B1(new_n321), .B2(new_n340), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(G214), .B1(G237), .B2(G902), .ZN(new_n344));
  XOR2_X1   g158(.A(new_n344), .B(KEYINPUT91), .Z(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(G110), .B(G122), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n347), .B(KEYINPUT8), .ZN(new_n348));
  INV_X1    g162(.A(G107), .ZN(new_n349));
  OAI21_X1  g163(.A(KEYINPUT88), .B1(new_n349), .B2(G104), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT88), .ZN(new_n351));
  INV_X1    g165(.A(G104), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(new_n352), .A3(G107), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n350), .B(new_n353), .C1(new_n352), .C2(G107), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G101), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT87), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(new_n349), .A3(G104), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(KEYINPUT3), .ZN(new_n358));
  INV_X1    g172(.A(G101), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT3), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n356), .A2(new_n360), .A3(new_n349), .A4(G104), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n352), .A2(G107), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n358), .A2(new_n359), .A3(new_n361), .A4(new_n362), .ZN(new_n363));
  AND2_X1   g177(.A1(new_n355), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G119), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G116), .ZN(new_n366));
  INV_X1    g180(.A(G116), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G119), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  OR2_X1    g183(.A1(new_n369), .A2(new_n242), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT92), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n371), .B1(new_n366), .B2(KEYINPUT5), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT5), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n373), .A2(new_n365), .A3(KEYINPUT92), .A4(G116), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n372), .A2(G113), .A3(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n369), .A2(new_n373), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n370), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n348), .B1(new_n364), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT93), .B1(new_n369), .B2(new_n373), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT93), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n241), .A2(new_n380), .A3(KEYINPUT5), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n374), .A2(G113), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n379), .A2(new_n381), .A3(new_n382), .A4(new_n372), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT94), .B1(new_n383), .B2(new_n370), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n355), .A2(new_n363), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n383), .A2(KEYINPUT94), .A3(new_n370), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n378), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n297), .A2(G125), .ZN(new_n389));
  INV_X1    g203(.A(G125), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n390), .B(new_n228), .C1(new_n229), .C2(new_n232), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G224), .ZN(new_n393));
  OAI21_X1  g207(.A(KEYINPUT7), .B1(new_n393), .B2(G953), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n394), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n389), .A2(new_n391), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n388), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n358), .A2(new_n361), .A3(new_n362), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G101), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(KEYINPUT4), .A3(new_n363), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT4), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n400), .A2(new_n403), .A3(G101), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n402), .A2(new_n263), .A3(new_n404), .ZN(new_n405));
  OR2_X1    g219(.A1(new_n377), .A2(new_n385), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n406), .A3(new_n347), .ZN(new_n407));
  AOI21_X1  g221(.A(G902), .B1(new_n399), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n405), .A2(new_n406), .ZN(new_n409));
  INV_X1    g223(.A(new_n347), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(KEYINPUT6), .A3(new_n407), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT6), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n409), .A2(new_n413), .A3(new_n410), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n393), .A2(G953), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n392), .B(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n412), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(G210), .B1(G237), .B2(G902), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n408), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n418), .B1(new_n408), .B2(new_n417), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n346), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT95), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n408), .A2(new_n417), .ZN(new_n423));
  INV_X1    g237(.A(new_n418), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n408), .A2(new_n417), .A3(new_n418), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT95), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n428), .A3(new_n346), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n422), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(G116), .B(G122), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT14), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n367), .A2(KEYINPUT14), .A3(G122), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(G107), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n431), .A2(KEYINPUT102), .A3(new_n349), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n431), .A2(new_n349), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT102), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n435), .A2(new_n436), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n198), .A2(G128), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n226), .A2(G143), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n205), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n441), .A2(new_n442), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G134), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n444), .A2(KEYINPUT101), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n444), .A2(new_n446), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT101), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n440), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n441), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n453), .A2(KEYINPUT13), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n442), .B1(new_n453), .B2(KEYINPUT13), .ZN(new_n455));
  OAI21_X1  g269(.A(G134), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n431), .B(new_n349), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n444), .A3(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT9), .B(G234), .ZN(new_n459));
  INV_X1    g273(.A(G217), .ZN(new_n460));
  NOR3_X1   g274(.A1(new_n459), .A2(new_n460), .A3(G953), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n452), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n461), .ZN(new_n463));
  INV_X1    g277(.A(new_n458), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n463), .B1(new_n451), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(G902), .ZN(new_n467));
  INV_X1    g281(.A(G478), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(KEYINPUT15), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n466), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n470), .B1(new_n466), .B2(new_n467), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(G952), .ZN(new_n475));
  AOI211_X1 g289(.A(G953), .B(new_n475), .C1(G234), .C2(G237), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  AOI211_X1 g291(.A(new_n467), .B(new_n248), .C1(G234), .C2(G237), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(KEYINPUT21), .B(G898), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n480), .B(KEYINPUT103), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n477), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n474), .A2(new_n482), .ZN(new_n483));
  OR2_X1    g297(.A1(KEYINPUT69), .A2(G953), .ZN(new_n484));
  NAND2_X1  g298(.A1(KEYINPUT69), .A2(G953), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n484), .A2(G214), .A3(new_n249), .A4(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n198), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n248), .A2(G143), .A3(G214), .A4(new_n249), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n217), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT17), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n487), .A2(new_n488), .A3(new_n217), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT99), .ZN(new_n494));
  INV_X1    g308(.A(G140), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(G125), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n390), .A2(G140), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT78), .ZN(new_n498));
  OR3_X1    g312(.A1(new_n390), .A2(KEYINPUT78), .A3(G140), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n499), .A3(KEYINPUT16), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT16), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n500), .A2(new_n189), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n189), .B1(new_n500), .B2(new_n502), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n494), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n489), .A2(KEYINPUT17), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n500), .A2(new_n502), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(G146), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(KEYINPUT99), .A3(new_n503), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n493), .A2(new_n506), .A3(new_n507), .A4(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(G113), .B(G122), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT98), .B(G104), .ZN(new_n513));
  XOR2_X1   g327(.A(new_n512), .B(new_n513), .Z(new_n514));
  NAND2_X1  g328(.A1(new_n487), .A2(new_n488), .ZN(new_n515));
  NAND2_X1  g329(.A1(KEYINPUT96), .A2(KEYINPUT18), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n515), .A2(G131), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n498), .A2(new_n499), .A3(G146), .ZN(new_n519));
  XNOR2_X1  g333(.A(G125), .B(G140), .ZN(new_n520));
  AND3_X1   g334(.A1(new_n269), .A2(new_n520), .A3(KEYINPUT80), .ZN(new_n521));
  AOI21_X1  g335(.A(KEYINPUT80), .B1(new_n269), .B2(new_n520), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n519), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n487), .B(new_n488), .C1(new_n217), .C2(new_n516), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n518), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n511), .A2(new_n514), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n514), .B1(new_n511), .B2(new_n525), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n467), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(G475), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT20), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT19), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n532), .B1(new_n498), .B2(new_n499), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n520), .A2(KEYINPUT19), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n269), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n487), .A2(new_n488), .A3(new_n217), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n509), .B(new_n535), .C1(new_n536), .C2(new_n489), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n525), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT97), .ZN(new_n539));
  INV_X1    g353(.A(new_n514), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT97), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n537), .A2(new_n525), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n526), .ZN(new_n544));
  NOR2_X1   g358(.A1(G475), .A2(G902), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n531), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n545), .ZN(new_n547));
  AOI211_X1 g361(.A(KEYINPUT20), .B(new_n547), .C1(new_n543), .C2(new_n526), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n530), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT100), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT100), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n530), .B(new_n551), .C1(new_n546), .C2(new_n548), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n483), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(G469), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n248), .A2(G227), .ZN(new_n555));
  XOR2_X1   g369(.A(new_n555), .B(KEYINPUT86), .Z(new_n556));
  XNOR2_X1  g370(.A(G110), .B(G140), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n556), .B(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT10), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n226), .B1(new_n202), .B2(KEYINPUT1), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n228), .B1(new_n270), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n559), .B1(new_n562), .B2(new_n385), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n402), .A2(new_n204), .A3(new_n404), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n364), .A2(KEYINPUT10), .A3(new_n233), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n289), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n289), .A2(KEYINPUT89), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT89), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n288), .A2(new_n569), .A3(new_n237), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n571), .A2(new_n564), .A3(new_n563), .A4(new_n565), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n558), .B1(new_n567), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT90), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT12), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n216), .A2(new_n224), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n271), .A2(new_n385), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n364), .A2(new_n561), .ZN(new_n578));
  AOI211_X1 g392(.A(new_n575), .B(new_n576), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n578), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT12), .B1(new_n580), .B2(new_n289), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n572), .A2(new_n558), .ZN(new_n583));
  OAI22_X1  g397(.A1(new_n573), .A2(new_n574), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AOI211_X1 g398(.A(KEYINPUT90), .B(new_n558), .C1(new_n567), .C2(new_n572), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n554), .B(new_n467), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n558), .ZN(new_n587));
  INV_X1    g401(.A(new_n572), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n587), .B1(new_n582), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n567), .A2(new_n572), .A3(new_n558), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n589), .A2(G469), .A3(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n554), .A2(new_n467), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n586), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(G221), .B1(new_n459), .B2(G902), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n430), .A2(new_n553), .A3(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT82), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n226), .A2(G119), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n365), .A2(G128), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT76), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n602), .B1(new_n600), .B2(new_n601), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g419(.A(KEYINPUT24), .B(G110), .Z(new_n606));
  INV_X1    g420(.A(KEYINPUT77), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n600), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT23), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n609), .B1(new_n365), .B2(G128), .ZN(new_n610));
  NOR2_X1   g424(.A1(KEYINPUT77), .A2(KEYINPUT23), .ZN(new_n611));
  OAI22_X1  g425(.A1(new_n608), .A2(new_n610), .B1(new_n600), .B2(new_n611), .ZN(new_n612));
  OAI22_X1  g426(.A1(new_n605), .A2(new_n606), .B1(G110), .B2(new_n612), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n613), .B(new_n509), .C1(new_n522), .C2(new_n521), .ZN(new_n614));
  AOI22_X1  g428(.A1(new_n605), .A2(new_n606), .B1(new_n612), .B2(G110), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT79), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n615), .B(new_n616), .C1(new_n504), .C2(new_n505), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n509), .A2(new_n503), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n616), .B1(new_n619), .B2(new_n615), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n614), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n248), .A2(G221), .A3(G234), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT22), .B(G137), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n599), .B1(new_n621), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n619), .A2(new_n615), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(KEYINPUT79), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n617), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n629), .A2(KEYINPUT82), .A3(new_n614), .A4(new_n624), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n621), .A2(KEYINPUT81), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT81), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n633), .B(new_n614), .C1(new_n618), .C2(new_n620), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n632), .A2(new_n634), .A3(new_n625), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n631), .A2(new_n467), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(KEYINPUT25), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT25), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n631), .A2(new_n635), .A3(new_n638), .A4(new_n467), .ZN(new_n639));
  INV_X1    g453(.A(G234), .ZN(new_n640));
  OAI21_X1  g454(.A(G217), .B1(new_n640), .B2(G902), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT75), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n637), .A2(new_n639), .A3(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT83), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n642), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n646), .B1(new_n636), .B2(KEYINPUT25), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(KEYINPUT83), .A3(new_n639), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n642), .A2(G902), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n631), .A2(new_n635), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT84), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n645), .A2(new_n648), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(KEYINPUT85), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT85), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n645), .A2(new_n654), .A3(new_n648), .A4(new_n651), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n343), .A2(new_n598), .A3(new_n653), .A4(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G101), .ZN(G3));
  AND2_X1   g471(.A1(new_n653), .A2(new_n655), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n468), .A2(new_n467), .ZN(new_n659));
  INV_X1    g473(.A(new_n466), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n660), .A2(G902), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n659), .B1(new_n661), .B2(new_n468), .ZN(new_n662));
  OR2_X1    g476(.A1(new_n466), .A2(KEYINPUT33), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n466), .A2(KEYINPUT33), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n663), .A2(G478), .A3(new_n664), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n550), .A2(new_n552), .A3(new_n666), .ZN(new_n667));
  OAI211_X1 g481(.A(new_n346), .B(new_n482), .C1(new_n419), .C2(new_n420), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(G472), .B1(new_n306), .B2(G902), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n670), .B1(new_n308), .B2(new_n306), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n671), .A2(new_n596), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n658), .A2(new_n669), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT34), .B(G104), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G6));
  INV_X1    g489(.A(new_n473), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n471), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n677), .B(new_n530), .C1(new_n546), .C2(new_n548), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n345), .B1(new_n425), .B2(new_n426), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n679), .A2(KEYINPUT104), .A3(new_n680), .A4(new_n482), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT104), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n682), .B1(new_n668), .B2(new_n678), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n658), .A2(new_n672), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT35), .B(G107), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G9));
  NAND2_X1  g501(.A1(new_n550), .A2(new_n552), .ZN(new_n688));
  INV_X1    g502(.A(new_n483), .ZN(new_n689));
  AND4_X1   g503(.A1(new_n688), .A2(new_n689), .A3(new_n595), .A4(new_n594), .ZN(new_n690));
  INV_X1    g504(.A(new_n671), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n632), .A2(new_n634), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n692), .A2(KEYINPUT36), .A3(new_n625), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n625), .A2(KEYINPUT36), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n694), .B1(new_n632), .B2(new_n634), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n649), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n645), .A2(new_n648), .A3(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n690), .A2(new_n430), .A3(new_n691), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(KEYINPUT105), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT37), .B(G110), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G12));
  AND4_X1   g515(.A1(KEYINPUT83), .A2(new_n637), .A3(new_n639), .A4(new_n642), .ZN(new_n702));
  AOI21_X1  g516(.A(KEYINPUT83), .B1(new_n647), .B2(new_n639), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n421), .B1(new_n704), .B2(new_n696), .ZN(new_n705));
  INV_X1    g519(.A(G900), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n476), .B1(new_n478), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n678), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n343), .A2(new_n705), .A3(new_n597), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G128), .ZN(G30));
  INV_X1    g524(.A(new_n697), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n474), .A2(new_n345), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n711), .A2(new_n550), .A3(new_n552), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(KEYINPUT106), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n323), .A2(new_n244), .ZN(new_n715));
  AOI22_X1  g529(.A1(new_n285), .A2(new_n292), .B1(new_n282), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g530(.A(G472), .B1(new_n716), .B2(G902), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n321), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n427), .B(KEYINPUT38), .ZN(new_n719));
  XOR2_X1   g533(.A(KEYINPUT107), .B(KEYINPUT39), .Z(new_n720));
  XNOR2_X1  g534(.A(new_n707), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n597), .A2(new_n721), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n718), .B(new_n719), .C1(new_n722), .C2(KEYINPUT40), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n723), .B1(KEYINPUT40), .B2(new_n722), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n714), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G143), .ZN(G45));
  NOR2_X1   g540(.A1(new_n667), .A2(new_n707), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n343), .A2(new_n705), .A3(new_n597), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G146), .ZN(G48));
  NAND2_X1  g543(.A1(new_n653), .A2(new_n655), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n306), .A2(KEYINPUT32), .A3(new_n308), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n319), .B1(new_n318), .B2(new_n307), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n340), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(KEYINPUT74), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n321), .A2(new_n322), .A3(new_n340), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n467), .B1(new_n584), .B2(new_n585), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(G469), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n737), .A2(new_n595), .A3(new_n586), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n734), .A2(new_n735), .A3(new_n669), .A4(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n730), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g554(.A(KEYINPUT41), .B(G113), .Z(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G15));
  AND4_X1   g556(.A1(new_n734), .A2(new_n684), .A3(new_n735), .A4(new_n738), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n658), .A2(new_n743), .A3(KEYINPUT108), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT108), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n734), .A2(new_n684), .A3(new_n735), .A4(new_n738), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n745), .B1(new_n730), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G116), .ZN(G18));
  NAND4_X1  g563(.A1(new_n734), .A2(new_n735), .A3(new_n553), .A4(new_n697), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n680), .A2(new_n737), .A3(new_n595), .A4(new_n586), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT109), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(new_n365), .ZN(G21));
  AND2_X1   g569(.A1(new_n738), .A2(new_n482), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n550), .A2(new_n427), .A3(new_n552), .A4(new_n712), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n757), .A2(KEYINPUT112), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n757), .A2(KEYINPUT112), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n756), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n652), .ZN(new_n761));
  OR3_X1    g575(.A1(new_n314), .A2(KEYINPUT110), .A3(new_n324), .ZN(new_n762));
  OAI21_X1  g576(.A(KEYINPUT110), .B1(new_n314), .B2(new_n324), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(new_n282), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n280), .A2(new_n293), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n308), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n670), .A2(KEYINPUT111), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n768), .B(G472), .C1(new_n306), .C2(G902), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n766), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n761), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n760), .A2(new_n771), .ZN(new_n772));
  XOR2_X1   g586(.A(new_n772), .B(G122), .Z(G24));
  AND2_X1   g587(.A1(new_n770), .A2(new_n697), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n751), .B(KEYINPUT109), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(new_n775), .A3(new_n727), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G125), .ZN(G27));
  INV_X1    g591(.A(KEYINPUT42), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n653), .A2(new_n734), .A3(new_n735), .A4(new_n655), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n591), .A2(KEYINPUT113), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n591), .A2(KEYINPUT113), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n780), .A2(new_n586), .A3(new_n593), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n346), .A2(new_n595), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n427), .A2(new_n783), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n727), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n778), .B1(new_n779), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n652), .B1(new_n340), .B2(new_n321), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n788), .A2(KEYINPUT42), .A3(new_n727), .A4(new_n785), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G131), .ZN(G33));
  NAND2_X1  g605(.A1(new_n785), .A2(new_n708), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n779), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(new_n205), .ZN(G36));
  NAND2_X1  g608(.A1(new_n589), .A2(new_n590), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT45), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT114), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n554), .B1(new_n795), .B2(new_n796), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n592), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(KEYINPUT46), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n586), .B1(new_n800), .B2(KEYINPUT46), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n595), .B(new_n721), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n425), .A2(new_n346), .A3(new_n426), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n688), .A2(new_n666), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT43), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n809), .A2(new_n671), .A3(new_n697), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT44), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n806), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G137), .ZN(G39));
  NOR4_X1   g629(.A1(new_n343), .A2(new_n667), .A3(new_n707), .A4(new_n805), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n800), .A2(KEYINPUT46), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n817), .A2(new_n586), .A3(new_n801), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT47), .B1(new_n818), .B2(new_n595), .ZN(new_n819));
  OAI211_X1 g633(.A(KEYINPUT47), .B(new_n595), .C1(new_n802), .C2(new_n803), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n730), .B(new_n816), .C1(new_n819), .C2(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(G140), .ZN(G42));
  NAND2_X1  g637(.A1(new_n737), .A2(new_n586), .ZN(new_n824));
  XOR2_X1   g638(.A(new_n824), .B(KEYINPUT49), .Z(new_n825));
  NOR2_X1   g639(.A1(new_n718), .A2(new_n783), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n807), .A2(new_n719), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n825), .A2(new_n761), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n757), .B(KEYINPUT112), .ZN(new_n830));
  INV_X1    g644(.A(new_n707), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n831), .A2(new_n595), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n718), .A2(new_n782), .A3(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n830), .A2(new_n711), .A3(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n709), .A2(new_n728), .A3(new_n776), .A4(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n835), .A2(new_n836), .A3(KEYINPUT52), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT52), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT116), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n836), .A2(KEYINPUT52), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n837), .B1(new_n835), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n422), .A2(new_n429), .A3(new_n482), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT115), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n474), .B(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n688), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n843), .B1(new_n846), .B2(new_n667), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n847), .A2(new_n653), .A3(new_n655), .A4(new_n672), .ZN(new_n848));
  INV_X1    g662(.A(new_n598), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n848), .B1(new_n779), .B2(new_n849), .ZN(new_n850));
  OAI22_X1  g664(.A1(new_n760), .A2(new_n771), .B1(new_n750), .B2(new_n753), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n698), .B1(new_n730), .B2(new_n739), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NOR4_X1   g667(.A1(new_n845), .A2(new_n805), .A3(new_n549), .A4(new_n707), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n734), .A2(new_n854), .A3(new_n735), .A4(new_n597), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n785), .A2(new_n770), .A3(new_n727), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n711), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n793), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n853), .A2(new_n748), .A3(new_n790), .A4(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n829), .B1(new_n842), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n851), .A2(new_n852), .ZN(new_n861));
  INV_X1    g675(.A(new_n850), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(new_n748), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n790), .A2(new_n858), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n835), .B(new_n838), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n865), .A2(new_n866), .A3(KEYINPUT53), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n860), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT54), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n809), .A2(new_n476), .ZN(new_n870));
  INV_X1    g684(.A(new_n771), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n738), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n873), .A2(new_n719), .A3(new_n346), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT50), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n872), .A2(KEYINPUT50), .A3(new_n874), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT117), .ZN(new_n880));
  INV_X1    g694(.A(new_n805), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n819), .A2(new_n821), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n824), .A2(new_n595), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n881), .B(new_n872), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n873), .A2(new_n805), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n870), .A2(new_n774), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT118), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n870), .A2(KEYINPUT118), .A3(new_n774), .A4(new_n885), .ZN(new_n889));
  INV_X1    g703(.A(new_n885), .ZN(new_n890));
  NOR4_X1   g704(.A1(new_n730), .A2(new_n890), .A3(new_n477), .A4(new_n718), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n666), .B1(new_n550), .B2(new_n552), .ZN(new_n892));
  AOI22_X1  g706(.A1(new_n888), .A2(new_n889), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT117), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n877), .A2(new_n894), .A3(new_n878), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n880), .A2(new_n884), .A3(new_n893), .A4(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT51), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n835), .B(KEYINPUT52), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n829), .B1(new_n899), .B2(new_n859), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n709), .A2(new_n776), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n734), .A2(new_n735), .A3(new_n597), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n697), .A2(new_n680), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n718), .A2(new_n782), .A3(new_n832), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n905), .A2(new_n697), .ZN(new_n906));
  AOI22_X1  g720(.A1(new_n904), .A2(new_n727), .B1(new_n830), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n840), .B1(new_n901), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n835), .A2(new_n841), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n865), .A2(new_n910), .A3(KEYINPUT53), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT54), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n900), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI211_X1 g727(.A(new_n475), .B(G953), .C1(new_n872), .C2(new_n775), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n870), .A2(new_n788), .A3(new_n885), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT48), .ZN(new_n916));
  INV_X1    g730(.A(new_n667), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n891), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n914), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n884), .A2(new_n893), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n897), .B1(new_n877), .B2(new_n878), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AND4_X1   g736(.A1(new_n869), .A2(new_n898), .A3(new_n913), .A4(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(G952), .A2(G953), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n828), .B1(new_n923), .B2(new_n924), .ZN(G75));
  NOR2_X1   g739(.A1(new_n248), .A2(G952), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT119), .Z(new_n927));
  NAND2_X1  g741(.A1(new_n412), .A2(new_n414), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(new_n416), .Z(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT55), .ZN(new_n930));
  NAND2_X1  g744(.A1(G210), .A2(G902), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n842), .A2(new_n859), .A3(new_n829), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT53), .B1(new_n865), .B2(new_n866), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT56), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n930), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n931), .B1(new_n900), .B2(new_n911), .ZN(new_n938));
  INV_X1    g752(.A(new_n930), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n938), .A2(KEYINPUT56), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n927), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(KEYINPUT120), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT120), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n943), .B(new_n927), .C1(new_n937), .C2(new_n940), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n942), .A2(new_n944), .ZN(G51));
  NAND2_X1  g759(.A1(new_n900), .A2(new_n911), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(KEYINPUT54), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n913), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n592), .B(KEYINPUT57), .Z(new_n950));
  OAI22_X1  g764(.A1(new_n949), .A2(new_n950), .B1(new_n585), .B2(new_n584), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n467), .B1(new_n900), .B2(new_n911), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n952), .A2(new_n798), .A3(new_n799), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n926), .B1(new_n951), .B2(new_n953), .ZN(G54));
  NAND3_X1  g768(.A1(new_n952), .A2(KEYINPUT58), .A3(G475), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n543), .A2(new_n526), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n955), .A2(new_n956), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n957), .A2(new_n958), .A3(new_n926), .ZN(G60));
  INV_X1    g773(.A(KEYINPUT122), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n659), .B(KEYINPUT59), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n961), .B1(new_n869), .B2(new_n913), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n663), .A2(new_n664), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT121), .Z(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n960), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n961), .ZN(new_n967));
  INV_X1    g781(.A(new_n913), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n912), .B1(new_n860), .B2(new_n867), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n970), .A2(KEYINPUT122), .A3(new_n964), .ZN(new_n971));
  INV_X1    g785(.A(new_n927), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n964), .A2(new_n961), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n972), .B1(new_n948), .B2(new_n973), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n966), .A2(new_n971), .A3(new_n974), .ZN(G63));
  NAND2_X1  g789(.A1(G217), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT60), .Z(new_n977));
  NAND2_X1  g791(.A1(new_n946), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n631), .A2(new_n635), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n972), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n693), .A2(new_n695), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n980), .B1(new_n981), .B2(new_n978), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT61), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n980), .B(KEYINPUT61), .C1(new_n981), .C2(new_n978), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(G66));
  INV_X1    g800(.A(new_n481), .ZN(new_n987));
  OAI21_X1  g801(.A(G953), .B1(new_n987), .B2(new_n393), .ZN(new_n988));
  INV_X1    g802(.A(new_n863), .ZN(new_n989));
  INV_X1    g803(.A(new_n248), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n928), .B1(G898), .B2(new_n248), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n991), .B(new_n992), .ZN(G69));
  INV_X1    g807(.A(KEYINPUT125), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n788), .A2(new_n830), .ZN(new_n995));
  OR3_X1    g809(.A1(new_n804), .A2(KEYINPUT124), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(KEYINPUT124), .B1(new_n804), .B2(new_n995), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n793), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AND2_X1   g812(.A1(new_n901), .A2(new_n728), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n822), .A2(new_n814), .A3(new_n790), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n994), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  AND3_X1   g816(.A1(new_n822), .A2(new_n814), .A3(new_n790), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n1003), .A2(KEYINPUT125), .A3(new_n999), .A4(new_n998), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n1002), .A2(new_n1004), .A3(new_n248), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n286), .A2(new_n262), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1006), .B(KEYINPUT123), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n533), .A2(new_n534), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1009), .B1(G900), .B2(new_n990), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1005), .A2(new_n1010), .ZN(new_n1011));
  AND2_X1   g825(.A1(new_n846), .A2(new_n667), .ZN(new_n1012));
  OR4_X1    g826(.A1(new_n779), .A2(new_n722), .A3(new_n805), .A4(new_n1012), .ZN(new_n1013));
  AND3_X1   g827(.A1(new_n822), .A2(new_n814), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT62), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n999), .A2(new_n1015), .A3(new_n725), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n999), .A2(new_n725), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(KEYINPUT62), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1014), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(new_n248), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n248), .B1(G227), .B2(G900), .ZN(new_n1021));
  AOI22_X1  g835(.A1(new_n1020), .A2(new_n1009), .B1(KEYINPUT126), .B2(new_n1021), .ZN(new_n1022));
  OR2_X1    g836(.A1(new_n1021), .A2(KEYINPUT126), .ZN(new_n1023));
  AND3_X1   g837(.A1(new_n1011), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1023), .B1(new_n1011), .B2(new_n1022), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n1024), .A2(new_n1025), .ZN(G72));
  NAND3_X1  g840(.A1(new_n1002), .A2(new_n1004), .A3(new_n989), .ZN(new_n1027));
  NAND2_X1  g841(.A1(G472), .A2(G902), .ZN(new_n1028));
  XOR2_X1   g842(.A(new_n1028), .B(KEYINPUT63), .Z(new_n1029));
  AOI211_X1 g843(.A(new_n334), .B(new_n258), .C1(new_n1027), .C2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g844(.A1(new_n1014), .A2(new_n1018), .A3(new_n989), .A4(new_n1016), .ZN(new_n1031));
  AOI211_X1 g845(.A(new_n330), .B(new_n282), .C1(new_n1031), .C2(new_n1029), .ZN(new_n1032));
  NOR2_X1   g846(.A1(new_n261), .A2(new_n279), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1029), .B1(new_n336), .B2(new_n1033), .ZN(new_n1034));
  XOR2_X1   g848(.A(new_n1034), .B(KEYINPUT127), .Z(new_n1035));
  AOI21_X1  g849(.A(new_n1035), .B1(new_n860), .B2(new_n867), .ZN(new_n1036));
  NOR4_X1   g850(.A1(new_n1030), .A2(new_n1032), .A3(new_n926), .A4(new_n1036), .ZN(G57));
endmodule


