

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741;

  NOR2_X1 U369 ( .A1(n684), .A2(n683), .ZN(n598) );
  XNOR2_X1 U370 ( .A(KEYINPUT64), .B(KEYINPUT82), .ZN(n405) );
  NAND2_X1 U371 ( .A1(n355), .A2(n352), .ZN(n517) );
  INV_X1 U372 ( .A(G953), .ZN(n734) );
  NOR2_X2 U373 ( .A1(n614), .A2(n711), .ZN(n616) );
  NOR2_X1 U374 ( .A1(n588), .A2(n385), .ZN(n563) );
  XNOR2_X2 U375 ( .A(n522), .B(n380), .ZN(n741) );
  NOR2_X4 U376 ( .A1(n378), .A2(n691), .ZN(n706) );
  NOR2_X1 U377 ( .A1(n566), .A2(n565), .ZN(n568) );
  AND2_X2 U378 ( .A1(n602), .A2(n601), .ZN(n378) );
  NOR2_X1 U379 ( .A1(n364), .A2(n361), .ZN(n555) );
  XNOR2_X1 U380 ( .A(n504), .B(n503), .ZN(n573) );
  XNOR2_X1 U381 ( .A(n464), .B(n463), .ZN(n590) );
  BUF_X1 U382 ( .A(n505), .Z(n535) );
  XNOR2_X1 U383 ( .A(n422), .B(n421), .ZN(n505) );
  XNOR2_X1 U384 ( .A(n474), .B(n473), .ZN(n506) );
  OR2_X1 U385 ( .A1(n698), .A2(n600), .ZN(n422) );
  XNOR2_X1 U386 ( .A(n431), .B(n368), .ZN(n725) );
  INV_X1 U387 ( .A(n404), .ZN(n406) );
  XNOR2_X1 U388 ( .A(G128), .B(G143), .ZN(n404) );
  XNOR2_X2 U389 ( .A(n373), .B(KEYINPUT19), .ZN(n429) );
  XNOR2_X1 U390 ( .A(G146), .B(G125), .ZN(n431) );
  NAND2_X1 U391 ( .A1(n741), .A2(KEYINPUT46), .ZN(n362) );
  XNOR2_X1 U392 ( .A(KEYINPUT85), .B(KEYINPUT24), .ZN(n478) );
  XNOR2_X1 U393 ( .A(KEYINPUT67), .B(G101), .ZN(n408) );
  NOR2_X1 U394 ( .A1(n506), .A2(n384), .ZN(n383) );
  INV_X1 U395 ( .A(n665), .ZN(n384) );
  OR2_X1 U396 ( .A1(n611), .A2(G902), .ZN(n370) );
  XOR2_X1 U397 ( .A(KEYINPUT3), .B(G119), .Z(n410) );
  NOR2_X1 U398 ( .A1(n741), .A2(KEYINPUT46), .ZN(n366) );
  NAND2_X1 U399 ( .A1(n363), .A2(n362), .ZN(n361) );
  AND2_X1 U400 ( .A1(n357), .A2(n356), .ZN(n355) );
  NAND2_X1 U401 ( .A1(n499), .A2(n354), .ZN(n353) );
  XNOR2_X1 U402 ( .A(n472), .B(n471), .ZN(n473) );
  NOR2_X1 U403 ( .A1(n617), .A2(G902), .ZN(n474) );
  XNOR2_X1 U404 ( .A(G137), .B(G134), .ZN(n465) );
  XNOR2_X1 U405 ( .A(n390), .B(n483), .ZN(n611) );
  XNOR2_X1 U406 ( .A(n482), .B(n401), .ZN(n483) );
  XNOR2_X1 U407 ( .A(n484), .B(n485), .ZN(n390) );
  XNOR2_X1 U408 ( .A(n358), .B(n379), .ZN(n698) );
  XNOR2_X1 U409 ( .A(n717), .B(n419), .ZN(n379) );
  NOR2_X1 U410 ( .A1(n524), .A2(n523), .ZN(n526) );
  NOR2_X1 U411 ( .A1(n378), .A2(n397), .ZN(n393) );
  INV_X1 U412 ( .A(G217), .ZN(n397) );
  NAND2_X1 U413 ( .A1(n394), .A2(n395), .ZN(n389) );
  NOR2_X1 U414 ( .A1(n378), .A2(n396), .ZN(n395) );
  INV_X1 U415 ( .A(G210), .ZN(n396) );
  NAND2_X1 U416 ( .A1(n553), .A2(n365), .ZN(n364) );
  NAND2_X1 U417 ( .A1(n367), .A2(n366), .ZN(n365) );
  NAND2_X1 U418 ( .A1(G469), .A2(G902), .ZN(n356) );
  INV_X1 U419 ( .A(G472), .ZN(n471) );
  INV_X1 U420 ( .A(KEYINPUT4), .ZN(n407) );
  XOR2_X1 U421 ( .A(KEYINPUT23), .B(KEYINPUT96), .Z(n481) );
  XNOR2_X1 U422 ( .A(G128), .B(G119), .ZN(n476) );
  XOR2_X1 U423 ( .A(G110), .B(G137), .Z(n477) );
  XNOR2_X1 U424 ( .A(n369), .B(G140), .ZN(n368) );
  INV_X1 U425 ( .A(KEYINPUT10), .ZN(n369) );
  XOR2_X1 U426 ( .A(G146), .B(G140), .Z(n491) );
  XNOR2_X1 U427 ( .A(n376), .B(n412), .ZN(n493) );
  XNOR2_X1 U428 ( .A(n377), .B(G110), .ZN(n376) );
  XNOR2_X1 U429 ( .A(G107), .B(KEYINPUT92), .ZN(n377) );
  INV_X1 U430 ( .A(KEYINPUT94), .ZN(n494) );
  XNOR2_X1 U431 ( .A(n535), .B(n519), .ZN(n666) );
  INV_X1 U432 ( .A(KEYINPUT38), .ZN(n519) );
  XNOR2_X1 U433 ( .A(n517), .B(KEYINPUT1), .ZN(n375) );
  OR2_X1 U434 ( .A1(n684), .A2(n683), .ZN(n732) );
  XNOR2_X1 U435 ( .A(G116), .B(G107), .ZN(n448) );
  XNOR2_X1 U436 ( .A(n392), .B(n391), .ZN(n479) );
  INV_X1 U437 ( .A(KEYINPUT8), .ZN(n391) );
  NAND2_X1 U438 ( .A1(n734), .A2(G234), .ZN(n392) );
  AND2_X1 U439 ( .A1(n687), .A2(KEYINPUT2), .ZN(n596) );
  BUF_X1 U440 ( .A(n375), .Z(n374) );
  XNOR2_X1 U441 ( .A(n359), .B(KEYINPUT78), .ZN(n524) );
  NAND2_X1 U442 ( .A1(n561), .A2(n402), .ZN(n577) );
  INV_X1 U443 ( .A(KEYINPUT0), .ZN(n372) );
  XNOR2_X1 U444 ( .A(n506), .B(n475), .ZN(n588) );
  XNOR2_X1 U445 ( .A(n358), .B(n470), .ZN(n617) );
  XNOR2_X1 U446 ( .A(KEYINPUT42), .B(KEYINPUT109), .ZN(n380) );
  OR2_X1 U447 ( .A1(n540), .A2(n680), .ZN(n522) );
  XNOR2_X1 U448 ( .A(n381), .B(n528), .ZN(n740) );
  NOR2_X1 U449 ( .A1(n540), .A2(n398), .ZN(n635) );
  INV_X1 U450 ( .A(KEYINPUT56), .ZN(n386) );
  XOR2_X1 U451 ( .A(KEYINPUT69), .B(G131), .Z(n347) );
  AND2_X1 U452 ( .A1(n520), .A2(n402), .ZN(n348) );
  XOR2_X1 U453 ( .A(n488), .B(n487), .Z(n349) );
  INV_X1 U454 ( .A(n561), .ZN(n569) );
  XNOR2_X1 U455 ( .A(n370), .B(n349), .ZN(n561) );
  INV_X1 U456 ( .A(G902), .ZN(n354) );
  XNOR2_X1 U457 ( .A(n699), .B(n698), .ZN(n350) );
  XNOR2_X1 U458 ( .A(n564), .B(KEYINPUT34), .ZN(n566) );
  NAND2_X1 U459 ( .A1(n371), .A2(n580), .ZN(n564) );
  XNOR2_X2 U460 ( .A(n595), .B(n594), .ZN(n687) );
  XNOR2_X2 U461 ( .A(n351), .B(KEYINPUT77), .ZN(n691) );
  NAND2_X1 U462 ( .A1(n596), .A2(n598), .ZN(n351) );
  OR2_X1 U463 ( .A1(n700), .A2(n353), .ZN(n352) );
  NAND2_X1 U464 ( .A1(n700), .A2(G469), .ZN(n357) );
  NAND2_X1 U465 ( .A1(n653), .A2(n375), .ZN(n385) );
  XNOR2_X2 U466 ( .A(n497), .B(n716), .ZN(n358) );
  XNOR2_X2 U467 ( .A(n726), .B(n408), .ZN(n497) );
  XNOR2_X2 U468 ( .A(n447), .B(n407), .ZN(n726) );
  NAND2_X1 U469 ( .A1(n382), .A2(n360), .ZN(n359) );
  AND2_X1 U470 ( .A1(n512), .A2(n561), .ZN(n360) );
  NAND2_X1 U471 ( .A1(n740), .A2(KEYINPUT46), .ZN(n363) );
  INV_X1 U472 ( .A(n740), .ZN(n367) );
  INV_X1 U473 ( .A(n663), .ZN(n371) );
  NAND2_X1 U474 ( .A1(n580), .A2(n348), .ZN(n464) );
  NAND2_X1 U475 ( .A1(n580), .A2(n659), .ZN(n583) );
  XNOR2_X2 U476 ( .A(n430), .B(n372), .ZN(n580) );
  NAND2_X1 U477 ( .A1(n429), .A2(n403), .ZN(n430) );
  NAND2_X1 U478 ( .A1(n505), .A2(n665), .ZN(n373) );
  INV_X1 U479 ( .A(n374), .ZN(n586) );
  NOR2_X1 U480 ( .A1(n653), .A2(n374), .ZN(n654) );
  NOR2_X1 U481 ( .A1(n557), .A2(n374), .ZN(n558) );
  NAND2_X1 U482 ( .A1(n538), .A2(n374), .ZN(n645) );
  XNOR2_X1 U483 ( .A(n493), .B(n492), .ZN(n496) );
  XNOR2_X1 U484 ( .A(n493), .B(n414), .ZN(n717) );
  NAND2_X1 U485 ( .A1(n556), .A2(n638), .ZN(n381) );
  INV_X1 U486 ( .A(n506), .ZN(n578) );
  XNOR2_X1 U487 ( .A(n383), .B(KEYINPUT30), .ZN(n382) );
  NOR2_X1 U488 ( .A1(n385), .A2(n652), .ZN(n659) );
  XNOR2_X1 U489 ( .A(n387), .B(n386), .ZN(G51) );
  NAND2_X1 U490 ( .A1(n388), .A2(n620), .ZN(n387) );
  XNOR2_X1 U491 ( .A(n389), .B(n350), .ZN(n388) );
  NAND2_X1 U492 ( .A1(n394), .A2(n393), .ZN(n613) );
  INV_X1 U493 ( .A(n691), .ZN(n394) );
  NAND2_X1 U494 ( .A1(n706), .A2(G472), .ZN(n619) );
  NAND2_X1 U495 ( .A1(n706), .A2(G475), .ZN(n606) );
  INV_X1 U496 ( .A(n429), .ZN(n398) );
  AND2_X1 U497 ( .A1(n547), .A2(n546), .ZN(n399) );
  AND2_X1 U498 ( .A1(n592), .A2(n591), .ZN(n400) );
  XOR2_X1 U499 ( .A(n481), .B(n480), .Z(n401) );
  XOR2_X1 U500 ( .A(n462), .B(n461), .Z(n402) );
  NAND2_X1 U501 ( .A1(n509), .A2(n428), .ZN(n403) );
  INV_X1 U502 ( .A(KEYINPUT44), .ZN(n575) );
  XNOR2_X1 U503 ( .A(n725), .B(n478), .ZN(n484) );
  NAND2_X1 U504 ( .A1(n666), .A2(n665), .ZN(n670) );
  XNOR2_X1 U505 ( .A(n496), .B(n728), .ZN(n498) );
  XNOR2_X1 U506 ( .A(n495), .B(n494), .ZN(n728) );
  INV_X1 U507 ( .A(KEYINPUT35), .ZN(n567) );
  INV_X1 U508 ( .A(KEYINPUT40), .ZN(n528) );
  AND2_X1 U509 ( .A1(n607), .A2(G953), .ZN(n711) );
  XNOR2_X2 U510 ( .A(n406), .B(n405), .ZN(n447) );
  XNOR2_X1 U511 ( .A(G116), .B(G113), .ZN(n409) );
  XNOR2_X1 U512 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U513 ( .A(n411), .B(KEYINPUT71), .ZN(n716) );
  XNOR2_X1 U514 ( .A(G104), .B(KEYINPUT76), .ZN(n412) );
  XNOR2_X1 U515 ( .A(KEYINPUT16), .B(G122), .ZN(n413) );
  XNOR2_X1 U516 ( .A(n413), .B(KEYINPUT75), .ZN(n414) );
  XNOR2_X1 U517 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n415) );
  XNOR2_X1 U518 ( .A(n431), .B(n415), .ZN(n418) );
  NAND2_X1 U519 ( .A1(n734), .A2(G224), .ZN(n416) );
  XNOR2_X1 U520 ( .A(n416), .B(KEYINPUT80), .ZN(n417) );
  XNOR2_X1 U521 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U522 ( .A(KEYINPUT15), .B(G902), .ZN(n459) );
  INV_X1 U523 ( .A(n459), .ZN(n600) );
  INV_X1 U524 ( .A(G237), .ZN(n420) );
  NAND2_X1 U525 ( .A1(n354), .A2(n420), .ZN(n423) );
  AND2_X1 U526 ( .A1(n423), .A2(G210), .ZN(n421) );
  NAND2_X1 U527 ( .A1(n423), .A2(G214), .ZN(n665) );
  NAND2_X1 U528 ( .A1(G234), .A2(G237), .ZN(n424) );
  XNOR2_X1 U529 ( .A(n424), .B(KEYINPUT14), .ZN(n426) );
  NAND2_X1 U530 ( .A1(G952), .A2(n426), .ZN(n425) );
  XNOR2_X1 U531 ( .A(KEYINPUT93), .B(n425), .ZN(n679) );
  NAND2_X1 U532 ( .A1(n679), .A2(n734), .ZN(n509) );
  NAND2_X1 U533 ( .A1(G902), .A2(n426), .ZN(n507) );
  INV_X1 U534 ( .A(n507), .ZN(n427) );
  NOR2_X1 U535 ( .A1(G898), .A2(n734), .ZN(n721) );
  NAND2_X1 U536 ( .A1(n427), .A2(n721), .ZN(n428) );
  XOR2_X1 U537 ( .A(G131), .B(KEYINPUT98), .Z(n433) );
  NOR2_X1 U538 ( .A1(G953), .A2(G237), .ZN(n466) );
  NAND2_X1 U539 ( .A1(G214), .A2(n466), .ZN(n432) );
  XNOR2_X1 U540 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U541 ( .A(n725), .B(n434), .ZN(n442) );
  XOR2_X1 U542 ( .A(G122), .B(G104), .Z(n436) );
  XNOR2_X1 U543 ( .A(G143), .B(G113), .ZN(n435) );
  XNOR2_X1 U544 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U545 ( .A(KEYINPUT100), .B(KEYINPUT12), .Z(n438) );
  XNOR2_X1 U546 ( .A(KEYINPUT11), .B(KEYINPUT99), .ZN(n437) );
  XNOR2_X1 U547 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U548 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U549 ( .A(n442), .B(n441), .ZN(n604) );
  NOR2_X1 U550 ( .A1(G902), .A2(n604), .ZN(n444) );
  XNOR2_X1 U551 ( .A(KEYINPUT13), .B(KEYINPUT101), .ZN(n443) );
  XNOR2_X1 U552 ( .A(n444), .B(n443), .ZN(n446) );
  INV_X1 U553 ( .A(G475), .ZN(n445) );
  XNOR2_X1 U554 ( .A(n446), .B(n445), .ZN(n527) );
  XOR2_X1 U555 ( .A(KEYINPUT103), .B(G122), .Z(n449) );
  XNOR2_X1 U556 ( .A(n449), .B(n448), .ZN(n453) );
  XOR2_X1 U557 ( .A(KEYINPUT9), .B(KEYINPUT104), .Z(n451) );
  XNOR2_X1 U558 ( .A(G134), .B(KEYINPUT7), .ZN(n450) );
  XNOR2_X1 U559 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U560 ( .A(n453), .B(n452), .Z(n455) );
  NAND2_X1 U561 ( .A1(G217), .A2(n479), .ZN(n454) );
  XNOR2_X1 U562 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U563 ( .A(n447), .B(n456), .Z(n707) );
  NOR2_X1 U564 ( .A1(G902), .A2(n707), .ZN(n458) );
  XNOR2_X1 U565 ( .A(KEYINPUT105), .B(G478), .ZN(n457) );
  XNOR2_X1 U566 ( .A(n458), .B(n457), .ZN(n543) );
  NOR2_X1 U567 ( .A1(n527), .A2(n543), .ZN(n520) );
  NAND2_X1 U568 ( .A1(n459), .A2(G234), .ZN(n460) );
  XNOR2_X1 U569 ( .A(n460), .B(KEYINPUT20), .ZN(n486) );
  AND2_X1 U570 ( .A1(n486), .A2(G221), .ZN(n462) );
  XNOR2_X1 U571 ( .A(KEYINPUT97), .B(KEYINPUT21), .ZN(n461) );
  XNOR2_X1 U572 ( .A(KEYINPUT65), .B(KEYINPUT22), .ZN(n463) );
  XNOR2_X1 U573 ( .A(n347), .B(n465), .ZN(n495) );
  XOR2_X1 U574 ( .A(G146), .B(KEYINPUT5), .Z(n468) );
  NAND2_X1 U575 ( .A1(n466), .A2(G210), .ZN(n467) );
  XNOR2_X1 U576 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U577 ( .A(n495), .B(n469), .ZN(n470) );
  INV_X1 U578 ( .A(KEYINPUT74), .ZN(n472) );
  INV_X1 U579 ( .A(KEYINPUT6), .ZN(n475) );
  INV_X1 U580 ( .A(n588), .ZN(n531) );
  XNOR2_X1 U581 ( .A(n477), .B(n476), .ZN(n485) );
  NAND2_X1 U582 ( .A1(G221), .A2(n479), .ZN(n482) );
  XNOR2_X1 U583 ( .A(KEYINPUT72), .B(KEYINPUT95), .ZN(n480) );
  XOR2_X1 U584 ( .A(KEYINPUT79), .B(KEYINPUT25), .Z(n488) );
  NAND2_X1 U585 ( .A1(n486), .A2(G217), .ZN(n487) );
  INV_X1 U586 ( .A(KEYINPUT106), .ZN(n489) );
  XNOR2_X1 U587 ( .A(n569), .B(n489), .ZN(n649) );
  NAND2_X1 U588 ( .A1(G227), .A2(n734), .ZN(n490) );
  XNOR2_X1 U589 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U590 ( .A(n497), .B(n498), .ZN(n700) );
  INV_X1 U591 ( .A(G469), .ZN(n499) );
  NOR2_X1 U592 ( .A1(n649), .A2(n586), .ZN(n500) );
  XNOR2_X1 U593 ( .A(n500), .B(KEYINPUT107), .ZN(n501) );
  NOR2_X1 U594 ( .A1(n531), .A2(n501), .ZN(n502) );
  NAND2_X1 U595 ( .A1(n590), .A2(n502), .ZN(n504) );
  XOR2_X1 U596 ( .A(KEYINPUT81), .B(KEYINPUT32), .Z(n503) );
  XNOR2_X1 U597 ( .A(n573), .B(G119), .ZN(G21) );
  INV_X1 U598 ( .A(n517), .ZN(n582) );
  NOR2_X1 U599 ( .A1(G900), .A2(n507), .ZN(n508) );
  NAND2_X1 U600 ( .A1(n508), .A2(G953), .ZN(n510) );
  NAND2_X1 U601 ( .A1(n510), .A2(n509), .ZN(n511) );
  NAND2_X1 U602 ( .A1(n511), .A2(n402), .ZN(n514) );
  NOR2_X1 U603 ( .A1(n582), .A2(n514), .ZN(n512) );
  NAND2_X1 U604 ( .A1(n527), .A2(n543), .ZN(n565) );
  NOR2_X1 U605 ( .A1(n524), .A2(n565), .ZN(n513) );
  NAND2_X1 U606 ( .A1(n535), .A2(n513), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n539), .B(G143), .ZN(G45) );
  XNOR2_X1 U608 ( .A(KEYINPUT70), .B(n514), .ZN(n529) );
  NAND2_X1 U609 ( .A1(n569), .A2(n578), .ZN(n515) );
  NOR2_X1 U610 ( .A1(n529), .A2(n515), .ZN(n516) );
  XNOR2_X1 U611 ( .A(KEYINPUT28), .B(n516), .ZN(n518) );
  NAND2_X1 U612 ( .A1(n518), .A2(n517), .ZN(n540) );
  INV_X1 U613 ( .A(n520), .ZN(n669) );
  NOR2_X1 U614 ( .A1(n670), .A2(n669), .ZN(n521) );
  XNOR2_X1 U615 ( .A(KEYINPUT41), .B(n521), .ZN(n680) );
  INV_X1 U616 ( .A(n666), .ZN(n523) );
  XNOR2_X1 U617 ( .A(KEYINPUT73), .B(KEYINPUT39), .ZN(n525) );
  XNOR2_X1 U618 ( .A(n526), .B(n525), .ZN(n556) );
  XOR2_X1 U619 ( .A(KEYINPUT102), .B(n527), .Z(n544) );
  NOR2_X1 U620 ( .A1(n544), .A2(n543), .ZN(n638) );
  INV_X1 U621 ( .A(n529), .ZN(n530) );
  NAND2_X1 U622 ( .A1(n665), .A2(n530), .ZN(n533) );
  NAND2_X1 U623 ( .A1(n638), .A2(n531), .ZN(n532) );
  NOR2_X1 U624 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U625 ( .A1(n534), .A2(n569), .ZN(n557) );
  INV_X1 U626 ( .A(n535), .ZN(n559) );
  NOR2_X1 U627 ( .A1(n557), .A2(n559), .ZN(n537) );
  XNOR2_X1 U628 ( .A(KEYINPUT110), .B(KEYINPUT36), .ZN(n536) );
  XNOR2_X1 U629 ( .A(n537), .B(n536), .ZN(n538) );
  NAND2_X1 U630 ( .A1(n645), .A2(n539), .ZN(n552) );
  XOR2_X1 U631 ( .A(KEYINPUT47), .B(KEYINPUT68), .Z(n541) );
  NAND2_X1 U632 ( .A1(n635), .A2(n541), .ZN(n542) );
  NAND2_X1 U633 ( .A1(n542), .A2(KEYINPUT84), .ZN(n545) );
  AND2_X1 U634 ( .A1(n544), .A2(n543), .ZN(n641) );
  NOR2_X1 U635 ( .A1(n638), .A2(n641), .ZN(n671) );
  INV_X1 U636 ( .A(n671), .ZN(n584) );
  NAND2_X1 U637 ( .A1(n545), .A2(n584), .ZN(n547) );
  OR2_X1 U638 ( .A1(KEYINPUT84), .A2(KEYINPUT47), .ZN(n546) );
  NAND2_X1 U639 ( .A1(n671), .A2(KEYINPUT84), .ZN(n548) );
  NAND2_X1 U640 ( .A1(n635), .A2(n548), .ZN(n549) );
  NAND2_X1 U641 ( .A1(n549), .A2(KEYINPUT47), .ZN(n550) );
  NAND2_X1 U642 ( .A1(n399), .A2(n550), .ZN(n551) );
  NOR2_X1 U643 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U644 ( .A(KEYINPUT48), .B(KEYINPUT89), .ZN(n554) );
  XNOR2_X1 U645 ( .A(n555), .B(n554), .ZN(n684) );
  NAND2_X1 U646 ( .A1(n556), .A2(n641), .ZN(n646) );
  XOR2_X1 U647 ( .A(n558), .B(KEYINPUT43), .Z(n560) );
  NAND2_X1 U648 ( .A1(n560), .A2(n559), .ZN(n647) );
  NAND2_X1 U649 ( .A1(n646), .A2(n647), .ZN(n683) );
  INV_X1 U650 ( .A(n577), .ZN(n653) );
  XNOR2_X1 U651 ( .A(KEYINPUT108), .B(KEYINPUT33), .ZN(n562) );
  XNOR2_X1 U652 ( .A(n563), .B(n562), .ZN(n663) );
  XNOR2_X1 U653 ( .A(n568), .B(n567), .ZN(n738) );
  INV_X1 U654 ( .A(n578), .ZN(n652) );
  AND2_X1 U655 ( .A1(n586), .A2(n569), .ZN(n570) );
  AND2_X1 U656 ( .A1(n652), .A2(n570), .ZN(n571) );
  NAND2_X1 U657 ( .A1(n590), .A2(n571), .ZN(n630) );
  INV_X1 U658 ( .A(n630), .ZN(n572) );
  NOR2_X1 U659 ( .A1(n738), .A2(n572), .ZN(n574) );
  NAND2_X1 U660 ( .A1(n574), .A2(n573), .ZN(n576) );
  XNOR2_X1 U661 ( .A(n576), .B(n575), .ZN(n593) );
  NOR2_X1 U662 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U663 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U664 ( .A1(n582), .A2(n581), .ZN(n625) );
  XNOR2_X1 U665 ( .A(n583), .B(KEYINPUT31), .ZN(n642) );
  OR2_X1 U666 ( .A1(n625), .A2(n642), .ZN(n585) );
  NAND2_X1 U667 ( .A1(n585), .A2(n584), .ZN(n592) );
  AND2_X1 U668 ( .A1(n586), .A2(n649), .ZN(n587) );
  AND2_X1 U669 ( .A1(n588), .A2(n587), .ZN(n589) );
  AND2_X1 U670 ( .A1(n590), .A2(n589), .ZN(n623) );
  INV_X1 U671 ( .A(n623), .ZN(n591) );
  NAND2_X1 U672 ( .A1(n593), .A2(n400), .ZN(n595) );
  XNOR2_X1 U673 ( .A(KEYINPUT88), .B(KEYINPUT45), .ZN(n594) );
  NAND2_X1 U674 ( .A1(n687), .A2(n600), .ZN(n597) );
  XNOR2_X1 U675 ( .A(n597), .B(KEYINPUT87), .ZN(n599) );
  NAND2_X1 U676 ( .A1(n599), .A2(n598), .ZN(n602) );
  NAND2_X1 U677 ( .A1(n600), .A2(KEYINPUT2), .ZN(n601) );
  XOR2_X1 U678 ( .A(KEYINPUT91), .B(KEYINPUT59), .Z(n603) );
  XNOR2_X1 U679 ( .A(n604), .B(n603), .ZN(n605) );
  XNOR2_X1 U680 ( .A(n606), .B(n605), .ZN(n608) );
  INV_X1 U681 ( .A(G952), .ZN(n607) );
  INV_X1 U682 ( .A(n711), .ZN(n620) );
  NAND2_X1 U683 ( .A1(n608), .A2(n620), .ZN(n610) );
  XOR2_X1 U684 ( .A(KEYINPUT66), .B(KEYINPUT60), .Z(n609) );
  XNOR2_X1 U685 ( .A(n610), .B(n609), .ZN(G60) );
  XNOR2_X1 U686 ( .A(n611), .B(KEYINPUT122), .ZN(n612) );
  XNOR2_X1 U687 ( .A(n613), .B(n612), .ZN(n614) );
  INV_X1 U688 ( .A(KEYINPUT123), .ZN(n615) );
  XNOR2_X1 U689 ( .A(n616), .B(n615), .ZN(G66) );
  XOR2_X1 U690 ( .A(KEYINPUT62), .B(n617), .Z(n618) );
  XNOR2_X1 U691 ( .A(n619), .B(n618), .ZN(n621) );
  NAND2_X1 U692 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U693 ( .A(n622), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U694 ( .A(G101), .B(n623), .Z(G3) );
  NAND2_X1 U695 ( .A1(n625), .A2(n638), .ZN(n624) );
  XNOR2_X1 U696 ( .A(n624), .B(G104), .ZN(G6) );
  XOR2_X1 U697 ( .A(KEYINPUT27), .B(KEYINPUT111), .Z(n627) );
  NAND2_X1 U698 ( .A1(n625), .A2(n641), .ZN(n626) );
  XNOR2_X1 U699 ( .A(n627), .B(n626), .ZN(n629) );
  XOR2_X1 U700 ( .A(G107), .B(KEYINPUT26), .Z(n628) );
  XNOR2_X1 U701 ( .A(n629), .B(n628), .ZN(G9) );
  XNOR2_X1 U702 ( .A(G110), .B(n630), .ZN(G12) );
  XOR2_X1 U703 ( .A(KEYINPUT29), .B(KEYINPUT113), .Z(n632) );
  NAND2_X1 U704 ( .A1(n635), .A2(n641), .ZN(n631) );
  XNOR2_X1 U705 ( .A(n632), .B(n631), .ZN(n634) );
  XOR2_X1 U706 ( .A(G128), .B(KEYINPUT112), .Z(n633) );
  XNOR2_X1 U707 ( .A(n634), .B(n633), .ZN(G30) );
  NAND2_X1 U708 ( .A1(n635), .A2(n638), .ZN(n636) );
  XNOR2_X1 U709 ( .A(n636), .B(KEYINPUT114), .ZN(n637) );
  XNOR2_X1 U710 ( .A(G146), .B(n637), .ZN(G48) );
  XOR2_X1 U711 ( .A(G113), .B(KEYINPUT115), .Z(n640) );
  NAND2_X1 U712 ( .A1(n642), .A2(n638), .ZN(n639) );
  XNOR2_X1 U713 ( .A(n640), .B(n639), .ZN(G15) );
  NAND2_X1 U714 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U715 ( .A(n643), .B(G116), .ZN(G18) );
  XOR2_X1 U716 ( .A(G125), .B(KEYINPUT37), .Z(n644) );
  XNOR2_X1 U717 ( .A(n645), .B(n644), .ZN(G27) );
  XNOR2_X1 U718 ( .A(G134), .B(n646), .ZN(G36) );
  XNOR2_X1 U719 ( .A(n647), .B(G140), .ZN(n648) );
  XNOR2_X1 U720 ( .A(KEYINPUT116), .B(n648), .ZN(G42) );
  NOR2_X1 U721 ( .A1(n649), .A2(n402), .ZN(n650) );
  XNOR2_X1 U722 ( .A(n650), .B(KEYINPUT49), .ZN(n651) );
  NAND2_X1 U723 ( .A1(n652), .A2(n651), .ZN(n656) );
  XNOR2_X1 U724 ( .A(n654), .B(KEYINPUT50), .ZN(n655) );
  NOR2_X1 U725 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U726 ( .A(KEYINPUT117), .B(n657), .Z(n658) );
  NOR2_X1 U727 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U728 ( .A(KEYINPUT118), .B(n660), .Z(n661) );
  XNOR2_X1 U729 ( .A(n661), .B(KEYINPUT51), .ZN(n662) );
  NOR2_X1 U730 ( .A1(n680), .A2(n662), .ZN(n676) );
  BUF_X1 U731 ( .A(n663), .Z(n664) );
  NOR2_X1 U732 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U733 ( .A(KEYINPUT119), .B(n667), .Z(n668) );
  NOR2_X1 U734 ( .A1(n669), .A2(n668), .ZN(n673) );
  NOR2_X1 U735 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U736 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U737 ( .A1(n664), .A2(n674), .ZN(n675) );
  NOR2_X1 U738 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U739 ( .A(KEYINPUT52), .B(n677), .Z(n678) );
  NAND2_X1 U740 ( .A1(n679), .A2(n678), .ZN(n682) );
  OR2_X1 U741 ( .A1(n680), .A2(n664), .ZN(n681) );
  NAND2_X1 U742 ( .A1(n682), .A2(n681), .ZN(n693) );
  INV_X1 U743 ( .A(KEYINPUT2), .ZN(n685) );
  NAND2_X1 U744 ( .A1(n732), .A2(n685), .ZN(n686) );
  XNOR2_X1 U745 ( .A(n686), .B(KEYINPUT86), .ZN(n689) );
  OR2_X1 U746 ( .A1(n687), .A2(KEYINPUT2), .ZN(n688) );
  NAND2_X1 U747 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U748 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U749 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U750 ( .A1(n734), .A2(n694), .ZN(n695) );
  XOR2_X1 U751 ( .A(KEYINPUT53), .B(n695), .Z(G75) );
  XOR2_X1 U752 ( .A(KEYINPUT55), .B(KEYINPUT54), .Z(n697) );
  XNOR2_X1 U753 ( .A(KEYINPUT90), .B(KEYINPUT83), .ZN(n696) );
  XNOR2_X1 U754 ( .A(n697), .B(n696), .ZN(n699) );
  XNOR2_X1 U755 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n702) );
  XNOR2_X1 U756 ( .A(n700), .B(KEYINPUT57), .ZN(n701) );
  XNOR2_X1 U757 ( .A(n702), .B(n701), .ZN(n704) );
  NAND2_X1 U758 ( .A1(n706), .A2(G469), .ZN(n703) );
  XOR2_X1 U759 ( .A(n704), .B(n703), .Z(n705) );
  NOR2_X1 U760 ( .A1(n711), .A2(n705), .ZN(G54) );
  NAND2_X1 U761 ( .A1(n706), .A2(G478), .ZN(n709) );
  XOR2_X1 U762 ( .A(n707), .B(KEYINPUT121), .Z(n708) );
  XNOR2_X1 U763 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X1 U764 ( .A1(n711), .A2(n710), .ZN(G63) );
  NAND2_X1 U765 ( .A1(n687), .A2(n734), .ZN(n715) );
  NAND2_X1 U766 ( .A1(G953), .A2(G224), .ZN(n712) );
  XNOR2_X1 U767 ( .A(KEYINPUT61), .B(n712), .ZN(n713) );
  NAND2_X1 U768 ( .A1(n713), .A2(G898), .ZN(n714) );
  NAND2_X1 U769 ( .A1(n715), .A2(n714), .ZN(n723) );
  XNOR2_X1 U770 ( .A(n716), .B(KEYINPUT125), .ZN(n718) );
  XNOR2_X1 U771 ( .A(n718), .B(n717), .ZN(n719) );
  XNOR2_X1 U772 ( .A(n719), .B(G101), .ZN(n720) );
  NOR2_X1 U773 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U774 ( .A(n723), .B(n722), .ZN(n724) );
  XNOR2_X1 U775 ( .A(KEYINPUT124), .B(n724), .ZN(G69) );
  XOR2_X1 U776 ( .A(n726), .B(n725), .Z(n727) );
  XNOR2_X1 U777 ( .A(n728), .B(n727), .ZN(n733) );
  XNOR2_X1 U778 ( .A(KEYINPUT126), .B(n733), .ZN(n729) );
  XNOR2_X1 U779 ( .A(G227), .B(n729), .ZN(n730) );
  NAND2_X1 U780 ( .A1(n730), .A2(G900), .ZN(n731) );
  NAND2_X1 U781 ( .A1(n731), .A2(G953), .ZN(n737) );
  XNOR2_X1 U782 ( .A(n733), .B(n732), .ZN(n735) );
  NAND2_X1 U783 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U784 ( .A1(n737), .A2(n736), .ZN(G72) );
  BUF_X1 U785 ( .A(n738), .Z(n739) );
  XOR2_X1 U786 ( .A(n739), .B(G122), .Z(G24) );
  XOR2_X1 U787 ( .A(G131), .B(n740), .Z(G33) );
  XOR2_X1 U788 ( .A(G137), .B(n741), .Z(G39) );
endmodule

