//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 1 1 1 0 1 1 1 0 1 1 0 1 0 0 0 0 1 1 1 0 0 0 1 1 0 0 0 0 0 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n855, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931;
  INV_X1    g000(.A(KEYINPUT78), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n188));
  INV_X1    g002(.A(G107), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G104), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT77), .B1(new_n188), .B2(new_n190), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n189), .A2(G104), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n190), .B1(new_n192), .B2(KEYINPUT3), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT77), .ZN(new_n194));
  INV_X1    g008(.A(G104), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G107), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT3), .ZN(new_n197));
  AND2_X1   g011(.A1(new_n197), .A2(KEYINPUT76), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n197), .A2(KEYINPUT76), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n194), .B(new_n196), .C1(new_n198), .C2(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n191), .A2(new_n193), .A3(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G101), .ZN(new_n202));
  INV_X1    g016(.A(G101), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n191), .A2(new_n200), .A3(new_n203), .A4(new_n193), .ZN(new_n204));
  AND3_X1   g018(.A1(new_n202), .A2(KEYINPUT4), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT4), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n201), .A2(new_n206), .A3(G101), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G143), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n210), .B1(new_n211), .B2(G146), .ZN(new_n212));
  NOR3_X1   g026(.A1(new_n208), .A2(KEYINPUT64), .A3(G143), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n209), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  XOR2_X1   g028(.A(KEYINPUT0), .B(G128), .Z(new_n215));
  NAND2_X1  g029(.A1(new_n211), .A2(G146), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n209), .A2(new_n216), .A3(G128), .ZN(new_n217));
  AOI22_X1  g031(.A1(new_n214), .A2(new_n215), .B1(new_n217), .B2(KEYINPUT0), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n207), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n187), .B1(new_n205), .B2(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(G101), .B1(new_n196), .B2(new_n192), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n204), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT1), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n209), .A2(new_n216), .A3(new_n224), .A4(G128), .ZN(new_n225));
  INV_X1    g039(.A(new_n209), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n216), .A2(KEYINPUT64), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n210), .A2(new_n211), .A3(G146), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G128), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n230), .B1(new_n209), .B2(KEYINPUT1), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n225), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n232), .A2(KEYINPUT10), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n209), .A2(new_n216), .ZN(new_n234));
  OAI211_X1 g048(.A(KEYINPUT79), .B(KEYINPUT1), .C1(new_n211), .C2(G146), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G128), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT79), .B1(new_n209), .B2(KEYINPUT1), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n234), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n225), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(new_n204), .A3(new_n221), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT10), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n223), .A2(new_n233), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n202), .A2(KEYINPUT4), .A3(new_n204), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n243), .A2(KEYINPUT78), .A3(new_n218), .A4(new_n207), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n220), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT11), .ZN(new_n246));
  INV_X1    g060(.A(G134), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n246), .B1(new_n247), .B2(G137), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(G137), .ZN(new_n249));
  INV_X1    g063(.A(G137), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(KEYINPUT11), .A3(G134), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n248), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G131), .ZN(new_n253));
  INV_X1    g067(.A(G131), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n248), .A2(new_n251), .A3(new_n254), .A4(new_n249), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n245), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(G110), .B(G140), .ZN(new_n258));
  INV_X1    g072(.A(G953), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G227), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n258), .B(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n262));
  XOR2_X1   g076(.A(new_n261), .B(new_n262), .Z(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n256), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n220), .A2(new_n265), .A3(new_n242), .A4(new_n244), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n266), .A2(KEYINPUT80), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(KEYINPUT80), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n257), .B(new_n264), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT81), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n222), .B(new_n225), .C1(new_n231), .C2(new_n229), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n265), .B1(new_n271), .B2(new_n240), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT12), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n272), .B(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n244), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n207), .A2(new_n218), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT78), .B1(new_n276), .B2(new_n243), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT80), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n278), .A2(new_n279), .A3(new_n265), .A4(new_n242), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n266), .A2(KEYINPUT80), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n274), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n269), .B(new_n270), .C1(new_n264), .C2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n266), .B(new_n279), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n263), .B1(new_n285), .B2(new_n274), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n270), .B1(new_n286), .B2(new_n269), .ZN(new_n287));
  OAI21_X1  g101(.A(G469), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT82), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n280), .A2(new_n281), .B1(new_n256), .B2(new_n245), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n289), .B1(new_n290), .B2(new_n264), .ZN(new_n291));
  INV_X1    g105(.A(new_n257), .ZN(new_n292));
  OAI211_X1 g106(.A(KEYINPUT82), .B(new_n263), .C1(new_n285), .C2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n274), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n294), .B(new_n264), .C1(new_n267), .C2(new_n268), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n291), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G469), .ZN(new_n297));
  INV_X1    g111(.A(G902), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(G469), .A2(G902), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n288), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  XOR2_X1   g115(.A(KEYINPUT9), .B(G234), .Z(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(G221), .B1(new_n303), .B2(G902), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT83), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n301), .A2(KEYINPUT83), .A3(new_n304), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G472), .ZN(new_n310));
  INV_X1    g124(.A(new_n249), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n247), .A2(G137), .ZN(new_n312));
  OAI21_X1  g126(.A(G131), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n232), .A2(new_n255), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT30), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n218), .A2(new_n256), .ZN(new_n316));
  AND3_X1   g130(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT66), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n218), .A2(new_n318), .A3(new_n256), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n318), .B1(new_n218), .B2(new_n256), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n314), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n317), .B1(new_n321), .B2(KEYINPUT30), .ZN(new_n322));
  XOR2_X1   g136(.A(KEYINPUT2), .B(G113), .Z(new_n323));
  XNOR2_X1  g137(.A(G116), .B(G119), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT65), .ZN(new_n326));
  OR2_X1    g140(.A1(new_n323), .A2(new_n324), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n326), .B(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT67), .B1(new_n322), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT67), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n316), .A2(KEYINPUT66), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n218), .A2(new_n318), .A3(new_n256), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n315), .B1(new_n334), .B2(new_n314), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n331), .B(new_n328), .C1(new_n335), .C2(new_n317), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n334), .A2(new_n329), .A3(new_n314), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n330), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n339), .B(G101), .ZN(new_n340));
  INV_X1    g154(.A(G237), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(new_n259), .A3(G210), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n340), .B(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n338), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT29), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n314), .A2(new_n316), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n328), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT28), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n349), .B1(new_n347), .B2(new_n328), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n348), .B(new_n350), .C1(new_n337), .C2(new_n349), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n345), .B(new_n346), .C1(new_n344), .C2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n350), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n321), .A2(new_n328), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n337), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n353), .B1(new_n355), .B2(KEYINPUT28), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n344), .A2(new_n346), .ZN(new_n357));
  AOI21_X1  g171(.A(G902), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n310), .B1(new_n352), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n351), .A2(new_n344), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT69), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n360), .B(new_n361), .ZN(new_n362));
  AND4_X1   g176(.A1(new_n343), .A2(new_n330), .A3(new_n336), .A4(new_n337), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(KEYINPUT68), .A3(KEYINPUT31), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT31), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n330), .A2(new_n336), .A3(new_n343), .A4(new_n337), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT68), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n362), .B1(new_n364), .B2(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(G472), .A2(G902), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(KEYINPUT32), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n360), .B(KEYINPUT69), .ZN(new_n373));
  AOI21_X1  g187(.A(KEYINPUT31), .B1(new_n363), .B2(KEYINPUT68), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n366), .A2(new_n367), .A3(new_n365), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT32), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(new_n377), .A3(new_n370), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n359), .B1(new_n372), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(G125), .B(G140), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n208), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT71), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n381), .B(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G125), .ZN(new_n384));
  NOR3_X1   g198(.A1(new_n384), .A2(KEYINPUT16), .A3(G140), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n385), .B1(new_n380), .B2(KEYINPUT16), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G146), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT23), .ZN(new_n388));
  INV_X1    g202(.A(G119), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n388), .B1(new_n389), .B2(G128), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n230), .A2(KEYINPUT23), .A3(G119), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n390), .B(new_n391), .C1(G119), .C2(new_n230), .ZN(new_n392));
  XNOR2_X1  g206(.A(G119), .B(G128), .ZN(new_n393));
  XOR2_X1   g207(.A(KEYINPUT24), .B(G110), .Z(new_n394));
  OAI22_X1  g208(.A1(new_n392), .A2(G110), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n383), .A2(new_n387), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT72), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n392), .A2(G110), .B1(new_n393), .B2(new_n394), .ZN(new_n399));
  INV_X1    g213(.A(new_n387), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n386), .A2(G146), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n383), .A2(KEYINPUT72), .A3(new_n387), .A4(new_n395), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n398), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n259), .A2(G221), .A3(G234), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n405), .B(KEYINPUT22), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n406), .B(G137), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n398), .A2(new_n402), .A3(new_n403), .A4(new_n407), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT25), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(new_n412), .A3(new_n298), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n409), .A2(new_n410), .ZN(new_n414));
  OAI21_X1  g228(.A(KEYINPUT25), .B1(new_n414), .B2(G902), .ZN(new_n415));
  INV_X1    g229(.A(G217), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n416), .B1(G234), .B2(new_n298), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n417), .B(KEYINPUT70), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n413), .A2(new_n415), .A3(new_n418), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n417), .A2(G902), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n409), .A2(new_n410), .A3(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n421), .B(KEYINPUT73), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n379), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(G214), .B1(G237), .B2(G902), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  XOR2_X1   g240(.A(G110), .B(G122), .Z(new_n427));
  XOR2_X1   g241(.A(new_n427), .B(KEYINPUT8), .Z(new_n428));
  NAND2_X1  g242(.A1(new_n389), .A2(G116), .ZN(new_n429));
  OAI21_X1  g243(.A(G113), .B1(new_n429), .B2(KEYINPUT5), .ZN(new_n430));
  XOR2_X1   g244(.A(new_n430), .B(KEYINPUT85), .Z(new_n431));
  NAND2_X1  g245(.A1(new_n324), .A2(KEYINPUT5), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n223), .A2(new_n433), .A3(new_n325), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n434), .B(KEYINPUT86), .ZN(new_n435));
  INV_X1    g249(.A(new_n430), .ZN(new_n436));
  AOI22_X1  g250(.A1(new_n436), .A2(new_n432), .B1(new_n324), .B2(new_n323), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n223), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n428), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  OR2_X1    g253(.A1(new_n232), .A2(G125), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n218), .A2(new_n384), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT84), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NOR3_X1   g258(.A1(new_n218), .A2(KEYINPUT84), .A3(new_n384), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n441), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G224), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n447), .A2(G953), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n449), .A2(KEYINPUT7), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n449), .A2(KEYINPUT87), .ZN(new_n451));
  OR3_X1    g265(.A1(new_n446), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n328), .A2(new_n243), .A3(new_n207), .ZN(new_n453));
  INV_X1    g267(.A(new_n427), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n223), .A2(new_n437), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n450), .B1(new_n446), .B2(new_n451), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n439), .A2(new_n452), .A3(new_n456), .A4(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n446), .B(new_n449), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n453), .A2(new_n455), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT6), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n461), .A3(new_n427), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n427), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n463), .A2(KEYINPUT6), .A3(new_n456), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n459), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n458), .A2(new_n465), .A3(new_n298), .ZN(new_n466));
  OAI21_X1  g280(.A(G210), .B1(G237), .B2(G902), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n458), .A2(new_n465), .A3(new_n298), .A4(new_n467), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n426), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(G475), .A2(G902), .ZN(new_n473));
  XNOR2_X1  g287(.A(G113), .B(G122), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(new_n195), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n341), .A2(new_n259), .A3(G214), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(new_n211), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G131), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n477), .B(G143), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n254), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n387), .ZN(new_n483));
  NAND2_X1  g297(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n380), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n485), .B(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n483), .B1(new_n208), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n383), .B1(new_n208), .B2(new_n380), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT18), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n490), .A2(new_n254), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n480), .B(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n476), .B1(new_n488), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT89), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n496), .B1(new_n400), .B2(new_n401), .ZN(new_n497));
  INV_X1    g311(.A(new_n401), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(KEYINPUT89), .A3(new_n387), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n478), .A2(KEYINPUT17), .A3(G131), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT17), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n479), .A2(new_n481), .A3(new_n501), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n497), .A2(new_n499), .A3(new_n500), .A4(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(new_n475), .A3(new_n493), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n495), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n505), .A2(KEYINPUT90), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT90), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n507), .B1(new_n495), .B2(new_n504), .ZN(new_n508));
  OAI211_X1 g322(.A(KEYINPUT20), .B(new_n473), .C1(new_n506), .C2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n504), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n475), .B1(new_n503), .B2(new_n493), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n298), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT92), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT91), .B(G475), .ZN(new_n515));
  OAI211_X1 g329(.A(KEYINPUT92), .B(new_n298), .C1(new_n510), .C2(new_n511), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n505), .A2(new_n473), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT20), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n509), .A2(new_n517), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n259), .A2(G952), .ZN(new_n523));
  NAND2_X1  g337(.A1(G234), .A2(G237), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  XOR2_X1   g340(.A(KEYINPUT21), .B(G898), .Z(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n524), .A2(G902), .A3(G953), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n526), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(G478), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(KEYINPUT15), .ZN(new_n534));
  NOR3_X1   g348(.A1(new_n303), .A2(new_n416), .A3(G953), .ZN(new_n535));
  XNOR2_X1  g349(.A(G128), .B(G143), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(G134), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(KEYINPUT93), .ZN(new_n538));
  XNOR2_X1  g352(.A(G116), .B(G122), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n189), .ZN(new_n540));
  INV_X1    g354(.A(G116), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n541), .A2(KEYINPUT14), .A3(G122), .ZN(new_n542));
  INV_X1    g356(.A(new_n539), .ZN(new_n543));
  OAI211_X1 g357(.A(G107), .B(new_n542), .C1(new_n543), .C2(KEYINPUT14), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n538), .A2(new_n540), .A3(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n539), .B(new_n189), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n230), .A2(KEYINPUT13), .A3(G143), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n547), .B1(new_n536), .B2(KEYINPUT13), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(G134), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n536), .A2(new_n247), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n546), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n535), .B1(new_n545), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n545), .A2(new_n551), .A3(new_n535), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n298), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT94), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n534), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n557), .ZN(new_n559));
  AOI21_X1  g373(.A(G902), .B1(new_n553), .B2(new_n554), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT94), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n558), .B1(new_n562), .B2(new_n534), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n522), .A2(new_n532), .A3(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n472), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n309), .A2(new_n424), .A3(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(G101), .ZN(G3));
  NAND2_X1  g381(.A1(new_n471), .A2(new_n532), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT33), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n555), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT95), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n552), .B(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT96), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n554), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n545), .A2(KEYINPUT96), .A3(new_n551), .A4(new_n535), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(KEYINPUT33), .A3(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n570), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n298), .A2(G478), .ZN(new_n578));
  OAI22_X1  g392(.A1(new_n577), .A2(new_n578), .B1(G478), .B2(new_n560), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n521), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n568), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(G472), .B1(new_n369), .B2(G902), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n583), .B1(new_n371), .B2(new_n369), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n584), .A2(new_n423), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n309), .A2(new_n582), .A3(new_n585), .ZN(new_n586));
  XOR2_X1   g400(.A(KEYINPUT34), .B(G104), .Z(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(KEYINPUT97), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n586), .B(new_n588), .ZN(G6));
  AND2_X1   g403(.A1(new_n509), .A2(new_n517), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n506), .A2(new_n508), .ZN(new_n591));
  INV_X1    g405(.A(new_n473), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n519), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n568), .A2(new_n563), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n309), .A2(new_n585), .A3(new_n595), .ZN(new_n596));
  XOR2_X1   g410(.A(KEYINPUT35), .B(G107), .Z(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(G9));
  XNOR2_X1  g412(.A(new_n404), .B(KEYINPUT98), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n408), .A2(KEYINPUT36), .ZN(new_n600));
  XOR2_X1   g414(.A(new_n599), .B(new_n600), .Z(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n420), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n419), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n584), .A2(new_n604), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n301), .A2(KEYINPUT83), .A3(new_n304), .ZN(new_n606));
  AOI21_X1  g420(.A(KEYINPUT83), .B1(new_n301), .B2(new_n304), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n565), .B(new_n605), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  XOR2_X1   g422(.A(new_n608), .B(KEYINPUT37), .Z(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G110), .ZN(G12));
  INV_X1    g424(.A(new_n359), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n377), .B1(new_n376), .B2(new_n370), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n369), .A2(KEYINPUT32), .A3(new_n371), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n525), .B1(G900), .B2(new_n529), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n590), .A2(new_n593), .A3(new_n615), .ZN(new_n616));
  NOR4_X1   g430(.A1(new_n472), .A2(new_n604), .A3(new_n616), .A4(new_n563), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n614), .B(new_n617), .C1(new_n606), .C2(new_n607), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G128), .ZN(G30));
  XOR2_X1   g433(.A(new_n615), .B(KEYINPUT39), .Z(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n309), .A2(new_n621), .ZN(new_n622));
  OR2_X1    g436(.A1(new_n622), .A2(KEYINPUT40), .ZN(new_n623));
  INV_X1    g437(.A(new_n563), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n521), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n622), .B2(KEYINPUT40), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n372), .A2(new_n378), .ZN(new_n627));
  INV_X1    g441(.A(new_n355), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n366), .B1(new_n343), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n310), .B1(new_n629), .B2(new_n298), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n603), .B1(new_n627), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n469), .A2(new_n470), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT38), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n623), .A2(new_n626), .A3(new_n425), .A4(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G143), .ZN(G45));
  AND3_X1   g451(.A1(new_n521), .A2(new_n579), .A3(new_n615), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n471), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n379), .A2(new_n604), .A3(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n640), .B1(new_n606), .B2(new_n607), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT99), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(new_n208), .ZN(G48));
  AND3_X1   g457(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n297), .B1(new_n296), .B2(new_n298), .ZN(new_n645));
  INV_X1    g459(.A(new_n304), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n424), .A2(new_n582), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT41), .B(G113), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G15));
  NAND3_X1  g464(.A1(new_n424), .A2(new_n595), .A3(new_n647), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G116), .ZN(G18));
  NOR2_X1   g466(.A1(new_n644), .A2(new_n645), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT100), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n653), .A2(new_n654), .A3(new_n304), .A4(new_n471), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n296), .A2(new_n298), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(G469), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n657), .A2(new_n304), .A3(new_n299), .A4(new_n471), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(KEYINPUT100), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n564), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n379), .A2(new_n604), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G119), .ZN(G21));
  OAI22_X1  g478(.A1(new_n374), .A2(new_n375), .B1(new_n343), .B2(new_n356), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n370), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT101), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n423), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(KEYINPUT101), .B1(new_n419), .B2(new_n422), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n583), .A2(new_n666), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(KEYINPUT102), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT102), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n583), .A2(new_n666), .A3(new_n670), .A4(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n568), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n657), .A2(new_n304), .A3(new_n299), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n677), .A2(new_n625), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n675), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G122), .ZN(G24));
  NAND4_X1  g494(.A1(new_n583), .A2(new_n666), .A3(new_n638), .A4(new_n603), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n681), .B1(new_n655), .B2(new_n659), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT103), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G125), .ZN(G27));
  NAND2_X1  g498(.A1(new_n286), .A2(new_n269), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n299), .B(new_n300), .C1(new_n297), .C2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n304), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n687), .A2(new_n379), .A3(new_n423), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n689));
  INV_X1    g503(.A(new_n638), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n469), .A2(new_n425), .A3(new_n470), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n688), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n692), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n614), .A2(KEYINPUT104), .A3(new_n670), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n696));
  INV_X1    g510(.A(new_n670), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n696), .B1(new_n379), .B2(new_n697), .ZN(new_n698));
  AOI211_X1 g512(.A(new_n687), .B(new_n694), .C1(new_n695), .C2(new_n698), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n693), .B1(new_n699), .B2(new_n689), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n254), .ZN(G33));
  INV_X1    g515(.A(new_n616), .ZN(new_n702));
  INV_X1    g516(.A(new_n691), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n688), .A2(new_n624), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G134), .ZN(G36));
  AOI21_X1  g519(.A(KEYINPUT105), .B1(new_n522), .B2(new_n579), .ZN(new_n706));
  XOR2_X1   g520(.A(new_n706), .B(KEYINPUT43), .Z(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(new_n584), .A3(new_n603), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n703), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT106), .ZN(new_n711));
  OR3_X1    g525(.A1(new_n284), .A2(new_n287), .A3(KEYINPUT45), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT45), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n712), .B(G469), .C1(new_n713), .C2(new_n685), .ZN(new_n714));
  AOI21_X1  g528(.A(KEYINPUT46), .B1(new_n714), .B2(new_n300), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n715), .A2(new_n644), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(KEYINPUT46), .A3(new_n300), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n646), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n718), .A2(new_n621), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n708), .A2(new_n709), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n711), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G137), .ZN(G39));
  XOR2_X1   g536(.A(new_n718), .B(KEYINPUT47), .Z(new_n723));
  NAND3_X1  g537(.A1(new_n692), .A2(new_n379), .A3(new_n423), .ZN(new_n724));
  XOR2_X1   g538(.A(new_n724), .B(KEYINPUT107), .Z(new_n725));
  OR2_X1    g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G140), .ZN(G42));
  INV_X1    g541(.A(new_n653), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n627), .B(new_n631), .C1(new_n728), .C2(KEYINPUT49), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n728), .A2(KEYINPUT49), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n522), .A2(new_n579), .ZN(new_n731));
  NOR4_X1   g545(.A1(new_n729), .A2(new_n730), .A3(new_n634), .A4(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n732), .A2(new_n304), .A3(new_n425), .A4(new_n670), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n707), .A2(new_n526), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n734), .B1(new_n674), .B2(new_n672), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n660), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n723), .B1(new_n304), .B2(new_n728), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n737), .A2(new_n703), .A3(new_n735), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n647), .A2(new_n703), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n627), .A2(new_n631), .ZN(new_n740));
  NOR4_X1   g554(.A1(new_n739), .A2(new_n423), .A3(new_n740), .A4(new_n525), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n522), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n742), .A2(new_n579), .ZN(new_n743));
  NOR2_X1   g557(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n734), .A2(new_n739), .ZN(new_n745));
  AND4_X1   g559(.A1(new_n583), .A2(new_n745), .A3(new_n603), .A4(new_n666), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n634), .A2(new_n425), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n735), .A2(new_n647), .A3(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n748), .A2(new_n749), .ZN(new_n751));
  AOI211_X1 g565(.A(new_n744), .B(new_n746), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n738), .A2(new_n743), .A3(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT112), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT51), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n738), .A2(new_n757), .A3(new_n743), .A4(new_n752), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n756), .A2(new_n523), .A3(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n563), .A2(new_n521), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n568), .A2(new_n761), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n585), .B(new_n762), .C1(new_n606), .C2(new_n607), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT109), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n608), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n586), .ZN(new_n766));
  INV_X1    g580(.A(new_n566), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n764), .B1(new_n608), .B2(new_n763), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n693), .B(new_n704), .C1(new_n699), .C2(new_n689), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n703), .A2(new_n603), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n309), .A2(new_n614), .A3(new_n563), .A4(new_n702), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n686), .A2(new_n304), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n773), .A2(new_n583), .A3(new_n638), .A4(new_n666), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n771), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n770), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n639), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n614), .A2(new_n603), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n778), .B1(new_n307), .B2(new_n308), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n682), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n472), .A2(new_n625), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n773), .A2(new_n615), .A3(new_n632), .A4(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n780), .A2(KEYINPUT52), .A3(new_n618), .A4(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n681), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n654), .B1(new_n647), .B2(new_n471), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n658), .A2(KEYINPUT100), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n787), .A2(new_n618), .A3(new_n641), .A4(new_n782), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n783), .A2(new_n790), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n679), .A2(new_n648), .A3(new_n651), .ZN(new_n793));
  OAI21_X1  g607(.A(KEYINPUT108), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n568), .B1(new_n672), .B2(new_n674), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n677), .A2(new_n379), .A3(new_n423), .ZN(new_n796));
  AOI22_X1  g610(.A1(new_n795), .A2(new_n678), .B1(new_n796), .B2(new_n595), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT108), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n797), .A2(new_n663), .A3(new_n798), .A4(new_n648), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n794), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n769), .A2(new_n776), .A3(new_n791), .A4(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT53), .B1(new_n791), .B2(KEYINPUT110), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(KEYINPUT54), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n792), .A2(new_n793), .A3(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n769), .A2(new_n776), .A3(new_n791), .A4(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT111), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n801), .A2(new_n809), .A3(new_n806), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n809), .B1(new_n801), .B2(new_n806), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n805), .B(new_n808), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n804), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n759), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n741), .A2(new_n580), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n695), .A2(new_n698), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n745), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(KEYINPUT48), .ZN(new_n818));
  AND4_X1   g632(.A1(new_n736), .A2(new_n814), .A3(new_n815), .A4(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(G952), .A2(G953), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n733), .B1(new_n819), .B2(new_n820), .ZN(G75));
  OAI21_X1  g635(.A(new_n808), .B1(new_n810), .B2(new_n811), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n822), .A2(G210), .A3(G902), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT56), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(KEYINPUT114), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n464), .A2(new_n462), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(new_n459), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT113), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT55), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n259), .A2(G952), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n825), .A2(new_n829), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n830), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT115), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n830), .A2(KEYINPUT115), .A3(new_n832), .A4(new_n833), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(G51));
  NAND2_X1  g652(.A1(new_n822), .A2(KEYINPUT54), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n839), .A2(KEYINPUT116), .A3(new_n812), .ZN(new_n840));
  INV_X1    g654(.A(new_n822), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n841), .A2(new_n842), .A3(new_n805), .ZN(new_n843));
  XOR2_X1   g657(.A(new_n300), .B(KEYINPUT57), .Z(new_n844));
  NAND3_X1  g658(.A1(new_n840), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT117), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n840), .A2(new_n843), .A3(new_n847), .A4(new_n844), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n296), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n841), .A2(new_n298), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n714), .B(KEYINPUT118), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n831), .B1(new_n850), .B2(new_n853), .ZN(G54));
  NAND3_X1  g668(.A1(new_n851), .A2(KEYINPUT58), .A3(G475), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n855), .A2(new_n591), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n855), .A2(new_n591), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n856), .A2(new_n857), .A3(new_n831), .ZN(G60));
  NOR2_X1   g672(.A1(new_n572), .A2(new_n576), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n859), .B1(new_n569), .B2(new_n555), .ZN(new_n860));
  NAND2_X1  g674(.A1(G478), .A2(G902), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(KEYINPUT59), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n840), .A2(new_n843), .A3(new_n860), .A4(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n863), .A2(new_n864), .A3(new_n832), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n864), .B1(new_n863), .B2(new_n832), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n860), .B1(new_n813), .B2(new_n862), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(G63));
  NAND2_X1  g682(.A1(G217), .A2(G902), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT60), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n841), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n831), .B1(new_n872), .B2(new_n414), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT61), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n871), .A2(new_n601), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n873), .B(new_n876), .C1(new_n874), .C2(KEYINPUT61), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(G66));
  NAND2_X1  g694(.A1(new_n769), .A2(new_n800), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n259), .ZN(new_n882));
  OAI21_X1  g696(.A(G953), .B1(new_n528), .B2(new_n447), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n826), .B1(G898), .B2(new_n259), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n884), .B(new_n885), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT121), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(KEYINPUT122), .Z(G69));
  XOR2_X1   g702(.A(new_n322), .B(new_n487), .Z(new_n889));
  NAND2_X1  g703(.A1(G900), .A2(G953), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n726), .A2(new_n721), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n780), .A2(new_n618), .ZN(new_n892));
  INV_X1    g706(.A(new_n770), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n719), .A2(new_n816), .A3(new_n781), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n891), .A2(new_n892), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n889), .B(new_n890), .C1(new_n895), .C2(G953), .ZN(new_n896));
  INV_X1    g710(.A(new_n622), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n761), .A2(new_n581), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n897), .A2(new_n424), .A3(new_n703), .A4(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n636), .A2(new_n892), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT62), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n901), .A2(new_n902), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n900), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(G953), .B1(new_n891), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n896), .B1(new_n907), .B2(new_n889), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n259), .B1(G227), .B2(G900), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n907), .A2(new_n889), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n911), .A2(KEYINPUT123), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(KEYINPUT123), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n912), .A2(new_n896), .A3(new_n913), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n909), .B(KEYINPUT124), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n910), .B1(new_n914), .B2(new_n915), .ZN(G72));
  NAND2_X1  g730(.A1(G472), .A2(G902), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT63), .Z(new_n918));
  OAI21_X1  g732(.A(new_n918), .B1(new_n895), .B2(new_n881), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n338), .B(KEYINPUT125), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n920), .A2(new_n343), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT126), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n891), .A2(new_n906), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n918), .B1(new_n924), .B2(new_n881), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n925), .A2(new_n343), .A3(new_n920), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n345), .A2(new_n366), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n918), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(KEYINPUT127), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n928), .A2(KEYINPUT127), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n803), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  AND4_X1   g745(.A1(new_n832), .A2(new_n923), .A3(new_n926), .A4(new_n931), .ZN(G57));
endmodule


