//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 1 0 0 0 0 0 0 0 1 1 0 0 1 1 0 0 0 0 0 0 1 1 0 1 1 0 1 0 0 1 0 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(G113), .B(G122), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(G104), .ZN(new_n189));
  OR2_X1    g003(.A1(KEYINPUT68), .A2(G237), .ZN(new_n190));
  NAND2_X1  g004(.A1(KEYINPUT68), .A2(G237), .ZN(new_n191));
  AOI21_X1  g005(.A(G953), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(G143), .A3(G214), .ZN(new_n193));
  INV_X1    g007(.A(G953), .ZN(new_n194));
  AND2_X1   g008(.A1(KEYINPUT68), .A2(G237), .ZN(new_n195));
  NOR2_X1   g009(.A1(KEYINPUT68), .A2(G237), .ZN(new_n196));
  OAI211_X1 g010(.A(G214), .B(new_n194), .C1(new_n195), .C2(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n193), .A2(new_n199), .ZN(new_n200));
  AND2_X1   g014(.A1(KEYINPUT18), .A2(G131), .ZN(new_n201));
  OR2_X1    g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(G125), .B(G140), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XOR2_X1   g019(.A(G125), .B(G140), .Z(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G146), .ZN(new_n207));
  AOI22_X1  g021(.A1(new_n200), .A2(new_n201), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT91), .B1(new_n200), .B2(G131), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT17), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT91), .ZN(new_n211));
  INV_X1    g025(.A(G131), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n193), .A2(new_n199), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n200), .A2(G131), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n209), .A2(new_n210), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT16), .ZN(new_n217));
  INV_X1    g031(.A(G140), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT74), .A4(G125), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n217), .A2(new_n218), .A3(G125), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT74), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n216), .A2(new_n219), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n204), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n216), .A2(G146), .A3(new_n219), .A4(new_n222), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI211_X1 g040(.A(new_n210), .B(new_n212), .C1(new_n193), .C2(new_n199), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI221_X4 g042(.A(new_n189), .B1(new_n202), .B2(new_n208), .C1(new_n215), .C2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n189), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n215), .A2(new_n228), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n202), .A2(new_n208), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n187), .B1(new_n229), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT93), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT93), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n236), .B(new_n187), .C1(new_n229), .C2(new_n233), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n235), .A2(G475), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT20), .ZN(new_n239));
  NOR2_X1   g053(.A1(G475), .A2(G902), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n209), .A2(new_n213), .A3(new_n214), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n203), .B(KEYINPUT19), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n204), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n241), .A2(new_n225), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n230), .B1(new_n244), .B2(new_n232), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n239), .B(new_n240), .C1(new_n229), .C2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT92), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n240), .B1(new_n229), .B2(new_n245), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT90), .B(KEYINPUT20), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n246), .A2(KEYINPUT92), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n238), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT96), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT94), .B(G122), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G116), .ZN(new_n257));
  INV_X1    g071(.A(G107), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT95), .ZN(new_n259));
  INV_X1    g073(.A(G122), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n259), .B1(new_n260), .B2(G116), .ZN(new_n261));
  INV_X1    g075(.A(G116), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n262), .A2(KEYINPUT95), .A3(G122), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n257), .A2(new_n258), .A3(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G143), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT64), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT64), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G143), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n267), .A2(new_n269), .A3(G128), .ZN(new_n270));
  INV_X1    g084(.A(G134), .ZN(new_n271));
  INV_X1    g085(.A(G128), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G143), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n270), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n271), .B1(new_n270), .B2(new_n273), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n265), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AOI22_X1  g091(.A1(new_n264), .A2(KEYINPUT14), .B1(new_n256), .B2(G116), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT14), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n261), .A2(new_n279), .A3(new_n263), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n258), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n255), .B1(new_n277), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n264), .A2(KEYINPUT14), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n283), .A2(new_n280), .A3(new_n257), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G107), .ZN(new_n285));
  INV_X1    g099(.A(new_n276), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n274), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n285), .A2(new_n287), .A3(KEYINPUT96), .A4(new_n265), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n270), .A2(KEYINPUT13), .A3(new_n273), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n289), .B(G134), .C1(KEYINPUT13), .C2(new_n270), .ZN(new_n290));
  INV_X1    g104(.A(new_n265), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n258), .B1(new_n257), .B2(new_n264), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n290), .B(new_n274), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n282), .A2(new_n288), .A3(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT9), .B(G234), .ZN(new_n295));
  INV_X1    g109(.A(G217), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n295), .A2(new_n296), .A3(G953), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n282), .A2(new_n288), .A3(new_n293), .A4(new_n297), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n187), .ZN(new_n302));
  INV_X1    g116(.A(G478), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n303), .A2(KEYINPUT15), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n302), .A2(new_n304), .ZN(new_n306));
  OR2_X1    g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n254), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G952), .ZN(new_n309));
  AOI211_X1 g123(.A(G953), .B(new_n309), .C1(G234), .C2(G237), .ZN(new_n310));
  AOI211_X1 g124(.A(new_n187), .B(new_n194), .C1(G234), .C2(G237), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT21), .B(G898), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n308), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(G214), .B1(G237), .B2(G902), .ZN(new_n316));
  INV_X1    g130(.A(G104), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT3), .B1(new_n317), .B2(G107), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT3), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(new_n258), .A3(G104), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G101), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT77), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT77), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G101), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n317), .A2(G107), .ZN(new_n326));
  AND3_X1   g140(.A1(new_n323), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT78), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n321), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n318), .A2(new_n320), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n323), .A2(new_n325), .A3(new_n326), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT78), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT79), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n333), .B1(new_n317), .B2(G107), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n258), .A2(KEYINPUT79), .A3(G104), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(new_n326), .A3(new_n335), .ZN(new_n336));
  AOI22_X1  g150(.A1(new_n329), .A2(new_n332), .B1(G101), .B2(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n262), .A2(G119), .ZN(new_n338));
  INV_X1    g152(.A(G119), .ZN(new_n339));
  OAI21_X1  g153(.A(KEYINPUT66), .B1(new_n339), .B2(G116), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT66), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(new_n262), .A3(G119), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n338), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT5), .ZN(new_n344));
  INV_X1    g158(.A(G113), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT5), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n345), .B1(new_n338), .B2(new_n346), .ZN(new_n347));
  AND2_X1   g161(.A1(KEYINPUT2), .A2(G113), .ZN(new_n348));
  NOR2_X1   g162(.A1(KEYINPUT2), .A2(G113), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n344), .A2(new_n347), .B1(new_n343), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n337), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT4), .ZN(new_n353));
  AOI211_X1 g167(.A(new_n353), .B(new_n322), .C1(new_n321), .C2(new_n326), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n328), .B1(new_n321), .B2(new_n327), .ZN(new_n355));
  NOR3_X1   g169(.A1(new_n330), .A2(new_n331), .A3(KEYINPUT78), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT4), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n322), .B1(new_n321), .B2(new_n326), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n354), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n340), .A2(new_n342), .ZN(new_n361));
  INV_X1    g175(.A(new_n338), .ZN(new_n362));
  AND3_X1   g176(.A1(new_n361), .A2(new_n350), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n350), .B1(new_n361), .B2(new_n362), .ZN(new_n364));
  OAI21_X1  g178(.A(KEYINPUT67), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n361), .A2(new_n362), .ZN(new_n366));
  INV_X1    g180(.A(new_n350), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT67), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n343), .A2(new_n350), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n352), .B1(new_n360), .B2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(G110), .B(G122), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n352), .B(new_n374), .C1(new_n360), .C2(new_n372), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(KEYINPUT6), .A3(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n204), .A2(G143), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n380), .B1(new_n198), .B2(G146), .ZN(new_n381));
  AND2_X1   g195(.A1(KEYINPUT0), .A2(G128), .ZN(new_n382));
  NOR2_X1   g196(.A1(KEYINPUT0), .A2(G128), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n204), .A2(G143), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n386), .B1(new_n198), .B2(G146), .ZN(new_n387));
  AOI22_X1  g201(.A1(new_n381), .A2(new_n384), .B1(new_n387), .B2(new_n382), .ZN(new_n388));
  INV_X1    g202(.A(G125), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT83), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(G146), .B1(new_n267), .B2(new_n269), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n384), .B1(new_n391), .B2(new_n379), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n267), .A2(new_n269), .A3(G146), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(new_n385), .A3(new_n382), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n389), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT83), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n272), .B1(new_n385), .B2(KEYINPUT1), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n381), .A2(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n272), .A2(KEYINPUT1), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n393), .A2(new_n385), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n400), .A2(new_n389), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n390), .A2(new_n397), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G224), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n405), .A2(G953), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n404), .B(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT6), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n373), .A2(new_n408), .A3(new_n375), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n378), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n410), .A2(new_n187), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT85), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT7), .B1(new_n405), .B2(G953), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n412), .B1(new_n404), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n403), .B1(new_n395), .B2(new_n396), .ZN(new_n415));
  AOI211_X1 g229(.A(KEYINPUT83), .B(new_n389), .C1(new_n392), .C2(new_n394), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n412), .B(new_n413), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  OR3_X1    g233(.A1(new_n415), .A2(new_n416), .A3(new_n413), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT84), .B1(new_n337), .B2(new_n351), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n336), .A2(G101), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n355), .B2(new_n356), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n344), .A2(new_n347), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n370), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT84), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n423), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n421), .A2(new_n427), .B1(new_n337), .B2(new_n351), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n374), .B(KEYINPUT8), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n420), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(KEYINPUT86), .B1(new_n419), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n413), .B1(new_n415), .B2(new_n416), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(KEYINPUT85), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n417), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n421), .A2(new_n427), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n352), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n429), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT86), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n435), .A2(new_n438), .A3(new_n439), .A4(new_n420), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n432), .A2(new_n440), .A3(new_n377), .ZN(new_n441));
  OAI21_X1  g255(.A(G210), .B1(G237), .B2(G902), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n411), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n442), .B(KEYINPUT87), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n445), .B1(new_n411), .B2(new_n441), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n443), .B1(new_n446), .B2(KEYINPUT88), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT88), .ZN(new_n448));
  AOI211_X1 g262(.A(new_n448), .B(new_n445), .C1(new_n411), .C2(new_n441), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n316), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT89), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT89), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n452), .B(new_n316), .C1(new_n447), .C2(new_n449), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n315), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT65), .B1(new_n271), .B2(G137), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT11), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT11), .ZN(new_n457));
  OAI211_X1 g271(.A(KEYINPUT65), .B(new_n457), .C1(new_n271), .C2(G137), .ZN(new_n458));
  INV_X1    g272(.A(G137), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n459), .A2(G134), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AND4_X1   g275(.A1(new_n212), .A2(new_n456), .A3(new_n458), .A4(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n460), .B1(new_n455), .B2(KEYINPUT11), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n212), .B1(new_n463), .B2(new_n458), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n394), .B(new_n392), .C1(new_n462), .C2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n463), .A2(new_n212), .A3(new_n458), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n271), .A2(G137), .ZN(new_n467));
  OAI21_X1  g281(.A(G131), .B1(new_n467), .B2(new_n460), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n268), .A2(G143), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n266), .A2(KEYINPUT64), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n204), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n398), .B1(new_n471), .B2(new_n380), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n393), .A2(new_n385), .A3(new_n401), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n466), .B(new_n468), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n465), .A2(KEYINPUT30), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(KEYINPUT30), .B1(new_n465), .B2(new_n474), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n475), .A2(new_n476), .A3(new_n372), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n465), .A2(new_n474), .A3(new_n371), .A4(new_n365), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n192), .A2(G210), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT27), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT26), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT27), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n192), .A2(new_n482), .A3(G210), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n481), .B1(new_n480), .B2(new_n483), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n322), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n480), .A2(new_n483), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT26), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n488), .A2(G101), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n478), .A2(new_n486), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(KEYINPUT31), .B1(new_n477), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n486), .A2(new_n490), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT28), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n465), .A2(new_n474), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n365), .A2(new_n371), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n494), .B1(new_n497), .B2(new_n478), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n478), .A2(new_n494), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n493), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n492), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n491), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT30), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n495), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n465), .A2(KEYINPUT30), .A3(new_n474), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(new_n496), .A3(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT69), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT31), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n503), .A2(new_n507), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n486), .A2(new_n490), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n507), .A2(new_n511), .A3(new_n509), .A4(new_n478), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT69), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n502), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(G472), .A2(G902), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT70), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT32), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n513), .A2(new_n510), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n492), .A2(new_n501), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT70), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n521), .A2(new_n522), .A3(new_n515), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n517), .A2(new_n518), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n497), .A2(new_n478), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT28), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n486), .A2(new_n490), .A3(KEYINPUT29), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n499), .A2(KEYINPUT71), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT71), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n529), .B1(new_n478), .B2(new_n494), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n526), .B(new_n527), .C1(new_n528), .C2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n187), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n511), .B1(new_n498), .B2(new_n500), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n507), .A2(new_n478), .A3(new_n493), .ZN(new_n534));
  AOI21_X1  g348(.A(KEYINPUT29), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(G472), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT72), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT72), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n538), .B(G472), .C1(new_n532), .C2(new_n535), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n516), .B1(new_n519), .B2(new_n520), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT32), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n524), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(G234), .ZN(new_n544));
  OAI21_X1  g358(.A(G217), .B1(new_n544), .B2(G902), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n272), .B(G119), .C1(KEYINPUT73), .C2(KEYINPUT23), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT23), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n547), .B1(new_n339), .B2(G128), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT73), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(new_n339), .B2(G128), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n546), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(G119), .B(G128), .ZN(new_n552));
  XOR2_X1   g366(.A(KEYINPUT24), .B(G110), .Z(new_n553));
  AOI22_X1  g367(.A1(new_n551), .A2(G110), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n226), .A2(new_n554), .ZN(new_n555));
  OAI22_X1  g369(.A1(new_n551), .A2(G110), .B1(new_n552), .B2(new_n553), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n556), .A2(new_n205), .A3(new_n225), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT75), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n555), .A2(new_n557), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT75), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n194), .A2(G221), .A3(G234), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(KEYINPUT22), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(G137), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n560), .A2(new_n562), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n558), .A2(new_n565), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n567), .A2(new_n187), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n545), .B1(new_n569), .B2(KEYINPUT25), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n570), .B1(KEYINPUT25), .B2(new_n569), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n567), .A2(new_n568), .ZN(new_n572));
  AOI21_X1  g386(.A(G902), .B1(new_n544), .B2(G217), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n543), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n329), .A2(new_n332), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n358), .B1(new_n578), .B2(KEYINPUT4), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n388), .B1(new_n579), .B2(new_n354), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n471), .A2(KEYINPUT1), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n387), .B1(new_n581), .B2(G128), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n337), .B1(new_n473), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT10), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n462), .A2(new_n464), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n472), .A2(new_n473), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n587), .A2(new_n584), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n337), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n580), .A2(new_n585), .A3(new_n586), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n400), .A2(new_n402), .ZN(new_n591));
  OAI21_X1  g405(.A(KEYINPUT80), .B1(new_n337), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT80), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n423), .A2(new_n587), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n592), .A2(new_n594), .A3(new_n583), .ZN(new_n595));
  INV_X1    g409(.A(new_n586), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT81), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(KEYINPUT12), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n601), .B1(new_n595), .B2(new_n596), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n590), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(G110), .B(G140), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n194), .A2(G227), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n590), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n585), .A2(new_n589), .ZN(new_n609));
  INV_X1    g423(.A(new_n388), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n360), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n596), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g426(.A1(new_n603), .A2(new_n606), .B1(new_n608), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(G469), .B1(new_n613), .B2(G902), .ZN(new_n614));
  INV_X1    g428(.A(G469), .ZN(new_n615));
  INV_X1    g429(.A(new_n601), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n597), .A2(new_n616), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n595), .B(new_n596), .C1(new_n598), .C2(KEYINPUT12), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n619), .A2(new_n608), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n607), .B1(new_n612), .B2(new_n590), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n615), .B(new_n187), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n614), .A2(KEYINPUT82), .A3(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(G221), .B1(new_n295), .B2(G902), .ZN(new_n624));
  XOR2_X1   g438(.A(new_n624), .B(KEYINPUT76), .Z(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT82), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n627), .B(G469), .C1(new_n613), .C2(G902), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n623), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n577), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n454), .A2(new_n630), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n323), .A2(new_n325), .ZN(new_n632));
  XOR2_X1   g446(.A(new_n631), .B(new_n632), .Z(G3));
  AND4_X1   g447(.A1(new_n187), .A2(new_n441), .A3(new_n410), .A4(new_n442), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n442), .B1(new_n411), .B2(new_n441), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n316), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT98), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI211_X1 g452(.A(KEYINPUT98), .B(new_n316), .C1(new_n634), .C2(new_n635), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n638), .A2(new_n314), .A3(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(G472), .B1(new_n514), .B2(G902), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT97), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(G472), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n521), .B2(new_n187), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(KEYINPUT97), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n643), .A2(new_n646), .A3(new_n517), .A4(new_n523), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n647), .A2(new_n629), .A3(new_n575), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT33), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n301), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n299), .A2(KEYINPUT33), .A3(new_n300), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n650), .A2(G478), .A3(new_n187), .A4(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n302), .A2(new_n303), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n652), .A2(KEYINPUT99), .A3(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(KEYINPUT99), .B1(new_n652), .B2(new_n653), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n657), .A2(new_n254), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n640), .A2(new_n648), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT34), .B(G104), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G6));
  INV_X1    g475(.A(KEYINPUT101), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n238), .B(new_n662), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n248), .A2(new_n250), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n664), .A2(KEYINPUT100), .A3(new_n251), .ZN(new_n665));
  OR3_X1    g479(.A1(new_n248), .A2(KEYINPUT100), .A3(new_n250), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n665), .A2(new_n307), .A3(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n638), .A2(new_n314), .A3(new_n639), .A4(new_n668), .ZN(new_n669));
  AND2_X1   g483(.A1(new_n669), .A2(KEYINPUT102), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n669), .A2(KEYINPUT102), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n648), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT35), .B(G107), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT103), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n672), .B(new_n674), .ZN(G9));
  NAND2_X1  g489(.A1(new_n560), .A2(new_n562), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n566), .A2(KEYINPUT36), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n676), .B(new_n677), .Z(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n573), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n571), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n647), .A2(new_n629), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n454), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT37), .B(G110), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G12));
  NAND2_X1  g499(.A1(new_n638), .A2(new_n639), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n686), .A2(new_n629), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n543), .A2(new_n680), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(G900), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n311), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n310), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n668), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n687), .A2(new_n689), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G128), .ZN(G30));
  AND3_X1   g511(.A1(new_n623), .A2(new_n626), .A3(new_n628), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n693), .B(KEYINPUT39), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n700), .B(KEYINPUT40), .Z(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT106), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n254), .A2(new_n307), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n316), .A3(new_n681), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT105), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n493), .B1(new_n507), .B2(new_n478), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n187), .B1(new_n511), .B2(new_n525), .ZN(new_n707));
  OAI21_X1  g521(.A(G472), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n524), .A2(new_n542), .A3(new_n708), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n702), .A2(new_n705), .A3(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n447), .A2(new_n449), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT104), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT38), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n710), .B(new_n713), .C1(KEYINPUT106), .C2(new_n701), .ZN(new_n714));
  XOR2_X1   g528(.A(new_n714), .B(new_n198), .Z(G45));
  OAI211_X1 g529(.A(new_n254), .B(new_n693), .C1(new_n656), .C2(new_n655), .ZN(new_n716));
  NOR4_X1   g530(.A1(new_n686), .A2(new_n688), .A3(new_n629), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(new_n204), .ZN(G48));
  NAND2_X1  g532(.A1(new_n612), .A2(new_n590), .ZN(new_n719));
  AOI22_X1  g533(.A1(new_n619), .A2(new_n608), .B1(new_n719), .B2(new_n606), .ZN(new_n720));
  OAI21_X1  g534(.A(G469), .B1(new_n720), .B2(G902), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n622), .A3(new_n722), .ZN(new_n723));
  OAI211_X1 g537(.A(KEYINPUT107), .B(G469), .C1(new_n720), .C2(G902), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n625), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n543), .A2(new_n576), .A3(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT108), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n640), .A2(new_n726), .A3(new_n727), .A4(new_n658), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n638), .A2(new_n658), .A3(new_n639), .A4(new_n314), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n543), .A2(new_n725), .A3(new_n576), .ZN(new_n730));
  OAI21_X1  g544(.A(KEYINPUT108), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(KEYINPUT41), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G113), .ZN(G15));
  OAI21_X1  g548(.A(new_n726), .B1(new_n670), .B2(new_n671), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(KEYINPUT109), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n737), .B(new_n726), .C1(new_n670), .C2(new_n671), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  XOR2_X1   g553(.A(new_n739), .B(KEYINPUT110), .Z(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G116), .ZN(G18));
  INV_X1    g555(.A(new_n725), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n686), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n688), .A2(new_n315), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G119), .ZN(G21));
  AND3_X1   g560(.A1(new_n638), .A2(new_n639), .A3(new_n703), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n526), .B1(new_n528), .B2(new_n530), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n526), .B(KEYINPUT111), .C1(new_n528), .C2(new_n530), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(new_n493), .A3(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n519), .A3(new_n492), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n515), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n576), .A2(new_n754), .A3(new_n314), .A4(new_n641), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n742), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n747), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G122), .ZN(G24));
  INV_X1    g572(.A(new_n686), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n754), .A2(new_n680), .A3(new_n641), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n716), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n759), .A2(new_n725), .A3(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G125), .ZN(G27));
  INV_X1    g577(.A(new_n447), .ZN(new_n764));
  INV_X1    g578(.A(new_n449), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n614), .A2(new_n622), .ZN(new_n766));
  INV_X1    g580(.A(new_n316), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n625), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n764), .A2(new_n765), .A3(new_n766), .A4(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT42), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n716), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n541), .A2(KEYINPUT32), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT112), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n775), .B1(new_n541), .B2(KEYINPUT32), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n774), .B(new_n540), .C1(new_n773), .C2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT113), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n777), .A2(new_n778), .A3(new_n576), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n778), .B1(new_n777), .B2(new_n576), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n772), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n768), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n447), .A2(new_n449), .A3(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n783), .A2(new_n543), .A3(new_n576), .A4(new_n766), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n770), .B1(new_n784), .B2(new_n716), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G131), .ZN(G33));
  NOR3_X1   g601(.A1(new_n769), .A2(new_n577), .A3(new_n694), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(new_n271), .ZN(G36));
  NOR2_X1   g603(.A1(new_n655), .A2(new_n656), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n790), .A2(new_n254), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT43), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(new_n647), .A3(new_n680), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT44), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n613), .A2(KEYINPUT45), .ZN(new_n796));
  OAI21_X1  g610(.A(G469), .B1(new_n613), .B2(KEYINPUT45), .ZN(new_n797));
  OAI22_X1  g611(.A1(new_n796), .A2(new_n797), .B1(new_n615), .B2(new_n187), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT46), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n622), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n801), .B1(new_n798), .B2(new_n799), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n625), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n803), .A2(new_n699), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n795), .A2(new_n804), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n793), .A2(new_n794), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n447), .A2(new_n767), .A3(new_n449), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n806), .A2(KEYINPUT114), .A3(new_n807), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n805), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(new_n459), .ZN(G39));
  XNOR2_X1  g627(.A(new_n803), .B(KEYINPUT47), .ZN(new_n814));
  INV_X1    g628(.A(new_n807), .ZN(new_n815));
  NOR4_X1   g629(.A1(new_n815), .A2(new_n543), .A3(new_n576), .A4(new_n716), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n814), .A2(KEYINPUT115), .A3(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT115), .B1(new_n814), .B2(new_n816), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(new_n218), .ZN(G42));
  NOR2_X1   g635(.A1(G952), .A2(G953), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(KEYINPUT122), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n792), .A2(new_n310), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n825), .A2(new_n576), .A3(new_n641), .A4(new_n754), .ZN(new_n826));
  OR4_X1    g640(.A1(new_n316), .A2(new_n713), .A3(new_n826), .A4(new_n742), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT120), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT50), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n827), .A2(KEYINPUT120), .A3(KEYINPUT50), .ZN(new_n831));
  INV_X1    g645(.A(new_n826), .ZN(new_n832));
  INV_X1    g646(.A(new_n723), .ZN(new_n833));
  INV_X1    g647(.A(new_n724), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n835), .A2(new_n626), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n832), .B(new_n807), .C1(new_n814), .C2(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n783), .B1(new_n834), .B2(new_n833), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n824), .A2(new_n760), .A3(new_n838), .ZN(new_n839));
  NOR4_X1   g653(.A1(new_n838), .A2(new_n692), .A3(new_n575), .A4(new_n709), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n657), .A2(new_n254), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n830), .A2(new_n831), .A3(new_n837), .A4(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT51), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n843), .A2(new_n844), .ZN(new_n846));
  AOI211_X1 g660(.A(new_n309), .B(G953), .C1(new_n840), .C2(new_n658), .ZN(new_n847));
  INV_X1    g661(.A(new_n743), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n847), .B1(new_n848), .B2(new_n826), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n849), .A2(KEYINPUT121), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n849), .A2(KEYINPUT121), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n779), .A2(new_n780), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n852), .A2(new_n824), .A3(new_n838), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(KEYINPUT48), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n850), .A2(new_n851), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n845), .A2(new_n846), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n451), .A2(new_n453), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n308), .B1(new_n254), .B2(new_n790), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n858), .A2(new_n314), .A3(new_n648), .A4(new_n859), .ZN(new_n860));
  AOI22_X1  g674(.A1(new_n743), .A2(new_n744), .B1(new_n747), .B2(new_n756), .ZN(new_n861));
  INV_X1    g675(.A(new_n315), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n858), .B(new_n862), .C1(new_n630), .C2(new_n682), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n732), .A2(new_n860), .A3(new_n861), .A4(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n864), .B1(new_n738), .B2(new_n736), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n761), .A2(new_n783), .A3(new_n766), .ZN(new_n866));
  INV_X1    g680(.A(new_n307), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n867), .A2(new_n666), .A3(new_n665), .A4(new_n693), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(new_n663), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n807), .A2(new_n698), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n866), .B1(new_n870), .B2(new_n688), .ZN(new_n871));
  AOI211_X1 g685(.A(new_n788), .B(new_n871), .C1(new_n785), .C2(new_n781), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT118), .B1(new_n865), .B2(new_n872), .ZN(new_n873));
  AND4_X1   g687(.A1(new_n732), .A2(new_n860), .A3(new_n861), .A4(new_n863), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n739), .A2(new_n874), .A3(KEYINPUT118), .A4(new_n872), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n687), .A2(new_n658), .A3(new_n689), .A4(new_n693), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n696), .A2(new_n876), .A3(new_n762), .ZN(new_n877));
  AND4_X1   g691(.A1(new_n766), .A2(new_n681), .A3(new_n626), .A4(new_n693), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n747), .A2(new_n709), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n877), .A2(KEYINPUT52), .A3(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT52), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n876), .A2(new_n696), .A3(new_n762), .ZN(new_n882));
  INV_X1    g696(.A(new_n879), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n875), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n857), .B1(new_n873), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n739), .A2(new_n874), .A3(new_n872), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT118), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n890), .A2(KEYINPUT53), .A3(new_n885), .A4(new_n875), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n887), .A2(KEYINPUT119), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT119), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n893), .B(new_n857), .C1(new_n873), .C2(new_n886), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n892), .A2(KEYINPUT54), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n885), .A2(KEYINPUT53), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n896), .A2(new_n888), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT54), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n887), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n823), .B1(new_n856), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n835), .A2(KEYINPUT49), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n902), .A2(new_n576), .A3(new_n768), .A4(new_n791), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT116), .Z(new_n904));
  NOR2_X1   g718(.A1(new_n835), .A2(KEYINPUT49), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT117), .ZN(new_n906));
  OR3_X1    g720(.A1(new_n713), .A2(new_n709), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n901), .B1(new_n904), .B2(new_n907), .ZN(G75));
  NOR2_X1   g722(.A1(new_n194), .A2(G952), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n378), .A2(new_n409), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT123), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n407), .B(KEYINPUT55), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n911), .B(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n887), .A2(new_n897), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n914), .A2(G210), .A3(G902), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT56), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n913), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n914), .A2(G902), .A3(new_n444), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n913), .A2(new_n916), .ZN(new_n919));
  AOI211_X1 g733(.A(new_n909), .B(new_n917), .C1(new_n918), .C2(new_n919), .ZN(G51));
  NAND2_X1  g734(.A1(new_n914), .A2(KEYINPUT54), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n899), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n615), .A2(new_n187), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT57), .Z(new_n925));
  OAI22_X1  g739(.A1(new_n923), .A2(new_n925), .B1(new_n621), .B2(new_n620), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n914), .A2(G902), .ZN(new_n927));
  OR3_X1    g741(.A1(new_n927), .A2(new_n796), .A3(new_n797), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n909), .B1(new_n926), .B2(new_n928), .ZN(G54));
  NAND4_X1  g743(.A1(new_n914), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n229), .A2(new_n245), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n930), .A2(new_n931), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n932), .A2(new_n933), .A3(new_n909), .ZN(G60));
  INV_X1    g748(.A(KEYINPUT124), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n650), .A2(new_n651), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(G478), .A2(G902), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT59), .Z(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n937), .B1(new_n900), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n936), .A2(new_n939), .ZN(new_n942));
  INV_X1    g756(.A(new_n899), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n898), .B1(new_n887), .B2(new_n897), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n909), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n935), .B1(new_n941), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n909), .B1(new_n922), .B2(new_n942), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n939), .B1(new_n895), .B2(new_n899), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n949), .B(KEYINPUT124), .C1(new_n950), .C2(new_n937), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n948), .A2(new_n951), .ZN(G63));
  NAND2_X1  g766(.A1(G217), .A2(G902), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT60), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n954), .B1(new_n887), .B2(new_n897), .ZN(new_n955));
  OR2_X1    g769(.A1(new_n955), .A2(new_n572), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n678), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n956), .A2(new_n946), .A3(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT61), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(G66));
  NOR3_X1   g774(.A1(new_n312), .A2(new_n405), .A3(new_n194), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n961), .B1(new_n865), .B2(new_n194), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n911), .B1(G898), .B2(new_n194), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(G69));
  AOI21_X1  g778(.A(new_n194), .B1(G227), .B2(G900), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n475), .A2(new_n476), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n242), .B(KEYINPUT125), .Z(new_n967));
  XOR2_X1   g781(.A(new_n966), .B(new_n967), .Z(new_n968));
  INV_X1    g782(.A(new_n811), .ZN(new_n969));
  AOI21_X1  g783(.A(KEYINPUT114), .B1(new_n806), .B2(new_n807), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI211_X1 g785(.A(KEYINPUT126), .B(new_n877), .C1(new_n971), .C2(new_n805), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT126), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n973), .B1(new_n812), .B2(new_n882), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n804), .B(new_n747), .C1(new_n779), .C2(new_n780), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n788), .B1(new_n781), .B2(new_n785), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n820), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n975), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n194), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT127), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n194), .A2(G900), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n981), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(G953), .B1(new_n975), .B2(new_n979), .ZN(new_n986));
  OAI21_X1  g800(.A(KEYINPUT127), .B1(new_n986), .B2(new_n983), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n968), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n968), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n714), .A2(new_n877), .ZN(new_n990));
  OR2_X1    g804(.A1(new_n990), .A2(KEYINPUT62), .ZN(new_n991));
  INV_X1    g805(.A(new_n859), .ZN(new_n992));
  NOR4_X1   g806(.A1(new_n700), .A2(new_n815), .A3(new_n992), .A4(new_n577), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n812), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n820), .B1(new_n990), .B2(KEYINPUT62), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n991), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n989), .B1(new_n996), .B2(new_n194), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n965), .B1(new_n988), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n982), .B1(new_n981), .B2(new_n984), .ZN(new_n999));
  NOR3_X1   g813(.A1(new_n986), .A2(KEYINPUT127), .A3(new_n983), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n989), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n965), .ZN(new_n1002));
  INV_X1    g816(.A(new_n997), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n998), .A2(new_n1004), .ZN(G72));
  INV_X1    g819(.A(new_n706), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n991), .A2(new_n995), .A3(new_n865), .A4(new_n994), .ZN(new_n1007));
  NAND2_X1  g821(.A1(G472), .A2(G902), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT63), .Z(new_n1009));
  AOI21_X1  g823(.A(new_n1006), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  AND3_X1   g824(.A1(new_n1006), .A2(new_n534), .A3(new_n1009), .ZN(new_n1011));
  AND3_X1   g825(.A1(new_n892), .A2(new_n894), .A3(new_n1011), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n975), .A2(new_n865), .A3(new_n979), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n534), .B1(new_n1013), .B2(new_n1009), .ZN(new_n1014));
  NOR4_X1   g828(.A1(new_n1010), .A2(new_n1012), .A3(new_n1014), .A4(new_n909), .ZN(G57));
endmodule


