

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n735, n736, n737,
         n738, n739, n740, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790;

  INV_X1 U374 ( .A(n742), .ZN(n353) );
  OR2_X1 U375 ( .A1(G237), .A2(G902), .ZN(n526) );
  XNOR2_X1 U376 ( .A(G101), .B(G107), .ZN(n562) );
  XNOR2_X1 U377 ( .A(n352), .B(KEYINPUT116), .ZN(n735) );
  BUF_X1 U378 ( .A(G143), .Z(n412) );
  BUF_X1 U379 ( .A(n740), .Z(n366) );
  NAND2_X1 U380 ( .A1(n351), .A2(n437), .ZN(n439) );
  NAND2_X1 U381 ( .A1(n665), .A2(KEYINPUT120), .ZN(n351) );
  NAND2_X1 U382 ( .A1(n732), .A2(n733), .ZN(n352) );
  NAND2_X2 U383 ( .A1(n386), .A2(n453), .ZN(n399) );
  AND2_X2 U384 ( .A1(n399), .A2(n377), .ZN(n407) );
  XNOR2_X2 U385 ( .A(n400), .B(n434), .ZN(n411) );
  XNOR2_X2 U386 ( .A(n354), .B(n353), .ZN(n743) );
  NAND2_X1 U387 ( .A1(n740), .A2(G210), .ZN(n354) );
  XNOR2_X1 U388 ( .A(G134), .B(G122), .ZN(n491) );
  BUF_X1 U389 ( .A(G113), .Z(n693) );
  XOR2_X1 U390 ( .A(n560), .B(KEYINPUT21), .Z(n355) );
  AND2_X2 U391 ( .A1(n459), .A2(n458), .ZN(n475) );
  INV_X2 U392 ( .A(n512), .ZN(n514) );
  XNOR2_X2 U393 ( .A(G101), .B(G113), .ZN(n512) );
  INV_X4 U394 ( .A(G116), .ZN(n406) );
  XNOR2_X1 U395 ( .A(n767), .B(n519), .ZN(n523) );
  AND2_X1 U396 ( .A1(n666), .A2(G217), .ZN(n357) );
  INV_X1 U397 ( .A(KEYINPUT76), .ZN(n358) );
  INV_X1 U398 ( .A(KEYINPUT22), .ZN(n575) );
  AND2_X1 U399 ( .A1(n599), .A2(n463), .ZN(n458) );
  XNOR2_X1 U400 ( .A(n613), .B(KEYINPUT40), .ZN(n788) );
  NOR2_X1 U401 ( .A1(n691), .A2(n650), .ZN(n613) );
  AND2_X1 U402 ( .A1(n472), .A2(n469), .ZN(n468) );
  XNOR2_X1 U403 ( .A(n625), .B(n624), .ZN(n787) );
  NOR2_X1 U404 ( .A1(n593), .A2(n415), .ZN(n473) );
  XNOR2_X1 U405 ( .A(n576), .B(n575), .ZN(n593) );
  NAND2_X1 U406 ( .A1(n606), .A2(n489), .ZN(n359) );
  XNOR2_X1 U407 ( .A(n490), .B(KEYINPUT95), .ZN(n606) );
  AND2_X1 U408 ( .A1(n718), .A2(n355), .ZN(n416) );
  XNOR2_X1 U409 ( .A(n558), .B(n356), .ZN(n704) );
  XNOR2_X1 U410 ( .A(n523), .B(n522), .ZN(n737) );
  NOR2_X1 U411 ( .A1(n667), .A2(G902), .ZN(n356) );
  XNOR2_X1 U412 ( .A(n449), .B(n775), .ZN(n667) );
  XNOR2_X1 U413 ( .A(n750), .B(n749), .ZN(n751) );
  XNOR2_X1 U414 ( .A(n487), .B(n552), .ZN(n449) );
  XNOR2_X1 U415 ( .A(KEYINPUT20), .B(n554), .ZN(n559) );
  XNOR2_X1 U416 ( .A(n448), .B(n569), .ZN(n775) );
  XNOR2_X1 U417 ( .A(n550), .B(KEYINPUT82), .ZN(n488) );
  XNOR2_X1 U418 ( .A(n600), .B(KEYINPUT45), .ZN(n601) );
  XNOR2_X1 U419 ( .A(n546), .B(KEYINPUT10), .ZN(n448) );
  INV_X1 U420 ( .A(n553), .ZN(n664) );
  XNOR2_X1 U421 ( .A(G110), .B(KEYINPUT24), .ZN(n547) );
  XOR2_X2 U422 ( .A(KEYINPUT78), .B(G104), .Z(n563) );
  XNOR2_X1 U423 ( .A(G119), .B(G128), .ZN(n550) );
  XOR2_X1 U424 ( .A(KEYINPUT73), .B(G110), .Z(n568) );
  XOR2_X1 U425 ( .A(G902), .B(KEYINPUT15), .Z(n553) );
  OR2_X2 U426 ( .A1(n409), .A2(n408), .ZN(n395) );
  NAND2_X1 U427 ( .A1(n740), .A2(n357), .ZN(n437) );
  XNOR2_X1 U428 ( .A(n359), .B(n358), .ZN(n609) );
  XNOR2_X1 U429 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U430 ( .A(n549), .B(n488), .ZN(n487) );
  NAND2_X1 U431 ( .A1(n360), .A2(n433), .ZN(n432) );
  NAND2_X1 U432 ( .A1(n370), .A2(n369), .ZN(n360) );
  NOR2_X2 U433 ( .A1(n753), .A2(n760), .ZN(n754) );
  XOR2_X2 U434 ( .A(G122), .B(G104), .Z(n511) );
  XNOR2_X2 U435 ( .A(n776), .B(G146), .ZN(n571) );
  XNOR2_X2 U436 ( .A(n361), .B(n544), .ZN(n776) );
  NAND2_X1 U437 ( .A1(n363), .A2(n362), .ZN(n361) );
  NAND2_X1 U438 ( .A1(n542), .A2(G134), .ZN(n362) );
  NAND2_X1 U439 ( .A1(n388), .A2(n389), .ZN(n363) );
  BUF_X1 U440 ( .A(n538), .Z(n364) );
  BUF_X1 U441 ( .A(n767), .Z(n365) );
  OR2_X1 U442 ( .A1(n593), .A2(n466), .ZN(n465) );
  NOR2_X2 U443 ( .A1(n735), .A2(G953), .ZN(n736) );
  NAND2_X1 U444 ( .A1(n476), .A2(n601), .ZN(n369) );
  NAND2_X1 U445 ( .A1(n367), .A2(n368), .ZN(n370) );
  INV_X1 U446 ( .A(n476), .ZN(n367) );
  INV_X1 U447 ( .A(n601), .ZN(n368) );
  BUF_X1 U448 ( .A(n776), .Z(n371) );
  XNOR2_X1 U449 ( .A(n476), .B(n601), .ZN(n372) );
  NAND2_X1 U450 ( .A1(n379), .A2(n430), .ZN(n429) );
  AND2_X1 U451 ( .A1(n461), .A2(KEYINPUT85), .ZN(n460) );
  NOR2_X1 U452 ( .A1(G953), .A2(G237), .ZN(n539) );
  INV_X1 U453 ( .A(KEYINPUT33), .ZN(n434) );
  XNOR2_X1 U454 ( .A(n481), .B(KEYINPUT96), .ZN(n480) );
  INV_X1 U455 ( .A(G472), .ZN(n481) );
  XNOR2_X1 U456 ( .A(n418), .B(n543), .ZN(n503) );
  XNOR2_X1 U457 ( .A(n546), .B(KEYINPUT10), .ZN(n418) );
  NAND2_X1 U458 ( .A1(n424), .A2(n660), .ZN(n423) );
  INV_X1 U459 ( .A(n658), .ZN(n424) );
  NOR2_X1 U460 ( .A1(n415), .A2(KEYINPUT32), .ZN(n467) );
  NAND2_X1 U461 ( .A1(n470), .A2(KEYINPUT32), .ZN(n469) );
  NAND2_X1 U462 ( .A1(n594), .A2(n471), .ZN(n470) );
  INV_X1 U463 ( .A(n415), .ZN(n471) );
  BUF_X1 U464 ( .A(n704), .Z(n415) );
  XNOR2_X1 U465 ( .A(n570), .B(n404), .ZN(n403) );
  NOR2_X1 U466 ( .A1(G952), .A2(n782), .ZN(n760) );
  INV_X1 U467 ( .A(n787), .ZN(n447) );
  INV_X1 U468 ( .A(KEYINPUT46), .ZN(n446) );
  AND2_X1 U469 ( .A1(n464), .A2(KEYINPUT44), .ZN(n462) );
  INV_X1 U470 ( .A(G134), .ZN(n389) );
  INV_X1 U471 ( .A(n688), .ZN(n484) );
  NAND2_X1 U472 ( .A1(n787), .A2(KEYINPUT46), .ZN(n444) );
  XOR2_X1 U473 ( .A(KEYINPUT25), .B(KEYINPUT77), .Z(n556) );
  XNOR2_X1 U474 ( .A(G116), .B(G137), .ZN(n535) );
  XOR2_X1 U475 ( .A(KEYINPUT74), .B(KEYINPUT5), .Z(n536) );
  XOR2_X1 U476 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n517) );
  NOR2_X1 U477 ( .A1(n664), .A2(n486), .ZN(n485) );
  NAND2_X1 U478 ( .A1(G234), .A2(G237), .ZN(n529) );
  INV_X1 U479 ( .A(n614), .ZN(n489) );
  NAND2_X1 U480 ( .A1(n704), .A2(n355), .ZN(n561) );
  NAND2_X1 U481 ( .A1(n402), .A2(n410), .ZN(n409) );
  NAND2_X1 U482 ( .A1(n373), .A2(G902), .ZN(n410) );
  INV_X1 U483 ( .A(KEYINPUT92), .ZN(n564) );
  XNOR2_X1 U484 ( .A(n622), .B(n621), .ZN(n729) );
  XNOR2_X1 U485 ( .A(n612), .B(n611), .ZN(n650) );
  NOR2_X1 U486 ( .A1(n627), .A2(n717), .ZN(n612) );
  INV_X1 U487 ( .A(KEYINPUT6), .ZN(n401) );
  XNOR2_X1 U488 ( .A(n506), .B(n419), .ZN(n750) );
  XNOR2_X1 U489 ( .A(n374), .B(n507), .ZN(n419) );
  NAND2_X1 U490 ( .A1(n426), .A2(n425), .ZN(n663) );
  NAND2_X1 U491 ( .A1(n468), .A2(n465), .ZN(n790) );
  NAND2_X1 U492 ( .A1(n594), .A2(n467), .ZN(n466) );
  INV_X1 U493 ( .A(n760), .ZN(n451) );
  XNOR2_X1 U494 ( .A(n745), .B(n414), .ZN(n748) );
  XOR2_X1 U495 ( .A(n572), .B(G469), .Z(n373) );
  XOR2_X1 U496 ( .A(n505), .B(n504), .Z(n374) );
  NOR2_X1 U497 ( .A1(n659), .A2(n423), .ZN(n375) );
  XOR2_X1 U498 ( .A(n525), .B(n524), .Z(n376) );
  OR2_X1 U499 ( .A1(n605), .A2(n534), .ZN(n377) );
  AND2_X1 U500 ( .A1(n447), .A2(n446), .ZN(n378) );
  XNOR2_X1 U501 ( .A(n616), .B(n401), .ZN(n577) );
  INV_X1 U502 ( .A(n577), .ZN(n397) );
  AND2_X1 U503 ( .A1(n375), .A2(n485), .ZN(n379) );
  NOR2_X1 U504 ( .A1(n393), .A2(n724), .ZN(n380) );
  OR2_X1 U505 ( .A1(n373), .A2(G902), .ZN(n381) );
  XOR2_X1 U506 ( .A(KEYINPUT66), .B(KEYINPUT0), .Z(n382) );
  XOR2_X1 U507 ( .A(KEYINPUT48), .B(KEYINPUT70), .Z(n383) );
  INV_X1 U508 ( .A(n660), .ZN(n433) );
  BUF_X1 U509 ( .A(n520), .Z(n384) );
  INV_X1 U510 ( .A(n610), .ZN(n385) );
  NOR2_X1 U511 ( .A1(n593), .A2(n397), .ZN(n578) );
  INV_X1 U512 ( .A(n655), .ZN(n386) );
  INV_X1 U513 ( .A(n655), .ZN(n610) );
  NOR2_X2 U514 ( .A1(n456), .A2(n455), .ZN(n454) );
  NAND2_X1 U515 ( .A1(n574), .A2(n702), .ZN(n387) );
  INV_X1 U516 ( .A(n542), .ZN(n388) );
  NAND2_X1 U517 ( .A1(n574), .A2(n702), .ZN(n580) );
  XNOR2_X1 U518 ( .A(n395), .B(KEYINPUT1), .ZN(n390) );
  BUF_X1 U519 ( .A(n428), .Z(n391) );
  NAND2_X1 U520 ( .A1(n432), .A2(n431), .ZN(n428) );
  XNOR2_X1 U521 ( .A(n477), .B(KEYINPUT35), .ZN(n392) );
  BUF_X1 U522 ( .A(n411), .Z(n393) );
  XNOR2_X1 U523 ( .A(n477), .B(KEYINPUT35), .ZN(n786) );
  XNOR2_X1 U524 ( .A(n580), .B(n435), .ZN(n398) );
  XNOR2_X2 U525 ( .A(n394), .B(n382), .ZN(n396) );
  NAND2_X1 U526 ( .A1(n407), .A2(n454), .ZN(n394) );
  NAND2_X1 U527 ( .A1(n702), .A2(n395), .ZN(n490) );
  XNOR2_X2 U528 ( .A(n395), .B(KEYINPUT1), .ZN(n574) );
  NAND2_X1 U529 ( .A1(n619), .A2(n395), .ZN(n620) );
  NAND2_X1 U530 ( .A1(n396), .A2(n712), .ZN(n581) );
  AND2_X1 U531 ( .A1(n396), .A2(n416), .ZN(n576) );
  XNOR2_X2 U532 ( .A(n396), .B(KEYINPUT91), .ZN(n582) );
  NAND2_X1 U533 ( .A1(n398), .A2(n397), .ZN(n400) );
  XNOR2_X2 U534 ( .A(n482), .B(n480), .ZN(n616) );
  NAND2_X1 U535 ( .A1(n454), .A2(n399), .ZN(n629) );
  NAND2_X1 U536 ( .A1(n747), .A2(n373), .ZN(n402) );
  XNOR2_X2 U537 ( .A(n571), .B(n403), .ZN(n747) );
  INV_X1 U538 ( .A(n569), .ZN(n404) );
  XNOR2_X2 U539 ( .A(n405), .B(n376), .ZN(n655) );
  OR2_X2 U540 ( .A1(n737), .A2(n553), .ZN(n405) );
  XNOR2_X2 U541 ( .A(n406), .B(G107), .ZN(n510) );
  NOR2_X1 U542 ( .A1(n747), .A2(n381), .ZN(n408) );
  NOR2_X2 U543 ( .A1(n411), .A2(n582), .ZN(n573) );
  NOR2_X1 U544 ( .A1(n393), .A2(n729), .ZN(n730) );
  NAND2_X1 U545 ( .A1(n740), .A2(G217), .ZN(n665) );
  INV_X1 U546 ( .A(n626), .ZN(n478) );
  NAND2_X2 U547 ( .A1(n427), .A2(n429), .ZN(n740) );
  XNOR2_X1 U548 ( .A(n413), .B(n566), .ZN(n570) );
  XNOR2_X1 U549 ( .A(n567), .B(n568), .ZN(n413) );
  NAND2_X1 U550 ( .A1(n428), .A2(n485), .ZN(n427) );
  INV_X2 U551 ( .A(G143), .ZN(n422) );
  XNOR2_X1 U552 ( .A(n747), .B(n746), .ZN(n414) );
  XOR2_X2 U553 ( .A(KEYINPUT68), .B(G131), .Z(n543) );
  XNOR2_X2 U554 ( .A(G119), .B(KEYINPUT3), .ZN(n513) );
  XNOR2_X1 U555 ( .A(n417), .B(n672), .ZN(G57) );
  NOR2_X2 U556 ( .A1(n671), .A2(n760), .ZN(n417) );
  OR2_X2 U557 ( .A1(n659), .A2(n658), .ZN(n780) );
  NAND2_X1 U558 ( .A1(n483), .A2(n444), .ZN(n443) );
  NAND2_X1 U559 ( .A1(n420), .A2(n460), .ZN(n459) );
  OR2_X1 U560 ( .A1(n420), .A2(KEYINPUT85), .ZN(n474) );
  XNOR2_X1 U561 ( .A(n592), .B(n591), .ZN(n420) );
  XNOR2_X2 U562 ( .A(n520), .B(n421), .ZN(n542) );
  XNOR2_X2 U563 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n421) );
  XNOR2_X2 U564 ( .A(n422), .B(G128), .ZN(n520) );
  NAND2_X1 U565 ( .A1(n430), .A2(n375), .ZN(n425) );
  INV_X1 U566 ( .A(n391), .ZN(n426) );
  INV_X1 U567 ( .A(n372), .ZN(n430) );
  NAND2_X1 U568 ( .A1(n780), .A2(n433), .ZN(n431) );
  INV_X1 U569 ( .A(KEYINPUT100), .ZN(n435) );
  NAND2_X1 U570 ( .A1(n438), .A2(n451), .ZN(n450) );
  XNOR2_X1 U571 ( .A(n439), .B(n452), .ZN(n438) );
  NAND2_X1 U572 ( .A1(n441), .A2(n440), .ZN(n445) );
  NAND2_X1 U573 ( .A1(n788), .A2(KEYINPUT46), .ZN(n440) );
  NAND2_X1 U574 ( .A1(n442), .A2(n378), .ZN(n441) );
  INV_X1 U575 ( .A(n788), .ZN(n442) );
  NOR2_X2 U576 ( .A1(n445), .A2(n443), .ZN(n649) );
  XNOR2_X1 U577 ( .A(n450), .B(KEYINPUT121), .ZN(G66) );
  INV_X1 U578 ( .A(n667), .ZN(n452) );
  NAND2_X1 U579 ( .A1(n610), .A2(n653), .ZN(n638) );
  NOR2_X1 U580 ( .A1(n716), .A2(n528), .ZN(n453) );
  NOR2_X1 U581 ( .A1(n653), .A2(KEYINPUT19), .ZN(n455) );
  AND2_X1 U582 ( .A1(n655), .A2(n528), .ZN(n456) );
  XNOR2_X2 U583 ( .A(n457), .B(n515), .ZN(n767) );
  XNOR2_X2 U584 ( .A(n538), .B(KEYINPUT16), .ZN(n457) );
  XNOR2_X2 U585 ( .A(n514), .B(n513), .ZN(n538) );
  NAND2_X1 U586 ( .A1(n596), .A2(KEYINPUT44), .ZN(n461) );
  NAND2_X1 U587 ( .A1(n596), .A2(n462), .ZN(n463) );
  INV_X1 U588 ( .A(KEYINPUT85), .ZN(n464) );
  NAND2_X1 U589 ( .A1(n593), .A2(KEYINPUT32), .ZN(n472) );
  NAND2_X2 U590 ( .A1(n475), .A2(n474), .ZN(n476) );
  NAND2_X1 U591 ( .A1(n786), .A2(KEYINPUT44), .ZN(n590) );
  NAND2_X1 U592 ( .A1(n479), .A2(n478), .ZN(n477) );
  XNOR2_X1 U593 ( .A(n573), .B(KEYINPUT34), .ZN(n479) );
  OR2_X2 U594 ( .A1(n668), .A2(G902), .ZN(n482) );
  XNOR2_X1 U595 ( .A(n571), .B(n545), .ZN(n668) );
  NOR2_X1 U596 ( .A1(n648), .A2(n484), .ZN(n483) );
  NAND2_X1 U597 ( .A1(n663), .A2(n662), .ZN(n732) );
  INV_X1 U598 ( .A(n662), .ZN(n486) );
  NOR2_X2 U599 ( .A1(n760), .A2(n743), .ZN(n744) );
  INV_X1 U600 ( .A(KEYINPUT86), .ZN(n591) );
  INV_X1 U601 ( .A(n633), .ZN(n647) );
  XNOR2_X1 U602 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U603 ( .A(n518), .B(KEYINPUT79), .ZN(n519) );
  INV_X1 U604 ( .A(n700), .ZN(n657) );
  XNOR2_X1 U605 ( .A(n521), .B(n568), .ZN(n522) );
  NAND2_X1 U606 ( .A1(n657), .A2(n701), .ZN(n658) );
  INV_X1 U607 ( .A(KEYINPUT80), .ZN(n524) );
  XNOR2_X1 U608 ( .A(n668), .B(KEYINPUT62), .ZN(n669) );
  XNOR2_X1 U609 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U610 ( .A(n752), .B(n751), .ZN(n753) );
  XNOR2_X1 U611 ( .A(KEYINPUT99), .B(G478), .ZN(n501) );
  XOR2_X1 U612 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n492) );
  XNOR2_X1 U613 ( .A(n492), .B(n491), .ZN(n496) );
  XOR2_X1 U614 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n494) );
  XNOR2_X1 U615 ( .A(n384), .B(n510), .ZN(n493) );
  XNOR2_X1 U616 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U617 ( .A(n496), .B(n495), .Z(n499) );
  INV_X2 U618 ( .A(G953), .ZN(n782) );
  NAND2_X1 U619 ( .A1(G234), .A2(n782), .ZN(n497) );
  XOR2_X1 U620 ( .A(KEYINPUT8), .B(n497), .Z(n551) );
  NAND2_X1 U621 ( .A1(G217), .A2(n551), .ZN(n498) );
  XNOR2_X1 U622 ( .A(n499), .B(n498), .ZN(n755) );
  NOR2_X1 U623 ( .A1(G902), .A2(n755), .ZN(n500) );
  XNOR2_X1 U624 ( .A(n501), .B(n500), .ZN(n586) );
  XNOR2_X1 U625 ( .A(KEYINPUT13), .B(G475), .ZN(n509) );
  XOR2_X2 U626 ( .A(G146), .B(G125), .Z(n546) );
  XNOR2_X1 U627 ( .A(n693), .B(n412), .ZN(n502) );
  XNOR2_X1 U628 ( .A(n503), .B(n502), .ZN(n506) );
  XOR2_X1 U629 ( .A(G140), .B(KEYINPUT12), .Z(n505) );
  NAND2_X1 U630 ( .A1(G214), .A2(n539), .ZN(n504) );
  XNOR2_X1 U631 ( .A(n511), .B(KEYINPUT11), .ZN(n507) );
  NOR2_X1 U632 ( .A1(G902), .A2(n750), .ZN(n508) );
  XNOR2_X1 U633 ( .A(n509), .B(n508), .ZN(n584) );
  NAND2_X1 U634 ( .A1(n586), .A2(n584), .ZN(n626) );
  XOR2_X1 U635 ( .A(n511), .B(n510), .Z(n515) );
  NAND2_X1 U636 ( .A1(G224), .A2(n782), .ZN(n516) );
  XNOR2_X1 U637 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U638 ( .A(n542), .B(n546), .Z(n521) );
  NAND2_X1 U639 ( .A1(G210), .A2(n526), .ZN(n525) );
  NAND2_X1 U640 ( .A1(G214), .A2(n526), .ZN(n527) );
  XOR2_X1 U641 ( .A(KEYINPUT88), .B(n527), .Z(n716) );
  INV_X1 U642 ( .A(n716), .ZN(n653) );
  INV_X1 U643 ( .A(KEYINPUT19), .ZN(n528) );
  XOR2_X1 U644 ( .A(KEYINPUT14), .B(KEYINPUT89), .Z(n530) );
  XNOR2_X1 U645 ( .A(n530), .B(n529), .ZN(n531) );
  NAND2_X1 U646 ( .A1(G952), .A2(n531), .ZN(n728) );
  NOR2_X1 U647 ( .A1(G953), .A2(n728), .ZN(n605) );
  AND2_X1 U648 ( .A1(G953), .A2(n531), .ZN(n532) );
  NAND2_X1 U649 ( .A1(G902), .A2(n532), .ZN(n602) );
  NOR2_X1 U650 ( .A1(G898), .A2(n602), .ZN(n533) );
  XNOR2_X1 U651 ( .A(n533), .B(KEYINPUT90), .ZN(n534) );
  XNOR2_X1 U652 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U653 ( .A(n364), .B(n537), .Z(n541) );
  NAND2_X1 U654 ( .A1(n539), .A2(G210), .ZN(n540) );
  XNOR2_X1 U655 ( .A(n541), .B(n540), .ZN(n545) );
  XOR2_X1 U656 ( .A(KEYINPUT69), .B(n543), .Z(n544) );
  XOR2_X1 U657 ( .A(G137), .B(G140), .Z(n569) );
  XOR2_X1 U658 ( .A(KEYINPUT23), .B(KEYINPUT93), .Z(n548) );
  NAND2_X1 U659 ( .A1(G221), .A2(n551), .ZN(n552) );
  NAND2_X1 U660 ( .A1(G234), .A2(n664), .ZN(n554) );
  NAND2_X1 U661 ( .A1(G217), .A2(n559), .ZN(n555) );
  XNOR2_X1 U662 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U663 ( .A(KEYINPUT94), .B(n557), .ZN(n558) );
  NAND2_X1 U664 ( .A1(n559), .A2(G221), .ZN(n560) );
  XNOR2_X2 U665 ( .A(n561), .B(KEYINPUT67), .ZN(n702) );
  XNOR2_X1 U666 ( .A(n563), .B(n562), .ZN(n567) );
  NAND2_X1 U667 ( .A1(G227), .A2(n782), .ZN(n565) );
  XNOR2_X1 U668 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n572) );
  NOR2_X1 U669 ( .A1(n586), .A2(n584), .ZN(n718) );
  NAND2_X1 U670 ( .A1(n415), .A2(n578), .ZN(n579) );
  NOR2_X1 U671 ( .A1(n390), .A2(n579), .ZN(n673) );
  NOR2_X1 U672 ( .A1(n616), .A2(n387), .ZN(n712) );
  XOR2_X1 U673 ( .A(KEYINPUT31), .B(n581), .Z(n694) );
  INV_X1 U674 ( .A(n616), .ZN(n710) );
  NOR2_X1 U675 ( .A1(n710), .A2(n582), .ZN(n583) );
  NAND2_X1 U676 ( .A1(n606), .A2(n583), .ZN(n675) );
  NAND2_X1 U677 ( .A1(n694), .A2(n675), .ZN(n587) );
  INV_X1 U678 ( .A(n584), .ZN(n585) );
  OR2_X1 U679 ( .A1(n585), .A2(n586), .ZN(n691) );
  NAND2_X1 U680 ( .A1(n586), .A2(n585), .ZN(n695) );
  NAND2_X1 U681 ( .A1(n691), .A2(n695), .ZN(n721) );
  AND2_X1 U682 ( .A1(n587), .A2(n721), .ZN(n588) );
  NOR2_X1 U683 ( .A1(n673), .A2(n588), .ZN(n589) );
  NAND2_X1 U684 ( .A1(n590), .A2(n589), .ZN(n592) );
  XNOR2_X1 U685 ( .A(KEYINPUT87), .B(n390), .ZN(n643) );
  NOR2_X1 U686 ( .A1(n643), .A2(n397), .ZN(n594) );
  NOR2_X1 U687 ( .A1(n390), .A2(n710), .ZN(n595) );
  NAND2_X1 U688 ( .A1(n473), .A2(n595), .ZN(n681) );
  NAND2_X1 U689 ( .A1(n790), .A2(n681), .ZN(n596) );
  INV_X1 U690 ( .A(n596), .ZN(n598) );
  NOR2_X1 U691 ( .A1(n392), .A2(KEYINPUT44), .ZN(n597) );
  NAND2_X1 U692 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U693 ( .A(KEYINPUT64), .B(KEYINPUT83), .ZN(n600) );
  XOR2_X1 U694 ( .A(KEYINPUT101), .B(n602), .Z(n603) );
  NOR2_X1 U695 ( .A1(G900), .A2(n603), .ZN(n604) );
  NOR2_X1 U696 ( .A1(n605), .A2(n604), .ZN(n614) );
  NOR2_X1 U697 ( .A1(n616), .A2(n716), .ZN(n607) );
  XNOR2_X1 U698 ( .A(KEYINPUT30), .B(n607), .ZN(n608) );
  NAND2_X1 U699 ( .A1(n609), .A2(n608), .ZN(n627) );
  XNOR2_X1 U700 ( .A(KEYINPUT38), .B(n610), .ZN(n717) );
  XNOR2_X1 U701 ( .A(KEYINPUT84), .B(KEYINPUT39), .ZN(n611) );
  NOR2_X1 U702 ( .A1(n614), .A2(n704), .ZN(n615) );
  NAND2_X1 U703 ( .A1(n615), .A2(n355), .ZN(n639) );
  NOR2_X1 U704 ( .A1(n616), .A2(n639), .ZN(n618) );
  XNOR2_X1 U705 ( .A(KEYINPUT28), .B(KEYINPUT102), .ZN(n617) );
  XNOR2_X1 U706 ( .A(n618), .B(n617), .ZN(n619) );
  XOR2_X1 U707 ( .A(KEYINPUT103), .B(n620), .Z(n630) );
  XOR2_X1 U708 ( .A(KEYINPUT41), .B(KEYINPUT104), .Z(n622) );
  NOR2_X1 U709 ( .A1(n717), .A2(n716), .ZN(n720) );
  NAND2_X1 U710 ( .A1(n720), .A2(n718), .ZN(n621) );
  NOR2_X1 U711 ( .A1(n630), .A2(n729), .ZN(n625) );
  XOR2_X1 U712 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n623) );
  XNOR2_X1 U713 ( .A(KEYINPUT42), .B(n623), .ZN(n624) );
  NOR2_X1 U714 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U715 ( .A1(n628), .A2(n610), .ZN(n688) );
  NOR2_X1 U716 ( .A1(n630), .A2(n629), .ZN(n683) );
  AND2_X1 U717 ( .A1(n683), .A2(n721), .ZN(n631) );
  NOR2_X1 U718 ( .A1(KEYINPUT81), .A2(n631), .ZN(n632) );
  NOR2_X1 U719 ( .A1(KEYINPUT47), .A2(n632), .ZN(n633) );
  OR2_X1 U720 ( .A1(KEYINPUT81), .A2(n721), .ZN(n634) );
  NAND2_X1 U721 ( .A1(n634), .A2(n683), .ZN(n635) );
  NAND2_X1 U722 ( .A1(n635), .A2(KEYINPUT47), .ZN(n637) );
  NAND2_X1 U723 ( .A1(n721), .A2(KEYINPUT81), .ZN(n636) );
  NAND2_X1 U724 ( .A1(n637), .A2(n636), .ZN(n645) );
  NOR2_X1 U725 ( .A1(n691), .A2(n639), .ZN(n640) );
  NAND2_X1 U726 ( .A1(n640), .A2(n397), .ZN(n651) );
  NOR2_X1 U727 ( .A1(n638), .A2(n651), .ZN(n642) );
  XNOR2_X1 U728 ( .A(KEYINPUT107), .B(KEYINPUT36), .ZN(n641) );
  XNOR2_X1 U729 ( .A(n642), .B(n641), .ZN(n644) );
  NOR2_X1 U730 ( .A1(n644), .A2(n643), .ZN(n697) );
  NOR2_X1 U731 ( .A1(n645), .A2(n697), .ZN(n646) );
  NAND2_X1 U732 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U733 ( .A(n649), .B(n383), .ZN(n659) );
  NOR2_X1 U734 ( .A1(n650), .A2(n695), .ZN(n700) );
  NOR2_X1 U735 ( .A1(n390), .A2(n651), .ZN(n652) );
  NAND2_X1 U736 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U737 ( .A(KEYINPUT43), .B(n654), .ZN(n656) );
  NAND2_X1 U738 ( .A1(n656), .A2(n385), .ZN(n701) );
  INV_X1 U739 ( .A(KEYINPUT2), .ZN(n661) );
  OR2_X1 U740 ( .A1(n661), .A2(KEYINPUT75), .ZN(n660) );
  NAND2_X1 U741 ( .A1(KEYINPUT75), .A2(n661), .ZN(n662) );
  INV_X1 U742 ( .A(KEYINPUT120), .ZN(n666) );
  NAND2_X1 U743 ( .A1(n740), .A2(G472), .ZN(n670) );
  INV_X1 U744 ( .A(KEYINPUT63), .ZN(n672) );
  XOR2_X1 U745 ( .A(G101), .B(n673), .Z(G3) );
  NOR2_X1 U746 ( .A1(n691), .A2(n675), .ZN(n674) );
  XOR2_X1 U747 ( .A(G104), .B(n674), .Z(G6) );
  NOR2_X1 U748 ( .A1(n695), .A2(n675), .ZN(n680) );
  XOR2_X1 U749 ( .A(KEYINPUT109), .B(KEYINPUT27), .Z(n677) );
  XNOR2_X1 U750 ( .A(G107), .B(KEYINPUT26), .ZN(n676) );
  XNOR2_X1 U751 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U752 ( .A(KEYINPUT108), .B(n678), .ZN(n679) );
  XNOR2_X1 U753 ( .A(n680), .B(n679), .ZN(G9) );
  XNOR2_X1 U754 ( .A(G110), .B(KEYINPUT110), .ZN(n682) );
  XNOR2_X1 U755 ( .A(n682), .B(n681), .ZN(G12) );
  INV_X1 U756 ( .A(n683), .ZN(n689) );
  NOR2_X1 U757 ( .A1(n689), .A2(n695), .ZN(n687) );
  XOR2_X1 U758 ( .A(KEYINPUT111), .B(KEYINPUT29), .Z(n685) );
  XNOR2_X1 U759 ( .A(G128), .B(KEYINPUT112), .ZN(n684) );
  XNOR2_X1 U760 ( .A(n685), .B(n684), .ZN(n686) );
  XNOR2_X1 U761 ( .A(n687), .B(n686), .ZN(G30) );
  XNOR2_X1 U762 ( .A(n412), .B(n688), .ZN(G45) );
  NOR2_X1 U763 ( .A1(n691), .A2(n689), .ZN(n690) );
  XOR2_X1 U764 ( .A(G146), .B(n690), .Z(G48) );
  NOR2_X1 U765 ( .A1(n691), .A2(n694), .ZN(n692) );
  XOR2_X1 U766 ( .A(n693), .B(n692), .Z(G15) );
  NOR2_X1 U767 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U768 ( .A(G116), .B(n696), .Z(G18) );
  XOR2_X1 U769 ( .A(KEYINPUT37), .B(KEYINPUT113), .Z(n699) );
  XNOR2_X1 U770 ( .A(G125), .B(n697), .ZN(n698) );
  XNOR2_X1 U771 ( .A(n699), .B(n698), .ZN(G27) );
  XOR2_X1 U772 ( .A(G134), .B(n700), .Z(G36) );
  XNOR2_X1 U773 ( .A(G140), .B(n701), .ZN(G42) );
  OR2_X1 U774 ( .A1(n702), .A2(n390), .ZN(n703) );
  XNOR2_X1 U775 ( .A(KEYINPUT50), .B(n703), .ZN(n708) );
  NOR2_X1 U776 ( .A1(n415), .A2(n355), .ZN(n706) );
  XNOR2_X1 U777 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n705) );
  XNOR2_X1 U778 ( .A(n706), .B(n705), .ZN(n707) );
  NAND2_X1 U779 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U780 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U781 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U782 ( .A(n713), .B(KEYINPUT115), .ZN(n714) );
  XNOR2_X1 U783 ( .A(KEYINPUT51), .B(n714), .ZN(n715) );
  NOR2_X1 U784 ( .A1(n729), .A2(n715), .ZN(n725) );
  NAND2_X1 U785 ( .A1(n717), .A2(n716), .ZN(n719) );
  NAND2_X1 U786 ( .A1(n719), .A2(n718), .ZN(n723) );
  NAND2_X1 U787 ( .A1(n721), .A2(n720), .ZN(n722) );
  AND2_X1 U788 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U789 ( .A1(n725), .A2(n380), .ZN(n726) );
  XNOR2_X1 U790 ( .A(n726), .B(KEYINPUT52), .ZN(n727) );
  NOR2_X1 U791 ( .A1(n728), .A2(n727), .ZN(n731) );
  NOR2_X1 U792 ( .A1(n731), .A2(n730), .ZN(n733) );
  XNOR2_X1 U793 ( .A(n736), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U794 ( .A(KEYINPUT55), .B(KEYINPUT54), .Z(n739) );
  XNOR2_X1 U795 ( .A(n737), .B(KEYINPUT117), .ZN(n738) );
  XNOR2_X1 U796 ( .A(n739), .B(n738), .ZN(n742) );
  XNOR2_X1 U797 ( .A(KEYINPUT56), .B(n744), .ZN(G51) );
  XOR2_X1 U798 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n746) );
  NAND2_X1 U799 ( .A1(n366), .A2(G469), .ZN(n745) );
  NOR2_X1 U800 ( .A1(n760), .A2(n748), .ZN(G54) );
  NAND2_X1 U801 ( .A1(n740), .A2(G475), .ZN(n752) );
  XOR2_X1 U802 ( .A(KEYINPUT118), .B(KEYINPUT59), .Z(n749) );
  XNOR2_X1 U803 ( .A(n754), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U804 ( .A(n755), .B(KEYINPUT119), .Z(n758) );
  NAND2_X1 U805 ( .A1(n366), .A2(G478), .ZN(n757) );
  XNOR2_X1 U806 ( .A(n758), .B(n757), .ZN(n759) );
  NOR2_X1 U807 ( .A1(n760), .A2(n759), .ZN(G63) );
  INV_X1 U808 ( .A(G898), .ZN(n763) );
  NAND2_X1 U809 ( .A1(G953), .A2(G224), .ZN(n761) );
  XOR2_X1 U810 ( .A(KEYINPUT61), .B(n761), .Z(n762) );
  NOR2_X1 U811 ( .A1(n763), .A2(n762), .ZN(n765) );
  NOR2_X1 U812 ( .A1(G953), .A2(n372), .ZN(n764) );
  NOR2_X1 U813 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U814 ( .A(n766), .B(KEYINPUT125), .ZN(n773) );
  XOR2_X1 U815 ( .A(KEYINPUT124), .B(KEYINPUT123), .Z(n769) );
  XNOR2_X1 U816 ( .A(n365), .B(G110), .ZN(n768) );
  XNOR2_X1 U817 ( .A(n769), .B(n768), .ZN(n771) );
  NOR2_X1 U818 ( .A1(G898), .A2(n782), .ZN(n770) );
  NOR2_X1 U819 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U820 ( .A(n773), .B(n772), .ZN(n774) );
  XNOR2_X1 U821 ( .A(KEYINPUT122), .B(n774), .ZN(G69) );
  XNOR2_X1 U822 ( .A(n371), .B(n775), .ZN(n781) );
  XNOR2_X1 U823 ( .A(G227), .B(n781), .ZN(n777) );
  NAND2_X1 U824 ( .A1(n777), .A2(G900), .ZN(n778) );
  NAND2_X1 U825 ( .A1(G953), .A2(n778), .ZN(n779) );
  XNOR2_X1 U826 ( .A(n779), .B(KEYINPUT126), .ZN(n785) );
  XNOR2_X1 U827 ( .A(n781), .B(n780), .ZN(n783) );
  NAND2_X1 U828 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U829 ( .A1(n785), .A2(n784), .ZN(G72) );
  XOR2_X1 U830 ( .A(n392), .B(G122), .Z(G24) );
  XOR2_X1 U831 ( .A(G137), .B(n787), .Z(G39) );
  XNOR2_X1 U832 ( .A(G131), .B(KEYINPUT127), .ZN(n789) );
  XNOR2_X1 U833 ( .A(n789), .B(n788), .ZN(G33) );
  XNOR2_X1 U834 ( .A(G119), .B(n790), .ZN(G21) );
endmodule

