//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 0 0 1 0 0 0 1 1 0 0 0 0 0 1 1 0 1 1 0 0 1 0 0 1 1 1 0 0 0 1 0 0 0 0 0 1 1 1 0 0 0 0 0 1 0 0 1 1 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n822, new_n824, new_n825, new_n826, new_n827, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951;
  INV_X1    g000(.A(KEYINPUT82), .ZN(new_n202));
  XOR2_X1   g001(.A(G155gat), .B(G162gat), .Z(new_n203));
  INV_X1    g002(.A(KEYINPUT76), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G155gat), .B(G162gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT76), .ZN(new_n207));
  INV_X1    g006(.A(G155gat), .ZN(new_n208));
  INV_X1    g007(.A(G162gat), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT2), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  XOR2_X1   g009(.A(G141gat), .B(G148gat), .Z(new_n211));
  NAND4_X1  g010(.A1(new_n205), .A2(new_n207), .A3(new_n210), .A4(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(KEYINPUT75), .ZN(new_n214));
  XNOR2_X1  g013(.A(G141gat), .B(G148gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT75), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT2), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n206), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT3), .B1(new_n213), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n214), .A2(new_n217), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(new_n203), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(new_n222), .A3(new_n212), .ZN(new_n223));
  INV_X1    g022(.A(G120gat), .ZN(new_n224));
  OR3_X1    g023(.A1(new_n224), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT69), .B1(new_n224), .B2(G113gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(KEYINPUT68), .B(G120gat), .ZN(new_n227));
  INV_X1    g026(.A(G113gat), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n225), .B(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT1), .ZN(new_n230));
  INV_X1    g029(.A(G127gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G134gat), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n231), .A2(G134gat), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n229), .A2(new_n230), .A3(new_n232), .A4(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT67), .B(G134gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n232), .B1(new_n235), .B2(new_n231), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n224), .A2(G113gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n228), .A2(G120gat), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n230), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n234), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n219), .A2(new_n223), .A3(new_n241), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n213), .A2(new_n218), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n234), .A2(new_n240), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n243), .A2(new_n244), .A3(KEYINPUT4), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n221), .A2(new_n212), .A3(new_n234), .A4(new_n240), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT4), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n242), .A2(new_n245), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(G225gat), .A2(G233gat), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT39), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n221), .A2(new_n212), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(new_n241), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT77), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(new_n256), .A3(new_n246), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n254), .A2(KEYINPUT77), .A3(new_n241), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n251), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n253), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G1gat), .B(G29gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(KEYINPUT0), .ZN(new_n262));
  XNOR2_X1  g061(.A(G57gat), .B(G85gat), .ZN(new_n263));
  XOR2_X1   g062(.A(new_n262), .B(new_n263), .Z(new_n264));
  OAI21_X1  g063(.A(new_n264), .B1(new_n252), .B2(KEYINPUT39), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n202), .B1(new_n260), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT40), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n257), .A2(new_n251), .A3(new_n258), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT78), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n242), .A2(new_n245), .A3(new_n250), .A4(new_n248), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n257), .A2(KEYINPUT78), .A3(new_n251), .A4(new_n258), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n270), .A2(KEYINPUT5), .A3(new_n271), .A4(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT79), .B1(new_n271), .B2(KEYINPUT5), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  AND3_X1   g075(.A1(new_n272), .A2(KEYINPUT5), .A3(new_n271), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n277), .A2(new_n274), .A3(new_n270), .ZN(new_n278));
  INV_X1    g077(.A(new_n264), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n276), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT40), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n202), .B(new_n281), .C1(new_n260), .C2(new_n265), .ZN(new_n282));
  AND3_X1   g081(.A1(new_n267), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G211gat), .B(G218gat), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT22), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT72), .B(G211gat), .ZN(new_n286));
  INV_X1    g085(.A(G218gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G197gat), .B(G204gat), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n284), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n290), .A2(new_n291), .A3(new_n284), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G226gat), .ZN(new_n296));
  INV_X1    g095(.A(G233gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n298), .A2(KEYINPUT29), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(KEYINPUT27), .B(G183gat), .ZN(new_n301));
  INV_X1    g100(.A(G190gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT28), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT65), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n301), .B(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n302), .A2(KEYINPUT28), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n305), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OR3_X1    g108(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n311));
  INV_X1    g110(.A(G169gat), .ZN(new_n312));
  INV_X1    g111(.A(G176gat), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n310), .B(new_n311), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(G183gat), .A2(G190gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n314), .A2(KEYINPUT66), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n315), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT66), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n309), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT64), .B1(new_n312), .B2(new_n313), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n321), .B(KEYINPUT23), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(new_n315), .ZN(new_n324));
  NAND3_X1  g123(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n325));
  AOI22_X1  g124(.A1(new_n324), .A2(new_n325), .B1(G169gat), .B2(G176gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT25), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n322), .A2(KEYINPUT25), .A3(new_n326), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n320), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT74), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT74), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n320), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n300), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n298), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n295), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n294), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n340), .A2(new_n292), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n332), .A2(new_n299), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n333), .A2(new_n335), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n341), .B(new_n342), .C1(new_n343), .C2(new_n337), .ZN(new_n344));
  XNOR2_X1  g143(.A(G8gat), .B(G36gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(G64gat), .B(G92gat), .ZN(new_n346));
  XOR2_X1   g145(.A(new_n345), .B(new_n346), .Z(new_n347));
  NAND3_X1  g146(.A1(new_n339), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT30), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n347), .B1(new_n339), .B2(new_n344), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n339), .A2(new_n344), .A3(KEYINPUT30), .A4(new_n347), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n350), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G78gat), .B(G106gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(G50gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n356), .B(KEYINPUT80), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n357), .B(KEYINPUT31), .Z(new_n358));
  INV_X1    g157(.A(G22gat), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT29), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n360), .B1(new_n340), .B2(new_n292), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n243), .B1(new_n361), .B2(new_n222), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n295), .B1(new_n360), .B2(new_n223), .ZN(new_n363));
  INV_X1    g162(.A(G228gat), .ZN(new_n364));
  OAI22_X1  g163(.A1(new_n362), .A2(new_n363), .B1(new_n364), .B2(new_n297), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT29), .B1(new_n293), .B2(new_n294), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n254), .B1(new_n366), .B2(KEYINPUT3), .ZN(new_n367));
  INV_X1    g166(.A(new_n223), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n341), .B1(KEYINPUT29), .B2(new_n368), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n367), .A2(G228gat), .A3(G233gat), .A4(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n359), .B1(new_n365), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT81), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n358), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n365), .A2(new_n370), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(G22gat), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n365), .A2(new_n370), .A3(new_n359), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n375), .A2(new_n372), .A3(new_n376), .A4(new_n358), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n283), .A2(new_n354), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n348), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT37), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n347), .A2(new_n382), .ZN(new_n383));
  OR2_X1    g182(.A1(new_n351), .A2(new_n383), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n295), .B(new_n342), .C1(new_n343), .C2(new_n337), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n385), .A2(KEYINPUT37), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n341), .B1(new_n336), .B2(new_n338), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT38), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n381), .B1(new_n384), .B2(new_n388), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n273), .A2(new_n275), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n274), .B1(new_n277), .B2(new_n270), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n264), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT6), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(new_n393), .A3(new_n280), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n351), .A2(new_n383), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n382), .B1(new_n339), .B2(new_n344), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT38), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n276), .A2(new_n278), .A3(KEYINPUT6), .A4(new_n279), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n389), .A2(new_n394), .A3(new_n397), .A4(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n394), .A2(new_n398), .ZN(new_n400));
  INV_X1    g199(.A(new_n354), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n378), .A2(new_n379), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n380), .A2(new_n399), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n320), .A2(new_n331), .A3(new_n244), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT70), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n332), .A2(new_n241), .ZN(new_n407));
  NAND2_X1  g206(.A1(G227gat), .A2(G233gat), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT70), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n320), .A2(new_n331), .A3(new_n409), .A4(new_n244), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n406), .A2(new_n407), .A3(new_n408), .A4(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(KEYINPUT34), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT32), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n406), .A2(new_n407), .A3(new_n410), .ZN(new_n414));
  INV_X1    g213(.A(new_n408), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT33), .B1(new_n414), .B2(new_n415), .ZN(new_n417));
  XOR2_X1   g216(.A(G15gat), .B(G43gat), .Z(new_n418));
  XNOR2_X1  g217(.A(G71gat), .B(G99gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NOR3_X1   g220(.A1(new_n416), .A2(new_n417), .A3(new_n421), .ZN(new_n422));
  AOI221_X4 g221(.A(new_n413), .B1(KEYINPUT33), .B2(new_n420), .C1(new_n414), .C2(new_n415), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n412), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n417), .A2(new_n421), .ZN(new_n425));
  INV_X1    g224(.A(new_n416), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n412), .ZN(new_n428));
  INV_X1    g227(.A(new_n423), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n424), .A2(new_n430), .A3(KEYINPUT71), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT71), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n432), .B(new_n412), .C1(new_n422), .C2(new_n423), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n431), .A2(new_n433), .A3(KEYINPUT36), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n424), .A2(new_n430), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT36), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n431), .A2(new_n433), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n354), .B1(new_n394), .B2(new_n398), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n378), .A2(new_n379), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT35), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT35), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n440), .A2(new_n441), .A3(new_n444), .A4(new_n435), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n404), .A2(new_n438), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  AND2_X1   g245(.A1(G43gat), .A2(G50gat), .ZN(new_n447));
  NOR2_X1   g246(.A1(G43gat), .A2(G50gat), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT83), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(G43gat), .ZN(new_n450));
  INV_X1    g249(.A(G50gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT83), .ZN(new_n453));
  NAND2_X1  g252(.A1(G43gat), .A2(G50gat), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n449), .A2(new_n455), .A3(KEYINPUT15), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT15), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n452), .A2(new_n457), .A3(new_n454), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT14), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n459), .B1(G29gat), .B2(G36gat), .ZN(new_n460));
  NAND2_X1  g259(.A1(G29gat), .A2(G36gat), .ZN(new_n461));
  NOR2_X1   g260(.A1(G29gat), .A2(G36gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT14), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n458), .A2(new_n460), .A3(new_n461), .A4(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT84), .B1(new_n456), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n455), .A3(KEYINPUT15), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT84), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n463), .A2(new_n460), .A3(new_n461), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n466), .A2(new_n467), .A3(new_n468), .A4(new_n458), .ZN(new_n469));
  INV_X1    g268(.A(new_n468), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n456), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n465), .A2(KEYINPUT17), .A3(new_n469), .A4(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT88), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n466), .A2(new_n468), .A3(new_n458), .ZN(new_n474));
  AOI22_X1  g273(.A1(new_n474), .A2(KEYINPUT84), .B1(new_n456), .B2(new_n470), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT88), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n475), .A2(new_n476), .A3(KEYINPUT17), .A4(new_n469), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n359), .A2(G15gat), .ZN(new_n479));
  INV_X1    g278(.A(G15gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(G22gat), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT16), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n479), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n479), .A2(new_n481), .A3(KEYINPUT86), .ZN(new_n484));
  INV_X1    g283(.A(G1gat), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(G15gat), .B(G22gat), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n487), .B(KEYINPUT86), .C1(new_n482), .C2(G1gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(KEYINPUT87), .B(G8gat), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n486), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n486), .A2(new_n488), .ZN(new_n491));
  NOR2_X1   g290(.A1(KEYINPUT87), .A2(G8gat), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n465), .A2(new_n469), .A3(new_n471), .ZN(new_n494));
  XOR2_X1   g293(.A(KEYINPUT85), .B(KEYINPUT17), .Z(new_n495));
  AOI21_X1  g294(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n478), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n494), .A2(new_n493), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT18), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n499), .B1(G229gat), .B2(G233gat), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n497), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT89), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n502), .B1(new_n494), .B2(new_n493), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n492), .B1(new_n486), .B2(new_n488), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n504), .B1(new_n491), .B2(new_n489), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n505), .A2(new_n475), .A3(KEYINPUT89), .A4(new_n469), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n503), .A2(new_n506), .A3(new_n498), .ZN(new_n507));
  NAND2_X1  g306(.A1(G229gat), .A2(G233gat), .ZN(new_n508));
  XOR2_X1   g307(.A(new_n508), .B(KEYINPUT13), .Z(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n501), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n498), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n512), .B1(new_n478), .B2(new_n496), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT18), .B1(new_n513), .B2(new_n508), .ZN(new_n514));
  XNOR2_X1  g313(.A(G113gat), .B(G141gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(G197gat), .ZN(new_n516));
  XOR2_X1   g315(.A(KEYINPUT11), .B(G169gat), .Z(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(new_n517), .ZN(new_n518));
  XOR2_X1   g317(.A(new_n518), .B(KEYINPUT12), .Z(new_n519));
  NOR3_X1   g318(.A1(new_n511), .A2(new_n514), .A3(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n519), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n497), .A2(new_n508), .A3(new_n498), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(new_n499), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n513), .A2(new_n500), .B1(new_n509), .B2(new_n507), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(G57gat), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n527), .A2(G64gat), .ZN(new_n528));
  INV_X1    g327(.A(G64gat), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n529), .A2(G57gat), .ZN(new_n530));
  OAI22_X1  g329(.A1(new_n528), .A2(new_n530), .B1(KEYINPUT90), .B2(KEYINPUT9), .ZN(new_n531));
  INV_X1    g330(.A(G71gat), .ZN(new_n532));
  INV_X1    g331(.A(G78gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OR3_X1    g333(.A1(new_n532), .A2(new_n533), .A3(KEYINPUT90), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT90), .B1(new_n532), .B2(new_n533), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n531), .A2(new_n534), .A3(new_n535), .A4(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n532), .A2(new_n533), .A3(KEYINPUT9), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n538), .B1(new_n532), .B2(new_n533), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n527), .A2(KEYINPUT91), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT91), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(G57gat), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n540), .A2(new_n542), .A3(G64gat), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT92), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n544), .B1(new_n527), .B2(G64gat), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n529), .A2(KEYINPUT92), .A3(G57gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n539), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n537), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT21), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(G231gat), .A2(G233gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  OR2_X1    g352(.A1(new_n553), .A2(new_n231), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n231), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n505), .B1(new_n550), .B2(new_n549), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n554), .A2(new_n557), .A3(new_n555), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(new_n208), .ZN(new_n563));
  XNOR2_X1  g362(.A(G183gat), .B(G211gat), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n563), .B(new_n564), .Z(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n559), .A2(new_n560), .A3(new_n565), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G99gat), .A2(G106gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(KEYINPUT8), .ZN(new_n571));
  NAND2_X1  g370(.A1(G85gat), .A2(G92gat), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT7), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(G85gat), .ZN(new_n575));
  INV_X1    g374(.A(G92gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n571), .A2(new_n574), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G99gat), .B(G106gat), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  AOI22_X1  g381(.A1(KEYINPUT8), .A2(new_n570), .B1(new_n575), .B2(new_n576), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n583), .A2(new_n580), .A3(new_n574), .A4(new_n578), .ZN(new_n584));
  AOI21_X1  g383(.A(KEYINPUT94), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n584), .A2(KEYINPUT94), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n587), .B1(new_n494), .B2(new_n495), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n478), .A2(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(G232gat), .A2(G233gat), .ZN(new_n590));
  AOI22_X1  g389(.A1(new_n494), .A2(new_n587), .B1(KEYINPUT41), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(G190gat), .B(G218gat), .Z(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n590), .A2(KEYINPUT41), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT93), .ZN(new_n596));
  XNOR2_X1  g395(.A(G134gat), .B(G162gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n593), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n589), .A2(new_n599), .A3(new_n591), .ZN(new_n600));
  AND3_X1   g399(.A1(new_n594), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n598), .B1(new_n594), .B2(new_n600), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n569), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n549), .B1(new_n585), .B2(new_n586), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n537), .A2(new_n548), .A3(new_n584), .A4(new_n582), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT10), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n587), .A2(KEYINPUT10), .A3(new_n548), .A4(new_n537), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G230gat), .A2(G233gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n611), .B(KEYINPUT95), .Z(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n605), .A2(new_n606), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(new_n612), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G120gat), .B(G148gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(G176gat), .B(G204gat), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n619), .B(new_n620), .Z(new_n621));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n621), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n617), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NOR4_X1   g424(.A1(new_n446), .A2(new_n526), .A3(new_n604), .A4(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n400), .B(KEYINPUT96), .Z(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n354), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT42), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT16), .B(G8gat), .ZN(new_n632));
  OR3_X1    g431(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n630), .A2(G8gat), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n631), .B1(new_n630), .B2(new_n632), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(G1325gat));
  INV_X1    g435(.A(new_n626), .ZN(new_n637));
  OAI21_X1  g436(.A(G15gat), .B1(new_n637), .B2(new_n438), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n626), .A2(new_n480), .A3(new_n435), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(G1326gat));
  OR3_X1    g439(.A1(new_n637), .A2(KEYINPUT97), .A3(new_n441), .ZN(new_n641));
  OAI21_X1  g440(.A(KEYINPUT97), .B1(new_n637), .B2(new_n441), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT43), .B(G22gat), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n643), .B1(new_n641), .B2(new_n642), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n644), .A2(new_n645), .ZN(G1327gat));
  NAND2_X1  g445(.A1(new_n443), .A2(new_n445), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n283), .A2(new_n354), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n399), .A2(new_n441), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n402), .A2(new_n403), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n438), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n526), .ZN(new_n653));
  INV_X1    g452(.A(new_n569), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n601), .A2(new_n602), .ZN(new_n655));
  INV_X1    g454(.A(new_n625), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT98), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n400), .B(KEYINPUT96), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n659), .A2(G29gat), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n652), .A2(new_n653), .A3(new_n658), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT45), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n663), .B1(new_n446), .B2(new_n603), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n652), .A2(KEYINPUT44), .A3(new_n655), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n625), .B(KEYINPUT99), .Z(new_n666));
  NOR3_X1   g465(.A1(new_n666), .A2(new_n569), .A3(new_n526), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n664), .A2(new_n665), .A3(new_n627), .A4(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(G29gat), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n662), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT100), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(G1328gat));
  NOR2_X1   g471(.A1(new_n446), .A2(new_n526), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n658), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n674), .A2(G36gat), .A3(new_n401), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT46), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n664), .A2(new_n665), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n677), .A2(new_n354), .A3(new_n667), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT101), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(G36gat), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n678), .A2(new_n679), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n676), .B1(new_n681), .B2(new_n682), .ZN(G1329gat));
  INV_X1    g482(.A(new_n435), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n450), .B1(new_n674), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n677), .A2(new_n667), .ZN(new_n686));
  INV_X1    g485(.A(new_n438), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(G43gat), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n685), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT102), .B(KEYINPUT47), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  OAI211_X1 g491(.A(new_n685), .B(new_n690), .C1(new_n686), .C2(new_n688), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(G1330gat));
  NAND4_X1  g493(.A1(new_n673), .A2(new_n451), .A3(new_n403), .A4(new_n658), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n695), .A2(KEYINPUT104), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n664), .A2(new_n665), .A3(new_n403), .A4(new_n667), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(G50gat), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n695), .A2(KEYINPUT104), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n696), .A2(new_n698), .A3(KEYINPUT48), .A4(new_n699), .ZN(new_n700));
  OR2_X1    g499(.A1(new_n695), .A2(KEYINPUT103), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n695), .A2(KEYINPUT103), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n701), .A2(new_n698), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n700), .B1(new_n703), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g503(.A(new_n666), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n705), .A2(new_n653), .A3(new_n604), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n652), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(new_n659), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT105), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n540), .A2(new_n542), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1332gat));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n707), .B(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n354), .B(KEYINPUT107), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n715), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT108), .B1(new_n713), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n707), .B(KEYINPUT106), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT108), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n719), .A2(new_n720), .A3(new_n716), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n718), .A2(new_n723), .A3(new_n721), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(G1333gat));
  NAND3_X1  g526(.A1(new_n719), .A2(G71gat), .A3(new_n687), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n532), .B1(new_n707), .B2(new_n684), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n728), .A2(KEYINPUT50), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT50), .B1(new_n728), .B2(new_n729), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(G1334gat));
  NAND2_X1  g531(.A1(new_n719), .A2(new_n403), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g533(.A1(new_n653), .A2(new_n569), .A3(new_n656), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n664), .A2(new_n665), .A3(new_n627), .A4(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(G85gat), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n603), .B1(new_n647), .B2(new_n651), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n653), .A2(new_n569), .ZN(new_n739));
  AOI21_X1  g538(.A(KEYINPUT51), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n740), .A2(KEYINPUT109), .ZN(new_n741));
  INV_X1    g540(.A(new_n740), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n738), .A2(KEYINPUT51), .A3(new_n739), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n741), .B1(new_n744), .B2(KEYINPUT109), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n627), .A2(new_n575), .A3(new_n625), .ZN(new_n746));
  OAI211_X1 g545(.A(KEYINPUT110), .B(new_n737), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT110), .ZN(new_n748));
  INV_X1    g547(.A(new_n741), .ZN(new_n749));
  AND3_X1   g548(.A1(new_n738), .A2(KEYINPUT51), .A3(new_n739), .ZN(new_n750));
  OAI21_X1  g549(.A(KEYINPUT109), .B1(new_n750), .B2(new_n740), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n746), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n737), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n748), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n747), .A2(new_n754), .ZN(G1336gat));
  NAND4_X1  g554(.A1(new_n664), .A2(new_n665), .A3(new_n714), .A4(new_n735), .ZN(new_n756));
  AOI21_X1  g555(.A(KEYINPUT52), .B1(new_n756), .B2(G92gat), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n714), .A2(new_n576), .A3(new_n666), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n757), .B1(new_n745), .B2(new_n758), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n664), .A2(new_n665), .A3(new_n354), .A4(new_n735), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(G92gat), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n758), .B(KEYINPUT111), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(new_n750), .B2(new_n740), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT112), .B1(new_n764), .B2(KEYINPUT52), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT112), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767));
  AOI211_X1 g566(.A(new_n766), .B(new_n767), .C1(new_n761), .C2(new_n763), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n759), .B1(new_n765), .B2(new_n768), .ZN(G1337gat));
  NAND3_X1  g568(.A1(new_n677), .A2(new_n687), .A3(new_n735), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(G99gat), .ZN(new_n771));
  OR3_X1    g570(.A1(new_n684), .A2(G99gat), .A3(new_n656), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n745), .B2(new_n772), .ZN(G1338gat));
  OR3_X1    g572(.A1(new_n441), .A2(new_n705), .A3(G106gat), .ZN(new_n774));
  XOR2_X1   g573(.A(new_n774), .B(KEYINPUT113), .Z(new_n775));
  NOR2_X1   g574(.A1(new_n745), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n664), .A2(new_n665), .A3(new_n403), .A4(new_n735), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(G106gat), .ZN(new_n778));
  XNOR2_X1  g577(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n781));
  INV_X1    g580(.A(new_n775), .ZN(new_n782));
  AOI22_X1  g581(.A1(new_n744), .A2(new_n782), .B1(new_n777), .B2(G106gat), .ZN(new_n783));
  OAI22_X1  g582(.A1(new_n776), .A2(new_n780), .B1(new_n781), .B2(new_n783), .ZN(G1339gat));
  NAND3_X1  g583(.A1(new_n608), .A2(new_n609), .A3(new_n612), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n608), .A2(new_n609), .A3(KEYINPUT115), .A4(new_n612), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n787), .A2(new_n614), .A3(KEYINPUT54), .A4(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n612), .B1(new_n608), .B2(new_n609), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n621), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AOI211_X1 g594(.A(new_n794), .B(new_n621), .C1(new_n790), .C2(new_n791), .ZN(new_n796));
  AOI22_X1  g595(.A1(new_n796), .A2(new_n789), .B1(new_n618), .B2(new_n621), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n795), .B(new_n797), .C1(new_n601), .C2(new_n602), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n523), .A2(new_n524), .A3(new_n521), .ZN(new_n799));
  OAI22_X1  g598(.A1(new_n513), .A2(new_n508), .B1(new_n509), .B2(new_n507), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n518), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n799), .A2(KEYINPUT116), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT116), .B1(new_n799), .B2(new_n801), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n798), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n795), .B(new_n797), .C1(new_n520), .C2(new_n525), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n625), .A2(new_n799), .A3(new_n801), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n655), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n654), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n569), .A2(new_n526), .A3(new_n603), .A4(new_n656), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n403), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n811), .A2(new_n627), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n714), .A2(new_n684), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n814), .A2(new_n228), .A3(new_n526), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n812), .A2(new_n439), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(new_n653), .A3(new_n715), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n815), .B1(new_n818), .B2(new_n228), .ZN(G1340gat));
  OAI21_X1  g618(.A(G120gat), .B1(new_n814), .B2(new_n705), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n817), .A2(new_n715), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n656), .A2(new_n227), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(G1341gat));
  NAND4_X1  g622(.A1(new_n812), .A2(G127gat), .A3(new_n569), .A4(new_n813), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n824), .A2(KEYINPUT117), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n824), .A2(KEYINPUT117), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n817), .A2(new_n569), .A3(new_n715), .ZN(new_n827));
  AOI211_X1 g626(.A(new_n825), .B(new_n826), .C1(new_n231), .C2(new_n827), .ZN(G1342gat));
  NOR2_X1   g627(.A1(new_n354), .A2(new_n603), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  OR3_X1    g629(.A1(new_n816), .A2(new_n235), .A3(new_n830), .ZN(new_n831));
  OR2_X1    g630(.A1(new_n831), .A2(KEYINPUT56), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(KEYINPUT56), .ZN(new_n833));
  OAI21_X1  g632(.A(G134gat), .B1(new_n814), .B2(new_n603), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(KEYINPUT118), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT118), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n832), .A2(new_n833), .A3(new_n837), .A4(new_n834), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(G1343gat));
  AOI21_X1  g638(.A(new_n441), .B1(new_n809), .B2(new_n810), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(KEYINPUT57), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n687), .A2(new_n659), .A3(new_n714), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n844), .A2(G141gat), .A3(new_n653), .ZN(new_n845));
  INV_X1    g644(.A(new_n842), .ZN(new_n846));
  INV_X1    g645(.A(new_n840), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n846), .A2(new_n526), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n845), .B1(G141gat), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT58), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n849), .B(new_n850), .ZN(G1344gat));
  NOR2_X1   g650(.A1(new_n846), .A2(new_n847), .ZN(new_n852));
  INV_X1    g651(.A(G148gat), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n852), .A2(new_n853), .A3(new_n625), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n656), .B1(new_n846), .B2(KEYINPUT119), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n797), .A2(new_n795), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n807), .B1(new_n526), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n603), .ZN(new_n859));
  INV_X1    g658(.A(new_n804), .ZN(new_n860));
  INV_X1    g659(.A(new_n857), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n860), .A2(new_n861), .A3(new_n655), .A4(new_n802), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n569), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n810), .ZN(new_n864));
  OAI211_X1 g663(.A(KEYINPUT57), .B(new_n403), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n865), .A2(KEYINPUT120), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT120), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n867), .B1(new_n840), .B2(KEYINPUT57), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n809), .A2(new_n810), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n441), .B1(new_n870), .B2(KEYINPUT121), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n809), .A2(new_n872), .A3(new_n810), .ZN(new_n873));
  AOI21_X1  g672(.A(KEYINPUT57), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  OAI221_X1 g673(.A(new_n856), .B1(KEYINPUT119), .B2(new_n846), .C1(new_n869), .C2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n855), .B1(new_n875), .B2(G148gat), .ZN(new_n876));
  AOI211_X1 g675(.A(KEYINPUT59), .B(new_n853), .C1(new_n844), .C2(new_n625), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n854), .B1(new_n876), .B2(new_n877), .ZN(G1345gat));
  OAI21_X1  g677(.A(G155gat), .B1(new_n843), .B2(new_n654), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n852), .A2(new_n208), .A3(new_n569), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(G1346gat));
  OAI21_X1  g680(.A(G162gat), .B1(new_n843), .B2(new_n603), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n659), .A2(G162gat), .A3(new_n830), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n883), .A2(new_n438), .A3(new_n840), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(G1347gat));
  NAND2_X1  g684(.A1(new_n659), .A2(new_n354), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n435), .A3(new_n811), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n888), .B(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n653), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n891), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n892));
  AOI21_X1  g691(.A(KEYINPUT123), .B1(new_n891), .B2(G169gat), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n870), .A2(new_n659), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n894), .A2(new_n441), .A3(new_n439), .A4(new_n714), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n653), .A2(new_n312), .ZN(new_n896));
  OAI22_X1  g695(.A1(new_n892), .A2(new_n893), .B1(new_n895), .B2(new_n896), .ZN(G1348gat));
  NAND3_X1  g696(.A1(new_n890), .A2(G176gat), .A3(new_n666), .ZN(new_n898));
  OR2_X1    g697(.A1(new_n898), .A2(KEYINPUT124), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n313), .B1(new_n895), .B2(new_n656), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n898), .A2(KEYINPUT124), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(G1349gat));
  XNOR2_X1  g701(.A(new_n888), .B(KEYINPUT122), .ZN(new_n903));
  OAI21_X1  g702(.A(G183gat), .B1(new_n903), .B2(new_n654), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT125), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n905), .A2(KEYINPUT60), .ZN(new_n906));
  OR3_X1    g705(.A1(new_n895), .A2(new_n307), .A3(new_n654), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n904), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n906), .B1(new_n904), .B2(new_n907), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(G1350gat));
  AOI21_X1  g709(.A(new_n302), .B1(new_n890), .B2(new_n655), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT61), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n911), .A2(new_n912), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n655), .A2(new_n302), .ZN(new_n915));
  OAI22_X1  g714(.A1(new_n913), .A2(new_n914), .B1(new_n895), .B2(new_n915), .ZN(G1351gat));
  NOR3_X1   g715(.A1(new_n687), .A2(new_n715), .A3(new_n441), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n894), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n918), .A2(G197gat), .A3(new_n526), .ZN(new_n919));
  XOR2_X1   g718(.A(new_n919), .B(KEYINPUT126), .Z(new_n920));
  NAND2_X1  g719(.A1(new_n887), .A2(new_n438), .ZN(new_n921));
  OAI21_X1  g720(.A(KEYINPUT121), .B1(new_n863), .B2(new_n864), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(new_n403), .A3(new_n873), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT57), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n865), .A2(KEYINPUT120), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n840), .A2(new_n867), .A3(KEYINPUT57), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n921), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(G197gat), .B1(new_n930), .B2(new_n526), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n920), .A2(new_n931), .ZN(G1352gat));
  NOR3_X1   g731(.A1(new_n918), .A2(G204gat), .A3(new_n656), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT62), .ZN(new_n934));
  OAI21_X1  g733(.A(G204gat), .B1(new_n930), .B2(new_n705), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1353gat));
  INV_X1    g735(.A(new_n918), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n937), .A2(new_n286), .A3(new_n569), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT63), .ZN(new_n939));
  INV_X1    g738(.A(G211gat), .ZN(new_n940));
  AOI211_X1 g739(.A(new_n939), .B(new_n940), .C1(new_n929), .C2(new_n569), .ZN(new_n941));
  INV_X1    g740(.A(new_n921), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n569), .B(new_n942), .C1(new_n869), .C2(new_n874), .ZN(new_n943));
  AOI21_X1  g742(.A(KEYINPUT63), .B1(new_n943), .B2(G211gat), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n938), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(KEYINPUT127), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT127), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n947), .B(new_n938), .C1(new_n941), .C2(new_n944), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n948), .ZN(G1354gat));
  OAI21_X1  g748(.A(G218gat), .B1(new_n930), .B2(new_n603), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n937), .A2(new_n287), .A3(new_n655), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(G1355gat));
endmodule


