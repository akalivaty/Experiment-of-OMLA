//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 1 1 1 0 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n444, new_n445, new_n449, new_n451, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n616, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1245,
    new_n1246, new_n1247;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  INV_X1    g017(.A(G2072), .ZN(new_n443));
  INV_X1    g018(.A(G2078), .ZN(new_n444));
  NOR2_X1   g019(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g020(.A1(new_n445), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  NAND2_X1  g023(.A1(G94), .A2(G452), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g027(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g028(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT2), .Z(new_n456));
  NAND4_X1  g031(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT67), .Z(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI211_X1 g042(.A(G137), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n467), .A2(new_n472), .ZN(G160));
  OR2_X1    g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n462), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n463), .A2(new_n464), .ZN(new_n479));
  OAI21_X1  g054(.A(KEYINPUT69), .B1(new_n479), .B2(new_n462), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  AOI21_X1  g057(.A(G2105), .B1(new_n474), .B2(new_n475), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT68), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n487));
  AND3_X1   g062(.A1(new_n482), .A2(new_n485), .A3(new_n487), .ZN(G162));
  AND2_X1   g063(.A1(KEYINPUT70), .A2(G138), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n462), .B(new_n489), .C1(new_n463), .C2(new_n464), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g067(.A(KEYINPUT3), .B(G2104), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .A3(new_n462), .A4(new_n489), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n493), .A2(G126), .A3(G2105), .ZN(new_n495));
  OR2_X1    g070(.A1(new_n462), .A2(G114), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n492), .A2(new_n494), .A3(new_n495), .A4(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  XNOR2_X1  g076(.A(KEYINPUT6), .B(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G50), .ZN(new_n504));
  AND3_X1   g079(.A1(KEYINPUT71), .A2(KEYINPUT5), .A3(G543), .ZN(new_n505));
  AOI21_X1  g080(.A(KEYINPUT5), .B1(KEYINPUT71), .B2(G543), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n505), .A2(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT72), .B(G88), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n503), .A2(new_n504), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  OAI21_X1  g087(.A(G62), .B1(new_n505), .B2(new_n506), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n511), .A2(new_n515), .ZN(G166));
  NAND2_X1  g091(.A1(KEYINPUT71), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(KEYINPUT71), .A2(KEYINPUT5), .A3(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(G51), .ZN(new_n525));
  OAI211_X1 g100(.A(new_n522), .B(new_n524), .C1(new_n525), .C2(new_n503), .ZN(new_n526));
  INV_X1    g101(.A(new_n509), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n527), .A2(G89), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n526), .A2(new_n528), .ZN(G168));
  AOI22_X1  g104(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n512), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT73), .B(G52), .ZN(new_n532));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n503), .A2(new_n532), .B1(new_n509), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n531), .A2(new_n534), .ZN(G171));
  AOI22_X1  g110(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n512), .ZN(new_n537));
  INV_X1    g112(.A(G43), .ZN(new_n538));
  INV_X1    g113(.A(G81), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n503), .A2(new_n538), .B1(new_n509), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  NAND4_X1  g117(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g118(.A1(G1), .A2(G3), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT74), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(G188));
  INV_X1    g122(.A(KEYINPUT77), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n502), .A2(G53), .A3(G543), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(KEYINPUT9), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT9), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n502), .A2(new_n551), .A3(G53), .A4(G543), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n509), .A2(KEYINPUT75), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n521), .A2(new_n555), .A3(new_n502), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n554), .A2(G91), .A3(new_n556), .ZN(new_n557));
  AND2_X1   g132(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g133(.A(G65), .B1(new_n505), .B2(new_n506), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G651), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT76), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT76), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n561), .A2(new_n564), .A3(G651), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n548), .B1(new_n558), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n564), .B1(new_n561), .B2(G651), .ZN(new_n568));
  AOI211_X1 g143(.A(KEYINPUT76), .B(new_n512), .C1(new_n559), .C2(new_n560), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n553), .A2(new_n557), .ZN(new_n571));
  NOR3_X1   g146(.A1(new_n570), .A2(new_n571), .A3(KEYINPUT77), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n567), .A2(new_n572), .ZN(G299));
  INV_X1    g148(.A(G171), .ZN(G301));
  INV_X1    g149(.A(G168), .ZN(G286));
  INV_X1    g150(.A(G166), .ZN(G303));
  NOR2_X1   g151(.A1(new_n505), .A2(new_n506), .ZN(new_n577));
  INV_X1    g152(.A(G74), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n512), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n503), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n579), .B1(G49), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n554), .A2(G87), .A3(new_n556), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G288));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G61), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n577), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n586), .A2(G651), .B1(new_n580), .B2(G48), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n554), .A2(G86), .A3(new_n556), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(G305));
  AOI22_X1  g164(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(new_n512), .ZN(new_n591));
  INV_X1    g166(.A(G47), .ZN(new_n592));
  INV_X1    g167(.A(G85), .ZN(new_n593));
  OAI22_X1  g168(.A1(new_n503), .A2(new_n592), .B1(new_n509), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G290));
  INV_X1    g171(.A(G868), .ZN(new_n597));
  NOR2_X1   g172(.A1(G301), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n577), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G651), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n580), .A2(G54), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n554), .A2(G92), .A3(new_n556), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g182(.A1(new_n554), .A2(new_n556), .A3(KEYINPUT10), .A4(G92), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n604), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT78), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n598), .B1(new_n610), .B2(new_n597), .ZN(G284));
  AOI21_X1  g186(.A(new_n598), .B1(new_n610), .B2(new_n597), .ZN(G321));
  NAND2_X1  g187(.A1(G299), .A2(new_n597), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(new_n597), .B2(G168), .ZN(G297));
  OAI21_X1  g189(.A(new_n613), .B1(new_n597), .B2(G168), .ZN(G280));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n610), .B1(new_n616), .B2(G860), .ZN(G148));
  OAI21_X1  g192(.A(new_n597), .B1(new_n537), .B2(new_n540), .ZN(new_n618));
  AND2_X1   g193(.A1(new_n610), .A2(new_n616), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n597), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n493), .A2(new_n470), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT12), .Z(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT13), .Z(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n625), .A2(G2100), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n481), .A2(G123), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT79), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(G111), .ZN(new_n631));
  AOI22_X1  g206(.A1(new_n628), .A2(new_n629), .B1(new_n631), .B2(G2105), .ZN(new_n632));
  AOI22_X1  g207(.A1(new_n630), .A2(new_n632), .B1(new_n483), .B2(G135), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n627), .A2(new_n633), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n634), .A2(G2096), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n625), .A2(G2100), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(G2096), .ZN(new_n637));
  NAND4_X1  g212(.A1(new_n626), .A2(new_n635), .A3(new_n636), .A4(new_n637), .ZN(G156));
  INV_X1    g213(.A(G14), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  INV_X1    g215(.A(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2427), .B(G2430), .Z(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT80), .B(KEYINPUT14), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n642), .A2(new_n643), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2443), .B(G2446), .Z(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AND2_X1   g224(.A1(new_n646), .A2(new_n645), .ZN(new_n650));
  INV_X1    g225(.A(new_n648), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(new_n651), .A3(new_n644), .ZN(new_n652));
  XOR2_X1   g227(.A(G2451), .B(G2454), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT81), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n649), .A2(new_n652), .A3(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n655), .B1(new_n649), .B2(new_n652), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n639), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n649), .A2(new_n652), .ZN(new_n662));
  INV_X1    g237(.A(new_n655), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(new_n656), .ZN(new_n665));
  INV_X1    g240(.A(new_n660), .ZN(new_n666));
  AOI21_X1  g241(.A(KEYINPUT82), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT82), .ZN(new_n668));
  AOI211_X1 g243(.A(new_n668), .B(new_n660), .C1(new_n664), .C2(new_n656), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n661), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G401));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT83), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(KEYINPUT18), .ZN(new_n676));
  NOR2_X1   g251(.A1(G2072), .A2(G2078), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n676), .B1(new_n445), .B2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT84), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT18), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n675), .A2(KEYINPUT17), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n673), .A2(new_n674), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G2096), .B(G2100), .Z(new_n685));
  XOR2_X1   g260(.A(new_n684), .B(new_n685), .Z(new_n686));
  NAND2_X1  g261(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n684), .B(new_n685), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(new_n679), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n687), .A2(new_n689), .ZN(G227));
  XOR2_X1   g265(.A(G1991), .B(G1996), .Z(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1956), .B(G2474), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT85), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G1961), .B(G1966), .Z(new_n696));
  OR2_X1    g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1971), .B(G1976), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT19), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n695), .A2(new_n696), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n697), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  OR3_X1    g276(.A1(new_n699), .A2(new_n695), .A3(new_n696), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(new_n700), .B2(new_n699), .ZN(new_n706));
  INV_X1    g281(.A(new_n699), .ZN(new_n707));
  NAND4_X1  g282(.A1(new_n707), .A2(new_n695), .A3(new_n696), .A4(new_n704), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n692), .B1(new_n703), .B2(new_n709), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n709), .A2(new_n702), .A3(new_n701), .ZN(new_n711));
  INV_X1    g286(.A(new_n692), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n691), .B1(new_n710), .B2(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(G1981), .B(G1986), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n703), .A2(new_n709), .A3(new_n692), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n711), .A2(new_n712), .ZN(new_n717));
  INV_X1    g292(.A(new_n691), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  AND3_X1   g294(.A1(new_n714), .A2(new_n715), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n715), .B1(new_n714), .B2(new_n719), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(G229));
  INV_X1    g298(.A(G16), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G6), .ZN(new_n725));
  INV_X1    g300(.A(G305), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(new_n724), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT89), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT32), .B(G1981), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n728), .A2(new_n730), .ZN(new_n732));
  INV_X1    g307(.A(G288), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(new_n724), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n724), .B2(G23), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT33), .B(G1976), .Z(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n724), .A2(G22), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G166), .B2(new_n724), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G1971), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n735), .B2(new_n737), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n731), .A2(new_n732), .A3(new_n738), .A4(new_n742), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n743), .A2(KEYINPUT34), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(KEYINPUT34), .ZN(new_n745));
  INV_X1    g320(.A(G29), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G25), .ZN(new_n747));
  OAI21_X1  g322(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n748));
  INV_X1    g323(.A(G107), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(G2105), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT87), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G131), .B2(new_n483), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n481), .A2(G119), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n747), .B1(new_n755), .B2(new_n746), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT35), .B(G1991), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT88), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n756), .A2(new_n758), .B1(KEYINPUT90), .B2(KEYINPUT36), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n758), .B2(new_n756), .ZN(new_n760));
  NOR2_X1   g335(.A1(G16), .A2(G24), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n595), .B2(G16), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G1986), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n744), .A2(new_n745), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT25), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n483), .A2(G139), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n493), .A2(G127), .ZN(new_n774));
  NAND2_X1  g349(.A1(G115), .A2(G2104), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n462), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT92), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR3_X1   g354(.A1(new_n773), .A2(new_n776), .A3(KEYINPUT92), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n781), .A2(new_n746), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n746), .B2(G33), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n783), .A2(new_n443), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n443), .ZN(new_n785));
  AND3_X1   g360(.A1(new_n478), .A2(new_n480), .A3(G129), .ZN(new_n786));
  NAND3_X1  g361(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT26), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n483), .A2(G141), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n470), .A2(G105), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n786), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n792), .A2(new_n746), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n746), .B2(G32), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT27), .B(G1996), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT93), .B(KEYINPUT24), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G34), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n797), .A2(G29), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G29), .B2(G160), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n794), .A2(new_n795), .B1(G2084), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n784), .A2(new_n785), .A3(new_n800), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT94), .ZN(new_n802));
  NOR2_X1   g377(.A1(G29), .A2(G35), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G162), .B2(G29), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT29), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(G2090), .Z(new_n806));
  NOR2_X1   g381(.A1(new_n799), .A2(G2084), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT95), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n746), .A2(G26), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT28), .Z(new_n810));
  NOR2_X1   g385(.A1(G104), .A2(G2105), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT91), .Z(new_n812));
  INV_X1    g387(.A(G116), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n469), .B1(new_n813), .B2(G2105), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n812), .A2(new_n814), .B1(G140), .B2(new_n483), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n478), .A2(new_n480), .A3(G128), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n810), .B1(new_n817), .B2(G29), .ZN(new_n818));
  INV_X1    g393(.A(G2067), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n724), .A2(G19), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n541), .B2(new_n724), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G1341), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n808), .A2(new_n820), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n724), .A2(G21), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(G168), .B2(new_n724), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n724), .A2(G5), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(G171), .B2(new_n724), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n826), .A2(G1966), .B1(new_n828), .B2(G1961), .ZN(new_n829));
  OAI221_X1 g404(.A(new_n829), .B1(G1961), .B2(new_n828), .C1(new_n794), .C2(new_n795), .ZN(new_n830));
  NOR2_X1   g405(.A1(G27), .A2(G29), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(G164), .B2(G29), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(G2078), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n826), .A2(G1966), .ZN(new_n834));
  INV_X1    g409(.A(G28), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n835), .A2(KEYINPUT30), .ZN(new_n836));
  AOI21_X1  g411(.A(G29), .B1(new_n835), .B2(KEYINPUT30), .ZN(new_n837));
  OR2_X1    g412(.A1(KEYINPUT31), .A2(G11), .ZN(new_n838));
  NAND2_X1  g413(.A1(KEYINPUT31), .A2(G11), .ZN(new_n839));
  AOI22_X1  g414(.A1(new_n836), .A2(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n634), .B2(new_n746), .ZN(new_n841));
  NOR4_X1   g416(.A1(new_n830), .A2(new_n833), .A3(new_n834), .A4(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n806), .A2(new_n824), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n724), .A2(G4), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n610), .B2(new_n724), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(G1348), .ZN(new_n846));
  NOR3_X1   g421(.A1(new_n802), .A2(new_n843), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(G299), .A2(G16), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n724), .A2(G20), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT23), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT96), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(G1956), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n767), .A2(new_n768), .A3(new_n847), .A4(new_n853), .ZN(G150));
  INV_X1    g429(.A(G150), .ZN(G311));
  NAND2_X1  g430(.A1(new_n610), .A2(G559), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT38), .ZN(new_n857));
  AOI22_X1  g432(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n858), .A2(new_n512), .ZN(new_n859));
  INV_X1    g434(.A(G55), .ZN(new_n860));
  XOR2_X1   g435(.A(KEYINPUT97), .B(G93), .Z(new_n861));
  OAI22_X1  g436(.A1(new_n503), .A2(new_n860), .B1(new_n509), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n541), .A2(new_n863), .ZN(new_n864));
  OAI22_X1  g439(.A1(new_n537), .A2(new_n540), .B1(new_n859), .B2(new_n862), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n857), .B(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT39), .ZN(new_n868));
  AOI21_X1  g443(.A(G860), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n869), .B1(new_n868), .B2(new_n867), .ZN(new_n870));
  INV_X1    g445(.A(new_n863), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(G860), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n872), .B(KEYINPUT37), .Z(new_n873));
  NAND2_X1  g448(.A1(new_n870), .A2(new_n873), .ZN(G145));
  XNOR2_X1  g449(.A(new_n634), .B(G160), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n875), .B(G162), .Z(new_n876));
  NAND2_X1  g451(.A1(new_n792), .A2(new_n817), .ZN(new_n877));
  OAI211_X1 g452(.A(new_n816), .B(new_n815), .C1(new_n786), .C2(new_n791), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n500), .A2(KEYINPUT98), .ZN(new_n880));
  AOI22_X1  g455(.A1(new_n476), .A2(G126), .B1(new_n496), .B2(new_n498), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT98), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n881), .A2(new_n882), .A3(new_n494), .A4(new_n492), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n879), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(KEYINPUT99), .B1(new_n779), .B2(new_n780), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n877), .A2(new_n880), .A3(new_n883), .A4(new_n878), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT99), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(new_n889), .A3(new_n781), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n478), .A2(new_n480), .A3(G130), .ZN(new_n891));
  OAI21_X1  g466(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n892));
  INV_X1    g467(.A(G118), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n892), .B1(new_n893), .B2(G2105), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n894), .B1(G142), .B2(new_n483), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(KEYINPUT100), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT100), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n891), .A2(new_n898), .A3(new_n895), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n623), .ZN(new_n901));
  INV_X1    g476(.A(new_n623), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n897), .A2(new_n902), .A3(new_n899), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n755), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n901), .A2(new_n903), .A3(new_n754), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n781), .A2(new_n889), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n885), .A2(new_n907), .A3(new_n886), .A4(new_n887), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n890), .A2(new_n905), .A3(new_n906), .A4(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n905), .A2(new_n906), .ZN(new_n910));
  INV_X1    g485(.A(new_n781), .ZN(new_n911));
  AOI211_X1 g486(.A(KEYINPUT99), .B(new_n911), .C1(new_n885), .C2(new_n887), .ZN(new_n912));
  INV_X1    g487(.A(new_n908), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n876), .B1(new_n909), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n915), .A2(G37), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n909), .A2(new_n914), .A3(new_n876), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g494(.A1(new_n871), .A2(new_n597), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n619), .B(new_n866), .ZN(new_n921));
  INV_X1    g496(.A(new_n609), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n922), .B1(new_n567), .B2(new_n572), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n558), .A2(new_n566), .A3(new_n548), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT77), .B1(new_n570), .B2(new_n571), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n924), .A2(new_n925), .A3(new_n609), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT101), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT41), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n924), .A2(new_n925), .A3(new_n609), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n609), .B1(new_n924), .B2(new_n925), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n923), .A2(KEYINPUT41), .A3(new_n926), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n933), .A2(new_n934), .A3(KEYINPUT101), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n921), .A2(new_n930), .A3(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n927), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n936), .B1(new_n921), .B2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(G305), .B(new_n595), .ZN(new_n939));
  XNOR2_X1  g514(.A(G288), .B(G166), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XOR2_X1   g518(.A(new_n943), .B(KEYINPUT42), .Z(new_n944));
  XNOR2_X1  g519(.A(new_n938), .B(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n920), .B1(new_n945), .B2(new_n597), .ZN(G295));
  OAI21_X1  g521(.A(new_n920), .B1(new_n945), .B2(new_n597), .ZN(G331));
  INV_X1    g522(.A(KEYINPUT102), .ZN(new_n948));
  OAI21_X1  g523(.A(G171), .B1(G286), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n948), .B1(new_n526), .B2(new_n528), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n864), .A2(new_n865), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n950), .B1(new_n864), .B2(new_n865), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n950), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n866), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(G301), .B1(KEYINPUT102), .B2(G168), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n864), .A2(new_n865), .A3(new_n950), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n953), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n959), .A2(new_n937), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n960), .A2(new_n943), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n935), .A2(new_n930), .A3(new_n959), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G37), .ZN(new_n964));
  AOI22_X1  g539(.A1(new_n933), .A2(new_n934), .B1(new_n958), .B2(new_n953), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n943), .B1(new_n960), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n963), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT103), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT43), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n966), .A2(new_n964), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT103), .B1(new_n970), .B2(new_n963), .ZN(new_n971));
  OAI21_X1  g546(.A(KEYINPUT104), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n967), .A2(new_n968), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n970), .A2(KEYINPUT103), .A3(new_n963), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT104), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n973), .A2(new_n974), .A3(new_n975), .A4(KEYINPUT43), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n977));
  INV_X1    g552(.A(new_n960), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n962), .ZN(new_n979));
  AOI21_X1  g554(.A(G37), .B1(new_n979), .B2(new_n943), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT43), .B1(new_n961), .B2(new_n962), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n977), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n972), .A2(new_n976), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n970), .A2(new_n981), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n961), .A2(new_n962), .ZN(new_n985));
  INV_X1    g560(.A(new_n943), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n986), .B1(new_n978), .B2(new_n962), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n985), .A2(new_n987), .A3(G37), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT43), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n984), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n977), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n983), .A2(new_n991), .ZN(G397));
  INV_X1    g567(.A(G1384), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n880), .A2(new_n993), .A3(new_n883), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G125), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n997), .B1(new_n474), .B2(new_n475), .ZN(new_n998));
  INV_X1    g573(.A(new_n466), .ZN(new_n999));
  OAI21_X1  g574(.A(G2105), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n1000), .A2(G40), .A3(new_n471), .A4(new_n468), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT105), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT105), .ZN(new_n1003));
  NAND3_X1  g578(.A1(G160), .A2(new_n1003), .A3(G40), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n996), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G1996), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n1007), .A2(new_n1008), .A3(new_n792), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT106), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n817), .B(new_n819), .ZN(new_n1013));
  INV_X1    g588(.A(new_n792), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1013), .B1(G1996), .B2(new_n1014), .ZN(new_n1015));
  AOI22_X1  g590(.A1(new_n1011), .A2(new_n1012), .B1(new_n1006), .B2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g591(.A(new_n754), .B(new_n758), .Z(new_n1017));
  OAI21_X1  g592(.A(new_n1016), .B1(new_n1007), .B2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g593(.A(new_n595), .B(G1986), .Z(new_n1019));
  AOI21_X1  g594(.A(new_n1018), .B1(new_n1006), .B2(new_n1019), .ZN(new_n1020));
  AND2_X1   g595(.A1(new_n500), .A2(new_n993), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1021), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1022));
  XOR2_X1   g597(.A(KEYINPUT108), .B(G8), .Z(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n581), .A2(G1976), .A3(new_n582), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1022), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT52), .ZN(new_n1027));
  XOR2_X1   g602(.A(KEYINPUT109), .B(G1976), .Z(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT52), .B1(G288), .B2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1029), .A2(new_n1022), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT49), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n586), .A2(G651), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n527), .A2(G86), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n580), .A2(G48), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT110), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1036), .A2(new_n1037), .A3(G1981), .ZN(new_n1038));
  INV_X1    g613(.A(G1981), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n587), .A2(new_n1039), .A3(new_n588), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1037), .B1(new_n1036), .B2(G1981), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1032), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1042), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1044), .A2(KEYINPUT49), .A3(new_n1040), .A4(new_n1038), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1003), .B1(G160), .B2(G40), .ZN(new_n1046));
  INV_X1    g621(.A(G40), .ZN(new_n1047));
  NOR4_X1   g622(.A1(new_n467), .A2(new_n472), .A3(KEYINPUT105), .A4(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1023), .B1(new_n1049), .B2(new_n1021), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1043), .A2(new_n1045), .A3(new_n1050), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n1031), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(G8), .B1(new_n511), .B2(new_n515), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  OAI211_X1 g630(.A(KEYINPUT55), .B(G8), .C1(new_n511), .C2(new_n515), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT45), .B1(new_n500), .B2(new_n993), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n1059), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n880), .A2(KEYINPUT45), .A3(new_n993), .A4(new_n883), .ZN(new_n1061));
  AOI21_X1  g636(.A(G1971), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n500), .A2(new_n993), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT50), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT50), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n500), .A2(new_n1065), .A3(new_n993), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1064), .A2(new_n1002), .A3(new_n1004), .A4(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1067), .A2(G2090), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1062), .A2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1058), .B1(new_n1069), .B2(new_n1023), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT107), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n1055), .A2(new_n1071), .A3(new_n1056), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1071), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1074), .B(G8), .C1(new_n1062), .C2(new_n1068), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1052), .A2(new_n1070), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1059), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1049), .A2(new_n1061), .A3(new_n444), .A4(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g653(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n1079));
  XOR2_X1   g654(.A(KEYINPUT120), .B(G1961), .Z(new_n1080));
  AOI22_X1  g655(.A1(new_n1078), .A2(new_n1079), .B1(new_n1067), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n993), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1049), .A2(new_n444), .A3(new_n1077), .A4(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT53), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n993), .ZN(new_n1086));
  NOR3_X1   g661(.A1(new_n1005), .A2(new_n1059), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT119), .B1(new_n1087), .B2(new_n444), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1081), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1089), .A2(KEYINPUT122), .A3(G171), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(G171), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1076), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT51), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1049), .A2(new_n1077), .A3(new_n1082), .ZN(new_n1096));
  INV_X1    g671(.A(G1966), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G2084), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1049), .A2(new_n1099), .A3(new_n1066), .A4(new_n1064), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1023), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1095), .B1(new_n1101), .B2(G286), .ZN(new_n1102));
  AOI21_X1  g677(.A(G1966), .B1(new_n1060), .B2(new_n1082), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1067), .A2(G2084), .ZN(new_n1104));
  OAI211_X1 g679(.A(KEYINPUT118), .B(G8), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(G286), .A2(new_n1024), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT118), .B1(new_n1108), .B2(G8), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1102), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1101), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1111), .A2(new_n1095), .A3(new_n1106), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT62), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1110), .A2(KEYINPUT62), .A3(new_n1112), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1094), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(G1976), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1051), .A2(new_n1118), .A3(new_n733), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n1040), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1075), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1120), .A2(new_n1050), .B1(new_n1052), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1067), .A2(new_n1080), .ZN(new_n1124));
  OAI21_X1  g699(.A(KEYINPUT53), .B1(KEYINPUT123), .B2(G2078), .ZN(new_n1125));
  AOI211_X1 g700(.A(new_n1125), .B(new_n1001), .C1(KEYINPUT123), .C2(G2078), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1126), .A2(new_n996), .A3(new_n1061), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1123), .A2(G301), .A3(new_n1124), .A4(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT124), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT124), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1081), .A2(new_n1130), .A3(G301), .A4(new_n1127), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1093), .A2(new_n1132), .A3(new_n1090), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT54), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1075), .A2(new_n1031), .A3(new_n1051), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1049), .A2(new_n1061), .A3(new_n1077), .ZN(new_n1137));
  INV_X1    g712(.A(G1971), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1139), .B1(G2090), .B2(new_n1067), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1057), .B1(new_n1140), .B2(new_n1024), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1136), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1123), .A2(new_n1124), .A3(new_n1127), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(G171), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1144), .B(KEYINPUT54), .C1(new_n1089), .C2(G171), .ZN(new_n1145));
  AND4_X1   g720(.A1(new_n1142), .A2(new_n1110), .A3(new_n1145), .A4(new_n1112), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1135), .A2(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g722(.A(KEYINPUT56), .B(G2072), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1049), .A2(new_n1061), .A3(new_n1077), .A4(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT114), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1060), .A2(KEYINPUT114), .A3(new_n1061), .A4(new_n1148), .ZN(new_n1152));
  INV_X1    g727(.A(G1956), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1067), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT57), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n558), .A2(new_n566), .A3(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(KEYINPUT57), .B1(new_n570), .B2(new_n571), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1151), .A2(new_n1152), .A3(new_n1154), .A4(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1158), .A2(KEYINPUT115), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT115), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1156), .A2(new_n1157), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  AND4_X1   g739(.A1(new_n1049), .A2(new_n1061), .A3(new_n1077), .A4(new_n1148), .ZN(new_n1165));
  AOI22_X1  g740(.A1(new_n1165), .A2(KEYINPUT114), .B1(new_n1153), .B2(new_n1067), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1164), .B1(new_n1166), .B2(new_n1151), .ZN(new_n1167));
  INV_X1    g742(.A(G1348), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1067), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1049), .A2(new_n819), .A3(new_n1021), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n922), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  OAI211_X1 g746(.A(KEYINPUT116), .B(new_n1160), .C1(new_n1167), .C2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT116), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1151), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1163), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1162), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1171), .B1(new_n1174), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1160), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1173), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1172), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1169), .A2(KEYINPUT60), .A3(new_n1170), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1182), .A2(KEYINPUT117), .A3(new_n922), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n922), .B1(new_n1182), .B2(KEYINPUT117), .ZN(new_n1184));
  OAI22_X1  g759(.A1(new_n1183), .A2(new_n1184), .B1(KEYINPUT117), .B2(new_n1182), .ZN(new_n1185));
  AND2_X1   g760(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1186));
  OR2_X1    g761(.A1(new_n1186), .A2(KEYINPUT60), .ZN(new_n1187));
  XOR2_X1   g762(.A(KEYINPUT58), .B(G1341), .Z(new_n1188));
  NAND2_X1  g763(.A1(new_n1022), .A2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1189), .B1(new_n1137), .B2(G1996), .ZN(new_n1190));
  AND2_X1   g765(.A1(new_n1190), .A2(new_n541), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT59), .ZN(new_n1192));
  OR2_X1    g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1194));
  AOI22_X1  g769(.A1(new_n1185), .A2(new_n1187), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1174), .A2(new_n1158), .ZN(new_n1196));
  AOI21_X1  g771(.A(KEYINPUT61), .B1(new_n1196), .B2(new_n1160), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1167), .ZN(new_n1198));
  AND2_X1   g773(.A1(new_n1160), .A2(KEYINPUT61), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1197), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1181), .B1(new_n1195), .B2(new_n1200), .ZN(new_n1201));
  OAI211_X1 g776(.A(new_n1117), .B(new_n1122), .C1(new_n1147), .C2(new_n1201), .ZN(new_n1202));
  INV_X1    g777(.A(G8), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n1069), .A2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1058), .B1(new_n1204), .B2(KEYINPUT113), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1205), .B1(KEYINPUT113), .B2(new_n1204), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1111), .A2(G286), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1207), .A2(KEYINPUT63), .ZN(new_n1208));
  NOR3_X1   g783(.A1(new_n1206), .A2(new_n1136), .A3(new_n1208), .ZN(new_n1209));
  AND2_X1   g784(.A1(new_n1142), .A2(new_n1207), .ZN(new_n1210));
  OR2_X1    g785(.A1(new_n1210), .A2(KEYINPUT111), .ZN(new_n1211));
  XOR2_X1   g786(.A(KEYINPUT112), .B(KEYINPUT63), .Z(new_n1212));
  AOI21_X1  g787(.A(new_n1212), .B1(new_n1210), .B2(KEYINPUT111), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1209), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1020), .B1(new_n1202), .B2(new_n1214), .ZN(new_n1215));
  NOR2_X1   g790(.A1(new_n817), .A2(G2067), .ZN(new_n1216));
  NOR2_X1   g791(.A1(new_n754), .A2(new_n758), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1216), .B1(new_n1016), .B2(new_n1217), .ZN(new_n1218));
  NOR3_X1   g793(.A1(new_n1007), .A2(G1986), .A3(G290), .ZN(new_n1219));
  XNOR2_X1  g794(.A(new_n1219), .B(KEYINPUT48), .ZN(new_n1220));
  OAI22_X1  g795(.A1(new_n1218), .A2(new_n1007), .B1(new_n1018), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT46), .ZN(new_n1223));
  NOR2_X1   g798(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  XOR2_X1   g799(.A(new_n1224), .B(KEYINPUT126), .Z(new_n1225));
  NAND2_X1  g800(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1226));
  XOR2_X1   g801(.A(new_n1226), .B(KEYINPUT125), .Z(new_n1227));
  AOI21_X1  g802(.A(new_n1007), .B1(new_n792), .B2(new_n1013), .ZN(new_n1228));
  OR3_X1    g803(.A1(new_n1225), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  OR2_X1    g804(.A1(new_n1229), .A2(KEYINPUT47), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1229), .A2(KEYINPUT47), .ZN(new_n1231));
  AOI21_X1  g806(.A(new_n1221), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g807(.A1(new_n1215), .A2(new_n1232), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g808(.A(KEYINPUT127), .ZN(new_n1235));
  AND3_X1   g809(.A1(new_n687), .A2(new_n689), .A3(G319), .ZN(new_n1236));
  OAI211_X1 g810(.A(new_n1236), .B(new_n670), .C1(new_n720), .C2(new_n721), .ZN(new_n1237));
  AOI21_X1  g811(.A(new_n1237), .B1(new_n916), .B2(new_n917), .ZN(new_n1238));
  AOI21_X1  g812(.A(new_n1235), .B1(new_n990), .B2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g813(.A(new_n989), .B1(new_n980), .B2(new_n963), .ZN(new_n1240));
  AND3_X1   g814(.A1(new_n981), .A2(new_n964), .A3(new_n966), .ZN(new_n1241));
  OAI211_X1 g815(.A(new_n1238), .B(new_n1235), .C1(new_n1240), .C2(new_n1241), .ZN(new_n1242));
  INV_X1    g816(.A(new_n1242), .ZN(new_n1243));
  NOR2_X1   g817(.A1(new_n1239), .A2(new_n1243), .ZN(G308));
  NOR2_X1   g818(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1245));
  INV_X1    g819(.A(new_n1238), .ZN(new_n1246));
  OAI21_X1  g820(.A(KEYINPUT127), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g821(.A1(new_n1247), .A2(new_n1242), .ZN(G225));
endmodule


