//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 1 0 0 0 1 1 0 1 0 1 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 0 1 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n658, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(G143), .B(G146), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT0), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n189), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT72), .B(G125), .ZN(new_n193));
  XOR2_X1   g007(.A(KEYINPUT0), .B(G128), .Z(new_n194));
  OAI211_X1 g008(.A(new_n192), .B(new_n193), .C1(new_n189), .C2(new_n194), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n191), .A2(KEYINPUT1), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G143), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G146), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n196), .A2(new_n198), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT72), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT72), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G125), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n191), .A2(new_n197), .A3(G143), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n199), .B(G146), .C1(new_n191), .C2(KEYINPUT1), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n201), .A2(new_n206), .A3(new_n207), .A4(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n195), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT78), .B(G224), .ZN(new_n211));
  INV_X1    g025(.A(G953), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XOR2_X1   g027(.A(new_n210), .B(new_n213), .Z(new_n214));
  XOR2_X1   g028(.A(G116), .B(G119), .Z(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT2), .B(G113), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XOR2_X1   g031(.A(KEYINPUT2), .B(G113), .Z(new_n218));
  XNOR2_X1  g032(.A(G116), .B(G119), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G104), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT3), .B1(new_n222), .B2(G107), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n224));
  INV_X1    g038(.A(G107), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(new_n225), .A3(G104), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n222), .A2(G107), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n223), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT4), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(new_n229), .A3(G101), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n228), .A2(G101), .ZN(new_n231));
  XOR2_X1   g045(.A(KEYINPUT75), .B(G101), .Z(new_n232));
  OAI21_X1  g046(.A(KEYINPUT4), .B1(new_n228), .B2(new_n232), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n221), .B(new_n230), .C1(new_n231), .C2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT5), .ZN(new_n235));
  INV_X1    g049(.A(G119), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(new_n236), .A3(G116), .ZN(new_n237));
  OAI211_X1 g051(.A(G113), .B(new_n237), .C1(new_n215), .C2(new_n235), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT75), .B(G101), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n239), .A2(new_n227), .A3(new_n226), .A4(new_n223), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n225), .A2(G104), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n222), .A2(G107), .ZN(new_n242));
  OAI21_X1  g056(.A(G101), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n238), .A2(new_n220), .A3(new_n240), .A4(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n234), .A2(new_n244), .ZN(new_n245));
  XOR2_X1   g059(.A(G110), .B(G122), .Z(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n246), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n234), .A2(new_n248), .A3(new_n244), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n247), .A2(KEYINPUT6), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT77), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT6), .ZN(new_n252));
  AND4_X1   g066(.A1(new_n251), .A2(new_n245), .A3(new_n252), .A4(new_n246), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n248), .B1(new_n234), .B2(new_n244), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n251), .B1(new_n254), .B2(new_n252), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n214), .B(new_n250), .C1(new_n253), .C2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G902), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n195), .A2(KEYINPUT7), .A3(new_n213), .A4(new_n209), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n258), .B(KEYINPUT80), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n238), .A2(new_n220), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n243), .B1(new_n228), .B2(new_n232), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n244), .ZN(new_n263));
  XOR2_X1   g077(.A(new_n246), .B(KEYINPUT8), .Z(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(KEYINPUT79), .A2(KEYINPUT7), .ZN(new_n266));
  NAND2_X1  g080(.A1(KEYINPUT79), .A2(KEYINPUT7), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n213), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n210), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n259), .A2(new_n265), .A3(new_n249), .A4(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n256), .A2(new_n257), .A3(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(G210), .B1(G237), .B2(G902), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n256), .A2(new_n257), .A3(new_n272), .A4(new_n270), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n188), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G952), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n277), .A2(KEYINPUT89), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n277), .A2(KEYINPUT89), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n212), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n280), .B1(G234), .B2(G237), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  XOR2_X1   g096(.A(KEYINPUT70), .B(G902), .Z(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  AOI211_X1 g098(.A(new_n212), .B(new_n284), .C1(G234), .C2(G237), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  XOR2_X1   g100(.A(KEYINPUT21), .B(G898), .Z(new_n287));
  OAI21_X1  g101(.A(new_n282), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n276), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G469), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n192), .B1(new_n189), .B2(new_n194), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n291), .B(new_n230), .C1(new_n231), .C2(new_n233), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n201), .A2(new_n207), .A3(new_n208), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(new_n240), .A3(new_n243), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT10), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT11), .ZN(new_n297));
  INV_X1    g111(.A(G134), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n297), .B1(new_n298), .B2(G137), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(G137), .ZN(new_n300));
  INV_X1    g114(.A(G137), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(KEYINPUT11), .A3(G134), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n299), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G131), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT64), .ZN(new_n305));
  INV_X1    g119(.A(G131), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n299), .A2(new_n302), .A3(new_n306), .A4(new_n300), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n304), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n303), .A2(KEYINPUT64), .A3(G131), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n293), .A2(new_n240), .A3(KEYINPUT10), .A4(new_n243), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n292), .A2(new_n296), .A3(new_n310), .A4(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(G110), .B(G140), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n212), .A2(G227), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n313), .B(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n261), .A2(new_n207), .A3(new_n208), .A4(new_n201), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n294), .ZN(new_n318));
  INV_X1    g132(.A(new_n310), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n318), .B(new_n319), .C1(KEYINPUT76), .C2(KEYINPUT12), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT12), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n308), .A2(KEYINPUT76), .A3(new_n309), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n261), .B(new_n293), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n321), .B(new_n322), .C1(new_n323), .C2(new_n310), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n316), .B1(new_n320), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n292), .A2(new_n296), .A3(new_n311), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n319), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n315), .B1(new_n327), .B2(new_n312), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n290), .B(new_n284), .C1(new_n325), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(G469), .A2(G902), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n327), .A2(new_n312), .A3(new_n315), .ZN(new_n331));
  INV_X1    g145(.A(new_n312), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n332), .B1(new_n320), .B2(new_n324), .ZN(new_n333));
  OAI211_X1 g147(.A(G469), .B(new_n331), .C1(new_n333), .C2(new_n315), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n329), .A2(new_n330), .A3(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT9), .B(G234), .ZN(new_n336));
  OAI21_X1  g150(.A(G221), .B1(new_n336), .B2(G902), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n289), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT20), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT85), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT84), .ZN(new_n342));
  INV_X1    g156(.A(G237), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(new_n212), .A3(G214), .ZN(new_n344));
  NOR2_X1   g158(.A1(KEYINPUT81), .A2(G143), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(G237), .A2(G953), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n347), .B(G214), .C1(KEYINPUT81), .C2(G143), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  AND4_X1   g163(.A1(new_n342), .A2(new_n349), .A3(KEYINPUT17), .A4(G131), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n306), .B1(new_n346), .B2(new_n348), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n342), .B1(new_n351), .B2(KEYINPUT17), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT16), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n203), .A2(new_n205), .A3(G140), .ZN(new_n355));
  NOR2_X1   g169(.A1(G125), .A2(G140), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n354), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  NOR3_X1   g172(.A1(new_n206), .A2(KEYINPUT16), .A3(G140), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n197), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G140), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n193), .A2(new_n354), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n356), .B1(new_n193), .B2(G140), .ZN(new_n363));
  OAI211_X1 g177(.A(G146), .B(new_n362), .C1(new_n363), .C2(new_n354), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n341), .B1(new_n353), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n349), .A2(KEYINPUT17), .A3(G131), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT84), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n351), .A2(new_n342), .A3(KEYINPUT17), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n370), .A2(KEYINPUT85), .A3(new_n360), .A4(new_n364), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n349), .A2(G131), .ZN(new_n372));
  OR3_X1    g186(.A1(new_n372), .A2(KEYINPUT17), .A3(new_n351), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n366), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(G113), .B(G122), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(new_n222), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n346), .A2(new_n348), .A3(KEYINPUT82), .ZN(new_n377));
  NAND2_X1  g191(.A1(KEYINPUT18), .A2(G131), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n377), .B(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(G125), .B(G140), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n197), .ZN(new_n381));
  INV_X1    g195(.A(new_n363), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n381), .B1(new_n382), .B2(new_n197), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n374), .A2(new_n376), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n376), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n372), .A2(new_n351), .ZN(new_n387));
  INV_X1    g201(.A(new_n364), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT19), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n380), .A2(new_n389), .ZN(new_n390));
  OR2_X1    g204(.A1(new_n390), .A2(KEYINPUT83), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(KEYINPUT83), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n363), .A2(KEYINPUT19), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  AOI211_X1 g208(.A(new_n387), .B(new_n388), .C1(new_n394), .C2(new_n197), .ZN(new_n395));
  INV_X1    g209(.A(new_n384), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n386), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n385), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g212(.A1(G475), .A2(G902), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n340), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n399), .ZN(new_n401));
  AOI211_X1 g215(.A(KEYINPUT20), .B(new_n401), .C1(new_n385), .C2(new_n397), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n374), .A2(new_n384), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n386), .ZN(new_n404));
  AOI21_X1  g218(.A(G902), .B1(new_n404), .B2(new_n385), .ZN(new_n405));
  INV_X1    g219(.A(G475), .ZN(new_n406));
  OAI22_X1  g220(.A1(new_n400), .A2(new_n402), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G478), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(KEYINPUT15), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT86), .B(KEYINPUT13), .ZN(new_n410));
  XNOR2_X1  g224(.A(G128), .B(G143), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n191), .A2(G143), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT13), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n414), .A2(KEYINPUT86), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n414), .A2(KEYINPUT86), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n413), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n412), .A2(new_n417), .A3(G134), .ZN(new_n418));
  INV_X1    g232(.A(G122), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G116), .ZN(new_n420));
  INV_X1    g234(.A(G116), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G122), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G107), .ZN(new_n424));
  XNOR2_X1  g238(.A(G116), .B(G122), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n225), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n411), .A2(new_n298), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n418), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n199), .A2(G128), .ZN(new_n430));
  OAI21_X1  g244(.A(G134), .B1(new_n413), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n426), .A2(KEYINPUT87), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n421), .A2(KEYINPUT14), .A3(G122), .ZN(new_n434));
  OAI211_X1 g248(.A(G107), .B(new_n434), .C1(new_n423), .C2(KEYINPUT14), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT87), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n425), .A2(new_n436), .A3(new_n225), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n432), .A2(new_n433), .A3(new_n435), .A4(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n429), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G217), .ZN(new_n440));
  NOR3_X1   g254(.A1(new_n336), .A2(new_n440), .A3(G953), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n429), .A2(new_n438), .A3(new_n441), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n284), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT88), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n409), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n446), .B(new_n447), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n448), .B1(new_n449), .B2(new_n409), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n407), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n339), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n221), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n301), .A2(G134), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n298), .A2(G137), .ZN(new_n456));
  OAI21_X1  g270(.A(G131), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n307), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT65), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT65), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n307), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n459), .A2(new_n293), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n308), .A2(new_n309), .A3(new_n291), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n454), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n458), .A2(KEYINPUT66), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT66), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n307), .A2(new_n457), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n465), .A2(new_n293), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT28), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n468), .A2(new_n463), .A3(new_n469), .A4(new_n454), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n463), .A3(new_n454), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT28), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n464), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(G101), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n347), .A2(G210), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n475), .B(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(KEYINPUT68), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT30), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n462), .A2(new_n463), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n480), .B1(new_n468), .B2(new_n463), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n221), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n471), .A2(new_n477), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT67), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT67), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n471), .A2(new_n486), .A3(new_n477), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT31), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n471), .A2(new_n486), .A3(new_n477), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n486), .B1(new_n471), .B2(new_n477), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n493), .A2(KEYINPUT31), .A3(new_n483), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n479), .B1(new_n490), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(G472), .A2(G902), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(KEYINPUT32), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n479), .ZN(new_n499));
  AOI21_X1  g313(.A(KEYINPUT31), .B1(new_n493), .B2(new_n483), .ZN(new_n500));
  AND4_X1   g314(.A1(KEYINPUT31), .A2(new_n483), .A3(new_n485), .A4(new_n487), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT32), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n503), .A3(new_n496), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n472), .A2(new_n470), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n468), .A2(new_n463), .ZN(new_n506));
  AOI21_X1  g320(.A(KEYINPUT69), .B1(new_n506), .B2(new_n221), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n468), .A2(new_n463), .A3(KEYINPUT69), .A4(new_n454), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(KEYINPUT29), .A3(new_n477), .ZN(new_n511));
  AOI21_X1  g325(.A(KEYINPUT29), .B1(new_n473), .B2(new_n478), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n483), .A2(new_n471), .ZN(new_n513));
  INV_X1    g327(.A(new_n477), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n511), .A2(new_n516), .A3(new_n284), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n498), .A2(new_n504), .B1(G472), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT71), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n519), .B1(new_n236), .B2(G128), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n236), .A2(G128), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n520), .A2(KEYINPUT23), .A3(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT23), .B1(new_n191), .B2(G119), .ZN(new_n523));
  AOI21_X1  g337(.A(KEYINPUT71), .B1(new_n191), .B2(G119), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(G110), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n522), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT73), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n522), .A2(new_n525), .A3(KEYINPUT73), .A4(new_n526), .ZN(new_n530));
  XNOR2_X1  g344(.A(G119), .B(G128), .ZN(new_n531));
  XOR2_X1   g345(.A(KEYINPUT24), .B(G110), .Z(new_n532));
  OAI211_X1 g346(.A(new_n529), .B(new_n530), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n533), .A2(new_n364), .A3(new_n381), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n526), .B1(new_n522), .B2(new_n525), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n535), .B1(new_n531), .B2(new_n532), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n365), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n212), .A2(G221), .A3(G234), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(KEYINPUT22), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(G137), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n534), .A2(new_n537), .A3(new_n541), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n284), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT25), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n440), .B1(new_n284), .B2(G234), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT25), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n543), .A2(new_n548), .A3(new_n284), .A4(new_n544), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n543), .A2(new_n544), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n547), .A2(G902), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT74), .B1(new_n518), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n517), .A2(G472), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n495), .A2(KEYINPUT32), .A3(new_n497), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n503), .B1(new_n502), .B2(new_n496), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT74), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n560), .A2(new_n561), .A3(new_n554), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n453), .B1(new_n556), .B2(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(new_n239), .ZN(G3));
  OAI21_X1  g378(.A(G472), .B1(new_n495), .B2(new_n283), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n502), .A2(new_n496), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n339), .A2(new_n554), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT33), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n445), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n283), .A2(new_n408), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n443), .A2(KEYINPUT90), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n429), .A2(new_n438), .A3(new_n441), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n441), .B1(new_n429), .B2(new_n438), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g389(.A(KEYINPUT33), .B(new_n572), .C1(new_n575), .C2(KEYINPUT90), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n576), .A2(KEYINPUT91), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT91), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT90), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n569), .B1(new_n445), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n578), .B1(new_n580), .B2(new_n572), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n570), .B(new_n571), .C1(new_n577), .C2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n446), .A2(new_n408), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n407), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n568), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT34), .B(G104), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(KEYINPUT92), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n586), .B(new_n588), .ZN(G6));
  INV_X1    g403(.A(new_n385), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n376), .B1(new_n374), .B2(new_n384), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n257), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(G475), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n398), .A2(new_n399), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(KEYINPUT20), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n398), .A2(new_n340), .A3(new_n399), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(KEYINPUT93), .A3(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT93), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n599), .B1(new_n400), .B2(new_n402), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n594), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n451), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n568), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT35), .B(G107), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G9));
  NOR2_X1   g419(.A1(new_n542), .A2(KEYINPUT36), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n538), .B(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n552), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n550), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n565), .A2(new_n566), .A3(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT94), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n453), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(KEYINPUT37), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G110), .ZN(G12));
  AOI21_X1  g430(.A(new_n338), .B1(new_n550), .B2(new_n608), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n560), .A2(new_n276), .A3(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n282), .B1(new_n286), .B2(G900), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n601), .A2(new_n451), .A3(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT95), .B(G128), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G30));
  INV_X1    g437(.A(new_n338), .ZN(new_n624));
  XOR2_X1   g438(.A(new_n619), .B(KEYINPUT96), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(KEYINPUT39), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT97), .B(KEYINPUT40), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n498), .A2(new_n504), .ZN(new_n630));
  INV_X1    g444(.A(new_n478), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n507), .A2(new_n471), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n631), .A2(new_n509), .A3(new_n632), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n633), .A2(new_n488), .ZN(new_n634));
  OAI21_X1  g448(.A(G472), .B1(new_n634), .B2(G902), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n609), .B1(new_n630), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n274), .A2(new_n275), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT38), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n274), .A2(KEYINPUT38), .A3(new_n275), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n407), .A2(new_n451), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n641), .A2(new_n642), .A3(new_n188), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n629), .A2(new_n636), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G143), .ZN(G45));
  NAND3_X1  g459(.A1(new_n407), .A2(new_n584), .A3(new_n619), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n618), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(new_n197), .ZN(G48));
  NAND2_X1  g462(.A1(new_n560), .A2(new_n554), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n284), .B1(new_n325), .B2(new_n328), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(G469), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n651), .A2(new_n337), .A3(new_n329), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  OR4_X1    g467(.A1(new_n649), .A2(new_n653), .A3(new_n289), .A4(new_n585), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT41), .B(G113), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT98), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n654), .B(new_n656), .ZN(G15));
  NOR4_X1   g471(.A1(new_n649), .A2(new_n602), .A3(new_n653), .A4(new_n289), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(new_n421), .ZN(G18));
  AND2_X1   g473(.A1(new_n452), .A2(new_n288), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n276), .A2(new_n652), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n660), .A2(new_n560), .A3(new_n609), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT99), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G119), .ZN(G21));
  INV_X1    g478(.A(new_n276), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n642), .A2(new_n665), .A3(new_n653), .ZN(new_n666));
  OAI22_X1  g480(.A1(new_n500), .A2(new_n501), .B1(new_n478), .B2(new_n510), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n496), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n565), .A2(new_n554), .A3(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n666), .A2(new_n288), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G122), .ZN(G24));
  AND3_X1   g486(.A1(new_n565), .A2(new_n609), .A3(new_n668), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n407), .A2(new_n584), .A3(new_n619), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n673), .A2(new_n674), .A3(new_n661), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(KEYINPUT100), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n565), .A2(new_n609), .A3(new_n668), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n677), .A2(new_n646), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT100), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n678), .A2(new_n679), .A3(new_n661), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G125), .ZN(G27));
  INV_X1    g496(.A(new_n337), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT101), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n335), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n329), .A2(new_n334), .A3(KEYINPUT101), .A4(new_n330), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n683), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n274), .A2(new_n187), .A3(new_n275), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT102), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n274), .A2(KEYINPUT102), .A3(new_n187), .A4(new_n275), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(KEYINPUT103), .B1(new_n688), .B2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT103), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n687), .A2(new_n691), .A3(new_n695), .A4(new_n692), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n649), .ZN(new_n698));
  AND4_X1   g512(.A1(KEYINPUT42), .A2(new_n697), .A3(new_n698), .A4(new_n674), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n649), .B1(new_n694), .B2(new_n696), .ZN(new_n700));
  AOI21_X1  g514(.A(KEYINPUT42), .B1(new_n700), .B2(new_n674), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT104), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G131), .ZN(G33));
  AND3_X1   g518(.A1(new_n601), .A2(new_n451), .A3(new_n619), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n700), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G134), .ZN(G36));
  INV_X1    g521(.A(KEYINPUT43), .ZN(new_n708));
  INV_X1    g522(.A(new_n583), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n576), .A2(KEYINPUT91), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n580), .A2(new_n578), .A3(new_n572), .ZN(new_n711));
  AOI22_X1  g525(.A1(new_n710), .A2(new_n711), .B1(new_n569), .B2(new_n445), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n709), .B1(new_n712), .B2(new_n571), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n708), .B1(new_n407), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n596), .A2(new_n597), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n715), .A2(new_n584), .A3(KEYINPUT43), .A4(new_n593), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  OR2_X1    g531(.A1(new_n717), .A2(KEYINPUT105), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n567), .B1(new_n717), .B2(KEYINPUT105), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(new_n609), .A3(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n693), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n324), .A2(new_n320), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n315), .B1(new_n724), .B2(new_n312), .ZN(new_n725));
  INV_X1    g539(.A(new_n331), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n723), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI211_X1 g541(.A(KEYINPUT45), .B(new_n331), .C1(new_n333), .C2(new_n315), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(G469), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(KEYINPUT46), .B1(new_n729), .B2(new_n330), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n729), .A2(KEYINPUT46), .A3(new_n330), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n731), .A2(new_n329), .A3(new_n732), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n733), .A2(new_n337), .A3(new_n626), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n722), .B(new_n734), .C1(new_n721), .C2(new_n720), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(KEYINPUT106), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G137), .ZN(G39));
  INV_X1    g551(.A(KEYINPUT47), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n729), .A2(KEYINPUT46), .A3(new_n330), .ZN(new_n739));
  INV_X1    g553(.A(new_n329), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n739), .A2(new_n730), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n738), .B1(new_n741), .B2(new_n683), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n733), .A2(KEYINPUT47), .A3(new_n337), .ZN(new_n743));
  AOI211_X1 g557(.A(new_n560), .B(new_n646), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n691), .A2(new_n692), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n744), .A2(new_n555), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G140), .ZN(G42));
  INV_X1    g561(.A(new_n651), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n748), .A2(new_n740), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n749), .A2(KEYINPUT111), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(KEYINPUT111), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(new_n683), .A3(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n742), .A2(new_n743), .A3(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n282), .B1(new_n714), .B2(new_n716), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT110), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n756), .A2(new_n757), .A3(new_n670), .A4(new_n745), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n717), .A2(new_n745), .A3(new_n281), .A4(new_n670), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT110), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n742), .A2(new_n743), .A3(KEYINPUT114), .A4(new_n752), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n755), .A2(new_n758), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n745), .A2(new_n554), .A3(new_n652), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n630), .A2(new_n281), .A3(new_n635), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n715), .A2(new_n713), .A3(new_n593), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  AOI211_X1 g580(.A(new_n282), .B(new_n669), .C1(new_n714), .C2(new_n716), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT113), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n641), .A2(new_n768), .A3(new_n188), .A4(new_n652), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n274), .A2(KEYINPUT38), .A3(new_n275), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT38), .B1(new_n274), .B2(new_n275), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n188), .B(new_n652), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(KEYINPUT113), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n767), .A2(KEYINPUT50), .A3(new_n769), .A4(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT50), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n773), .A2(new_n769), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n717), .A2(new_n281), .A3(new_n670), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n766), .B1(new_n774), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n693), .A2(new_n653), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n756), .A2(new_n780), .A3(new_n673), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n762), .A2(KEYINPUT51), .A3(new_n779), .A4(new_n781), .ZN(new_n782));
  OR3_X1    g596(.A1(new_n763), .A2(new_n585), .A3(new_n764), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n698), .A2(new_n756), .A3(new_n780), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n784), .A2(KEYINPUT48), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(KEYINPUT48), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n280), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n782), .A2(new_n783), .A3(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n753), .A2(new_n760), .A3(new_n758), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(KEYINPUT112), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n753), .A2(new_n760), .A3(new_n791), .A4(new_n758), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n790), .A2(new_n779), .A3(new_n781), .A4(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT51), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n767), .A2(new_n661), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n788), .A2(KEYINPUT115), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n782), .A2(new_n796), .A3(new_n783), .A4(new_n787), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n793), .A2(new_n794), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n803));
  INV_X1    g617(.A(new_n662), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n658), .A2(new_n804), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n805), .A2(new_n654), .A3(new_n671), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n618), .B1(new_n620), .B2(new_n646), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n807), .B1(new_n680), .B2(new_n676), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n407), .A2(new_n276), .A3(new_n451), .ZN(new_n809));
  XOR2_X1   g623(.A(new_n619), .B(KEYINPUT107), .Z(new_n810));
  NAND4_X1  g624(.A1(new_n636), .A2(new_n687), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT108), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n688), .A2(new_n665), .A3(new_n642), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n814), .A2(KEYINPUT108), .A3(new_n636), .A4(new_n810), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT52), .B1(new_n808), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n624), .A2(new_n609), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n518), .A2(new_n818), .A3(new_n665), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n819), .B1(new_n705), .B2(new_n674), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n681), .A2(new_n813), .A3(new_n815), .A4(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT52), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n806), .B1(new_n817), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n700), .A2(new_n674), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT42), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n700), .A2(KEYINPUT42), .A3(new_n674), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n691), .A2(new_n619), .A3(new_n692), .ZN(new_n830));
  NOR4_X1   g644(.A1(new_n830), .A2(new_n518), .A3(new_n818), .A4(new_n451), .ZN(new_n831));
  AOI22_X1  g645(.A1(new_n700), .A2(new_n705), .B1(new_n831), .B2(new_n601), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n697), .A2(new_n678), .ZN(new_n833));
  INV_X1    g647(.A(new_n585), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n407), .A2(new_n450), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n568), .A2(new_n836), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n563), .A2(new_n614), .A3(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n829), .A2(new_n832), .A3(new_n833), .A4(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n803), .B1(new_n824), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n805), .A2(new_n654), .A3(new_n671), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n808), .A2(new_n816), .A3(KEYINPUT52), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n821), .A2(new_n822), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n838), .A2(new_n832), .A3(new_n833), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n845), .A2(new_n702), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n844), .A2(new_n846), .A3(KEYINPUT53), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n840), .A2(KEYINPUT109), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT109), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n844), .A2(new_n846), .A3(new_n849), .A4(KEYINPUT53), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n848), .A2(KEYINPUT54), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n840), .A2(new_n852), .A3(new_n847), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n802), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n277), .A2(new_n212), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n749), .B(KEYINPUT49), .ZN(new_n857));
  AND4_X1   g671(.A1(new_n554), .A2(new_n857), .A3(new_n337), .A4(new_n641), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n630), .A2(new_n635), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n407), .A2(new_n713), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n858), .A2(new_n187), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n856), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT116), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n856), .A2(KEYINPUT116), .A3(new_n861), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(G75));
  OAI21_X1  g680(.A(new_n250), .B1(new_n253), .B2(new_n255), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(new_n214), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n868), .B(KEYINPUT55), .Z(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  AOI211_X1 g684(.A(new_n284), .B(new_n272), .C1(new_n840), .C2(new_n847), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT56), .B1(new_n871), .B2(KEYINPUT117), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n844), .A2(new_n846), .A3(KEYINPUT53), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT53), .B1(new_n844), .B2(new_n846), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n283), .B(new_n273), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT117), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n870), .B1(new_n872), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n212), .A2(G952), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(KEYINPUT120), .Z(new_n880));
  INV_X1    g694(.A(KEYINPUT56), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n881), .B1(new_n869), .B2(KEYINPUT118), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n882), .B1(KEYINPUT118), .B2(new_n869), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n875), .A2(KEYINPUT119), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT119), .B1(new_n875), .B2(new_n883), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n880), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(KEYINPUT121), .B1(new_n878), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n877), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n881), .B1(new_n875), .B2(new_n876), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n869), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n885), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n875), .A2(KEYINPUT119), .A3(new_n883), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n890), .A2(new_n893), .A3(new_n894), .A4(new_n880), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n887), .A2(new_n895), .ZN(G51));
  NAND2_X1  g710(.A1(new_n840), .A2(new_n847), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT54), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n853), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n330), .A2(KEYINPUT57), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n330), .A2(KEYINPUT57), .ZN(new_n902));
  OAI22_X1  g716(.A1(new_n901), .A2(new_n902), .B1(new_n328), .B2(new_n325), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n897), .A2(new_n283), .ZN(new_n904));
  OR2_X1    g718(.A1(new_n904), .A2(new_n729), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n879), .B1(new_n903), .B2(new_n905), .ZN(G54));
  NAND4_X1  g720(.A1(new_n897), .A2(KEYINPUT58), .A3(G475), .A4(new_n283), .ZN(new_n907));
  INV_X1    g721(.A(new_n398), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n907), .A2(new_n908), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n909), .A2(new_n910), .A3(new_n879), .ZN(G60));
  NAND2_X1  g725(.A1(G478), .A2(G902), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT59), .Z(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n899), .A2(new_n712), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n913), .B1(new_n851), .B2(new_n853), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n915), .B(new_n880), .C1(new_n916), .C2(new_n712), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(G63));
  XNOR2_X1  g732(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n440), .A2(new_n257), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n919), .B(new_n920), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n607), .B(KEYINPUT123), .Z(new_n922));
  NAND3_X1  g736(.A1(new_n897), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n897), .A2(new_n921), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n880), .B(new_n923), .C1(new_n924), .C2(new_n551), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT61), .Z(G66));
  NAND2_X1  g740(.A1(new_n287), .A2(new_n211), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(G953), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n806), .A2(new_n838), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n928), .B1(new_n930), .B2(G953), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n867), .B1(G898), .B2(new_n212), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(G69));
  OR2_X1    g747(.A1(new_n481), .A2(new_n482), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(new_n394), .Z(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT124), .Z(new_n936));
  NAND2_X1  g750(.A1(new_n808), .A2(new_n644), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT62), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n937), .A2(KEYINPUT125), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(KEYINPUT125), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n808), .A2(new_n644), .A3(new_n940), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  OR2_X1    g756(.A1(new_n938), .A2(KEYINPUT125), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n627), .B1(new_n556), .B2(new_n562), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n944), .B(new_n745), .C1(new_n834), .C2(new_n835), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n735), .A2(new_n746), .A3(new_n943), .A4(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n942), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n936), .B1(new_n947), .B2(G953), .ZN(new_n948));
  NAND2_X1  g762(.A1(G900), .A2(G953), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n735), .A2(new_n746), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n734), .A2(new_n698), .A3(new_n809), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n829), .A2(new_n706), .A3(new_n808), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n949), .B1(new_n953), .B2(G953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n948), .B1(new_n954), .B2(new_n935), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n212), .B1(G227), .B2(G900), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(G72));
  NAND2_X1  g771(.A1(G472), .A2(G902), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT63), .Z(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n947), .B2(new_n930), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n513), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n939), .A2(new_n941), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n950), .A2(new_n943), .A3(new_n945), .A4(new_n964), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n962), .B(new_n959), .C1(new_n965), .C2(new_n929), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n477), .ZN(new_n967));
  OAI21_X1  g781(.A(KEYINPUT127), .B1(new_n963), .B2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n513), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n959), .B1(new_n965), .B2(new_n929), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n969), .B1(new_n970), .B2(KEYINPUT126), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT127), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n971), .A2(new_n972), .A3(new_n477), .A4(new_n966), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n968), .A2(new_n973), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n848), .A2(new_n850), .A3(new_n959), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n515), .A2(new_n488), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n879), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n959), .B1(new_n953), .B2(new_n929), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n978), .A2(new_n514), .A3(new_n969), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n974), .A2(new_n977), .A3(new_n979), .ZN(G57));
endmodule


