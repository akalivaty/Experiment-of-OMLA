

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n720, n721, n722, n723, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756;

  XNOR2_X1 U363 ( .A(n723), .B(n344), .ZN(G75) );
  NOR2_X1 U364 ( .A1(G953), .A2(n722), .ZN(n723) );
  XNOR2_X1 U365 ( .A(n345), .B(KEYINPUT121), .ZN(n344) );
  INV_X1 U366 ( .A(KEYINPUT53), .ZN(n345) );
  NAND2_X1 U367 ( .A1(n342), .A2(n718), .ZN(n720) );
  XNOR2_X1 U368 ( .A(n714), .B(n343), .ZN(n342) );
  INV_X1 U369 ( .A(KEYINPUT2), .ZN(n343) );
  AND2_X1 U370 ( .A1(n348), .A2(n380), .ZN(n368) );
  NOR2_X1 U371 ( .A1(n566), .A2(n625), .ZN(n578) );
  AND2_X1 U372 ( .A1(n390), .A2(n574), .ZN(n348) );
  BUF_X1 U373 ( .A(n569), .Z(n625) );
  XNOR2_X1 U374 ( .A(n413), .B(KEYINPUT33), .ZN(n692) );
  NAND2_X1 U375 ( .A1(n570), .A2(n609), .ZN(n413) );
  OR2_X2 U376 ( .A1(n651), .A2(G902), .ZN(n388) );
  NOR2_X1 U377 ( .A1(G953), .A2(G237), .ZN(n532) );
  XNOR2_X1 U378 ( .A(G116), .B(G122), .ZN(n514) );
  NAND2_X1 U379 ( .A1(n475), .A2(n474), .ZN(n500) );
  XNOR2_X1 U380 ( .A(n405), .B(n404), .ZN(n566) );
  INV_X1 U381 ( .A(G953), .ZN(n739) );
  BUF_X1 U382 ( .A(G143), .Z(n415) );
  XNOR2_X2 U383 ( .A(n542), .B(n444), .ZN(n443) );
  AND2_X1 U384 ( .A1(n632), .A2(n631), .ZN(n416) );
  NOR2_X1 U385 ( .A1(n752), .A2(n756), .ZN(n450) );
  INV_X1 U386 ( .A(n676), .ZN(n419) );
  INV_X1 U387 ( .A(n601), .ZN(n374) );
  INV_X1 U388 ( .A(KEYINPUT22), .ZN(n404) );
  INV_X1 U389 ( .A(KEYINPUT3), .ZN(n446) );
  AND2_X1 U390 ( .A1(n402), .A2(n398), .ZN(n396) );
  AND2_X1 U391 ( .A1(n432), .A2(n754), .ZN(n431) );
  NOR2_X1 U392 ( .A1(n562), .A2(n561), .ZN(n663) );
  XNOR2_X1 U393 ( .A(n567), .B(n436), .ZN(n568) );
  XNOR2_X1 U394 ( .A(n422), .B(n420), .ZN(n756) );
  XNOR2_X1 U395 ( .A(n440), .B(n439), .ZN(n601) );
  XNOR2_X1 U396 ( .A(n446), .B(G119), .ZN(n464) );
  INV_X1 U397 ( .A(n554), .ZN(n444) );
  XNOR2_X2 U398 ( .A(G110), .B(KEYINPUT88), .ZN(n466) );
  XNOR2_X1 U399 ( .A(n635), .B(KEYINPUT65), .ZN(n346) );
  XNOR2_X1 U400 ( .A(n635), .B(KEYINPUT65), .ZN(n347) );
  XNOR2_X1 U401 ( .A(n635), .B(KEYINPUT65), .ZN(n725) );
  NAND2_X2 U402 ( .A1(n634), .A2(n633), .ZN(n635) );
  OR2_X1 U403 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U404 ( .A(n424), .B(n615), .ZN(n752) );
  AND2_X1 U405 ( .A1(n576), .A2(n642), .ZN(n435) );
  OR2_X1 U406 ( .A1(n581), .A2(n571), .ZN(n390) );
  NAND2_X1 U407 ( .A1(n715), .A2(n416), .ZN(n713) );
  NOR2_X1 U408 ( .A1(n608), .A2(KEYINPUT67), .ZN(n384) );
  XNOR2_X1 U409 ( .A(n451), .B(KEYINPUT101), .ZN(n616) );
  OR2_X1 U410 ( .A1(n585), .A2(n523), .ZN(n451) );
  NAND2_X1 U411 ( .A1(n364), .A2(n350), .ZN(n429) );
  NOR2_X1 U412 ( .A1(n385), .A2(n383), .ZN(n382) );
  NAND2_X1 U413 ( .A1(n641), .A2(n442), .ZN(n385) );
  XNOR2_X1 U414 ( .A(n384), .B(n441), .ZN(n383) );
  NOR2_X1 U415 ( .A1(G902), .A2(G237), .ZN(n487) );
  XNOR2_X1 U416 ( .A(G131), .B(n415), .ZN(n494) );
  XNOR2_X1 U417 ( .A(KEYINPUT70), .B(G137), .ZN(n554) );
  XNOR2_X1 U418 ( .A(n587), .B(n358), .ZN(n715) );
  NOR2_X1 U419 ( .A1(n699), .A2(n697), .ZN(n619) );
  XNOR2_X1 U420 ( .A(n603), .B(KEYINPUT1), .ZN(n569) );
  XNOR2_X1 U421 ( .A(n538), .B(n537), .ZN(n541) );
  XOR2_X1 U422 ( .A(KEYINPUT69), .B(KEYINPUT10), .Z(n502) );
  NAND2_X1 U423 ( .A1(n353), .A2(n376), .ZN(n624) );
  NOR2_X1 U424 ( .A1(n610), .A2(n454), .ZN(n376) );
  AND2_X1 U425 ( .A1(n379), .A2(n348), .ZN(n370) );
  INV_X1 U426 ( .A(n575), .ZN(n378) );
  INV_X1 U427 ( .A(n628), .ZN(n411) );
  NAND2_X1 U428 ( .A1(n621), .A2(n386), .ZN(n606) );
  AND2_X1 U429 ( .A1(n387), .A2(n620), .ZN(n386) );
  XNOR2_X1 U430 ( .A(n509), .B(n508), .ZN(n585) );
  XNOR2_X1 U431 ( .A(n572), .B(n409), .ZN(n584) );
  INV_X1 U432 ( .A(G478), .ZN(n409) );
  INV_X1 U433 ( .A(KEYINPUT32), .ZN(n436) );
  INV_X1 U434 ( .A(n700), .ZN(n433) );
  INV_X1 U435 ( .A(KEYINPUT47), .ZN(n441) );
  XNOR2_X1 U436 ( .A(n453), .B(n452), .ZN(n699) );
  INV_X1 U437 ( .A(KEYINPUT109), .ZN(n452) );
  OR2_X1 U438 ( .A1(n617), .A2(n454), .ZN(n453) );
  INV_X1 U439 ( .A(KEYINPUT92), .ZN(n535) );
  XNOR2_X1 U440 ( .A(G137), .B(G146), .ZN(n536) );
  INV_X1 U441 ( .A(KEYINPUT71), .ZN(n449) );
  INV_X1 U442 ( .A(KEYINPUT48), .ZN(n447) );
  XNOR2_X1 U443 ( .A(KEYINPUT87), .B(KEYINPUT15), .ZN(n455) );
  INV_X1 U444 ( .A(KEYINPUT17), .ZN(n479) );
  NAND2_X1 U445 ( .A1(G234), .A2(G237), .ZN(n458) );
  INV_X1 U446 ( .A(KEYINPUT76), .ZN(n445) );
  XNOR2_X1 U447 ( .A(n491), .B(n490), .ZN(n604) );
  INV_X1 U448 ( .A(KEYINPUT19), .ZN(n490) );
  XNOR2_X1 U449 ( .A(n522), .B(n521), .ZN(n572) );
  XOR2_X1 U450 ( .A(KEYINPUT73), .B(KEYINPUT23), .Z(n548) );
  XNOR2_X1 U451 ( .A(G119), .B(G128), .ZN(n551) );
  INV_X1 U452 ( .A(G128), .ZN(n469) );
  XNOR2_X1 U453 ( .A(G134), .B(G107), .ZN(n515) );
  XNOR2_X1 U454 ( .A(n406), .B(n744), .ZN(n636) );
  XNOR2_X1 U455 ( .A(n506), .B(n505), .ZN(n406) );
  NOR2_X1 U456 ( .A1(n613), .A2(n617), .ZN(n614) );
  INV_X1 U457 ( .A(G472), .ZN(n439) );
  AND2_X1 U458 ( .A1(n603), .A2(n417), .ZN(n588) );
  XNOR2_X1 U459 ( .A(n580), .B(n392), .ZN(n581) );
  INV_X1 U460 ( .A(n747), .ZN(n372) );
  XNOR2_X1 U461 ( .A(n443), .B(n352), .ZN(n651) );
  XNOR2_X1 U462 ( .A(G146), .B(G140), .ZN(n527) );
  NAND2_X1 U463 ( .A1(n716), .A2(n373), .ZN(n717) );
  XNOR2_X1 U464 ( .A(n622), .B(n421), .ZN(n420) );
  NAND2_X1 U465 ( .A1(n423), .A2(n354), .ZN(n422) );
  INV_X1 U466 ( .A(KEYINPUT111), .ZN(n421) );
  XNOR2_X1 U467 ( .A(n375), .B(KEYINPUT36), .ZN(n611) );
  NOR2_X1 U468 ( .A1(n624), .A2(n628), .ZN(n375) );
  NAND2_X1 U469 ( .A1(n377), .A2(n370), .ZN(n369) );
  XNOR2_X1 U470 ( .A(n365), .B(n414), .ZN(n671) );
  INV_X1 U471 ( .A(KEYINPUT31), .ZN(n414) );
  NOR2_X1 U472 ( .A1(n687), .A2(n580), .ZN(n365) );
  NOR2_X1 U473 ( .A1(n606), .A2(n605), .ZN(n667) );
  AND2_X1 U474 ( .A1(n597), .A2(n411), .ZN(n410) );
  NOR2_X1 U475 ( .A1(n607), .A2(n606), .ZN(n664) );
  INV_X1 U476 ( .A(n605), .ZN(n668) );
  XNOR2_X1 U477 ( .A(n568), .B(G119), .ZN(n755) );
  INV_X1 U478 ( .A(n677), .ZN(n418) );
  XOR2_X1 U479 ( .A(n546), .B(KEYINPUT25), .Z(n349) );
  OR2_X1 U480 ( .A1(n433), .A2(n430), .ZN(n350) );
  AND2_X1 U481 ( .A1(n433), .A2(n430), .ZN(n351) );
  XOR2_X1 U482 ( .A(n530), .B(n529), .Z(n352) );
  AND2_X1 U483 ( .A1(n609), .A2(n668), .ZN(n353) );
  AND2_X1 U484 ( .A1(n621), .A2(n620), .ZN(n354) );
  AND2_X1 U485 ( .A1(n659), .A2(n351), .ZN(n355) );
  NAND2_X1 U486 ( .A1(n419), .A2(n418), .ZN(n681) );
  AND2_X1 U487 ( .A1(n489), .A2(G210), .ZN(n356) );
  NOR2_X1 U488 ( .A1(n685), .A2(n374), .ZN(n357) );
  XOR2_X1 U489 ( .A(n586), .B(KEYINPUT64), .Z(n358) );
  XOR2_X1 U490 ( .A(n651), .B(n650), .Z(n359) );
  XOR2_X1 U491 ( .A(n655), .B(n654), .Z(n360) );
  XOR2_X1 U492 ( .A(n648), .B(KEYINPUT123), .Z(n361) );
  XNOR2_X1 U493 ( .A(KEYINPUT62), .B(n645), .ZN(n362) );
  XNOR2_X1 U494 ( .A(n636), .B(KEYINPUT59), .ZN(n363) );
  INV_X1 U495 ( .A(n730), .ZN(n398) );
  NAND2_X1 U496 ( .A1(n671), .A2(n351), .ZN(n364) );
  XNOR2_X2 U497 ( .A(n366), .B(n445), .ZN(n570) );
  NAND2_X1 U498 ( .A1(n569), .A2(n417), .ZN(n366) );
  XNOR2_X2 U499 ( .A(n388), .B(n531), .ZN(n603) );
  NAND2_X1 U500 ( .A1(n367), .A2(n575), .ZN(n371) );
  NAND2_X1 U501 ( .A1(n368), .A2(n379), .ZN(n367) );
  NAND2_X1 U502 ( .A1(n371), .A2(n369), .ZN(n642) );
  XNOR2_X1 U503 ( .A(n416), .B(n372), .ZN(n745) );
  INV_X1 U504 ( .A(n416), .ZN(n373) );
  NAND2_X1 U505 ( .A1(n374), .A2(n693), .ZN(n593) );
  XNOR2_X1 U506 ( .A(n601), .B(KEYINPUT6), .ZN(n609) );
  NOR2_X2 U507 ( .A1(n583), .A2(n374), .ZN(n659) );
  AND2_X1 U508 ( .A1(n380), .A2(n378), .ZN(n377) );
  NAND2_X1 U509 ( .A1(n381), .A2(n389), .ZN(n379) );
  NAND2_X1 U510 ( .A1(n391), .A2(n692), .ZN(n380) );
  INV_X1 U511 ( .A(n692), .ZN(n381) );
  XNOR2_X1 U512 ( .A(n382), .B(n449), .ZN(n408) );
  NAND2_X1 U513 ( .A1(n611), .A2(n625), .ZN(n641) );
  INV_X1 U514 ( .A(n604), .ZN(n387) );
  INV_X1 U515 ( .A(n571), .ZN(n389) );
  AND2_X1 U516 ( .A1(n581), .A2(n571), .ZN(n391) );
  INV_X1 U517 ( .A(KEYINPUT90), .ZN(n392) );
  XNOR2_X1 U518 ( .A(n393), .B(KEYINPUT124), .ZN(G63) );
  AND2_X2 U519 ( .A1(n399), .A2(n398), .ZN(n393) );
  XNOR2_X1 U520 ( .A(n394), .B(KEYINPUT56), .ZN(G51) );
  AND2_X2 U521 ( .A1(n400), .A2(n398), .ZN(n394) );
  XNOR2_X1 U522 ( .A(n395), .B(n639), .ZN(G60) );
  AND2_X2 U523 ( .A1(n401), .A2(n398), .ZN(n395) );
  XNOR2_X1 U524 ( .A(n396), .B(n647), .ZN(G57) );
  XNOR2_X1 U525 ( .A(n397), .B(KEYINPUT122), .ZN(G54) );
  AND2_X2 U526 ( .A1(n403), .A2(n398), .ZN(n397) );
  XNOR2_X1 U527 ( .A(n649), .B(n361), .ZN(n399) );
  XNOR2_X1 U528 ( .A(n656), .B(n360), .ZN(n400) );
  XNOR2_X1 U529 ( .A(n637), .B(n363), .ZN(n401) );
  XNOR2_X1 U530 ( .A(n646), .B(n362), .ZN(n402) );
  XNOR2_X1 U531 ( .A(n652), .B(n359), .ZN(n403) );
  NOR2_X2 U532 ( .A1(n438), .A2(n580), .ZN(n405) );
  BUF_X1 U533 ( .A(n603), .Z(n620) );
  NAND2_X1 U534 ( .A1(n407), .A2(n408), .ZN(n448) );
  XNOR2_X1 U535 ( .A(n450), .B(KEYINPUT46), .ZN(n407) );
  INV_X1 U536 ( .A(n753), .ZN(n442) );
  NAND2_X1 U537 ( .A1(n412), .A2(n410), .ZN(n598) );
  INV_X1 U538 ( .A(n613), .ZN(n412) );
  NAND2_X1 U539 ( .A1(n645), .A2(n544), .ZN(n440) );
  XNOR2_X1 U540 ( .A(n448), .B(n447), .ZN(n632) );
  XNOR2_X1 U541 ( .A(n435), .B(KEYINPUT44), .ZN(n434) );
  INV_X1 U542 ( .A(n681), .ZN(n417) );
  XNOR2_X2 U543 ( .A(n560), .B(n349), .ZN(n676) );
  INV_X1 U544 ( .A(n675), .ZN(n423) );
  NAND2_X1 U545 ( .A1(n623), .A2(n668), .ZN(n424) );
  XNOR2_X1 U546 ( .A(n614), .B(n425), .ZN(n623) );
  INV_X1 U547 ( .A(KEYINPUT39), .ZN(n425) );
  NAND2_X1 U548 ( .A1(n428), .A2(n426), .ZN(n432) );
  OR2_X1 U549 ( .A1(n659), .A2(n427), .ZN(n426) );
  OR2_X1 U550 ( .A1(n671), .A2(n430), .ZN(n427) );
  NOR2_X1 U551 ( .A1(n355), .A2(n429), .ZN(n428) );
  INV_X1 U552 ( .A(KEYINPUT100), .ZN(n430) );
  NAND2_X1 U553 ( .A1(n431), .A2(n434), .ZN(n587) );
  XNOR2_X2 U554 ( .A(n437), .B(n493), .ZN(n580) );
  NOR2_X2 U555 ( .A1(n604), .A2(n492), .ZN(n437) );
  NAND2_X1 U556 ( .A1(n616), .A2(n418), .ZN(n438) );
  NOR2_X1 U557 ( .A1(n663), .A2(n568), .ZN(n576) );
  XNOR2_X1 U558 ( .A(n542), .B(n543), .ZN(n645) );
  XNOR2_X1 U559 ( .A(n443), .B(n744), .ZN(n747) );
  NAND2_X1 U560 ( .A1(n570), .A2(n374), .ZN(n687) );
  INV_X1 U561 ( .A(n617), .ZN(n694) );
  INV_X1 U562 ( .A(n616), .ZN(n697) );
  INV_X1 U563 ( .A(n693), .ZN(n454) );
  BUF_X1 U564 ( .A(n653), .Z(n655) );
  NAND2_X1 U565 ( .A1(n612), .A2(n693), .ZN(n491) );
  XNOR2_X1 U566 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U567 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U568 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U569 ( .A(n507), .B(G475), .ZN(n508) );
  INV_X1 U570 ( .A(KEYINPUT42), .ZN(n622) );
  BUF_X1 U571 ( .A(n642), .Z(n644) );
  INV_X1 U572 ( .A(G902), .ZN(n544) );
  XNOR2_X1 U573 ( .A(n455), .B(n544), .ZN(n486) );
  NAND2_X1 U574 ( .A1(G234), .A2(n486), .ZN(n456) );
  XNOR2_X1 U575 ( .A(KEYINPUT20), .B(n456), .ZN(n545) );
  NAND2_X1 U576 ( .A1(n545), .A2(G221), .ZN(n457) );
  XNOR2_X1 U577 ( .A(n457), .B(KEYINPUT21), .ZN(n677) );
  INV_X1 U578 ( .A(KEYINPUT0), .ZN(n493) );
  XNOR2_X1 U579 ( .A(n458), .B(KEYINPUT14), .ZN(n461) );
  NAND2_X1 U580 ( .A1(G952), .A2(n461), .ZN(n709) );
  NOR2_X1 U581 ( .A1(G953), .A2(n709), .ZN(n459) );
  XOR2_X1 U582 ( .A(KEYINPUT89), .B(n459), .Z(n592) );
  AND2_X1 U583 ( .A1(G953), .A2(G902), .ZN(n460) );
  NAND2_X1 U584 ( .A1(n461), .A2(n460), .ZN(n589) );
  NOR2_X1 U585 ( .A1(G898), .A2(n589), .ZN(n462) );
  NOR2_X1 U586 ( .A1(n592), .A2(n462), .ZN(n492) );
  XOR2_X2 U587 ( .A(G122), .B(G104), .Z(n504) );
  XNOR2_X1 U588 ( .A(n504), .B(KEYINPUT16), .ZN(n465) );
  XNOR2_X1 U589 ( .A(G113), .B(G116), .ZN(n463) );
  XNOR2_X1 U590 ( .A(n464), .B(n463), .ZN(n539) );
  XNOR2_X1 U591 ( .A(n465), .B(n539), .ZN(n737) );
  INV_X1 U592 ( .A(n466), .ZN(n468) );
  XNOR2_X1 U593 ( .A(G101), .B(G107), .ZN(n467) );
  XNOR2_X1 U594 ( .A(n468), .B(n467), .ZN(n735) );
  XNOR2_X1 U595 ( .A(n735), .B(KEYINPUT74), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n737), .B(n530), .ZN(n485) );
  XNOR2_X2 U597 ( .A(KEYINPUT81), .B(G143), .ZN(n470) );
  XNOR2_X2 U598 ( .A(n470), .B(n469), .ZN(n512) );
  XNOR2_X2 U599 ( .A(n512), .B(KEYINPUT4), .ZN(n525) );
  INV_X1 U600 ( .A(G146), .ZN(n471) );
  NAND2_X1 U601 ( .A1(n471), .A2(G125), .ZN(n475) );
  INV_X1 U602 ( .A(G125), .ZN(n472) );
  NAND2_X1 U603 ( .A1(n472), .A2(G146), .ZN(n474) );
  AND2_X1 U604 ( .A1(n475), .A2(n474), .ZN(n473) );
  NAND2_X1 U605 ( .A1(n473), .A2(KEYINPUT18), .ZN(n478) );
  INV_X1 U606 ( .A(KEYINPUT18), .ZN(n476) );
  NAND2_X1 U607 ( .A1(n500), .A2(n476), .ZN(n477) );
  NAND2_X1 U608 ( .A1(n478), .A2(n477), .ZN(n482) );
  NAND2_X1 U609 ( .A1(G224), .A2(n739), .ZN(n480) );
  XNOR2_X1 U610 ( .A(n525), .B(n483), .ZN(n484) );
  XNOR2_X1 U611 ( .A(n485), .B(n484), .ZN(n653) );
  INV_X1 U612 ( .A(n486), .ZN(n633) );
  OR2_X2 U613 ( .A1(n653), .A2(n633), .ZN(n488) );
  XNOR2_X1 U614 ( .A(n487), .B(KEYINPUT77), .ZN(n489) );
  XNOR2_X2 U615 ( .A(n488), .B(n356), .ZN(n612) );
  NAND2_X1 U616 ( .A1(G214), .A2(n489), .ZN(n693) );
  XOR2_X1 U617 ( .A(KEYINPUT11), .B(KEYINPUT94), .Z(n495) );
  XNOR2_X1 U618 ( .A(n495), .B(n494), .ZN(n499) );
  XOR2_X1 U619 ( .A(G113), .B(KEYINPUT12), .Z(n497) );
  NAND2_X1 U620 ( .A1(G214), .A2(n532), .ZN(n496) );
  XNOR2_X1 U621 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U622 ( .A(n499), .B(n498), .ZN(n506) );
  XNOR2_X1 U623 ( .A(n500), .B(G140), .ZN(n501) );
  XNOR2_X1 U624 ( .A(n502), .B(n501), .ZN(n550) );
  BUF_X1 U625 ( .A(n550), .Z(n744) );
  XOR2_X1 U626 ( .A(KEYINPUT95), .B(KEYINPUT93), .Z(n503) );
  XNOR2_X1 U627 ( .A(n504), .B(n503), .ZN(n505) );
  NOR2_X1 U628 ( .A1(G902), .A2(n636), .ZN(n509) );
  XNOR2_X1 U629 ( .A(KEYINPUT96), .B(KEYINPUT13), .ZN(n507) );
  XOR2_X1 U630 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n511) );
  NAND2_X1 U631 ( .A1(G234), .A2(n739), .ZN(n510) );
  XNOR2_X1 U632 ( .A(n511), .B(n510), .ZN(n555) );
  NAND2_X1 U633 ( .A1(G217), .A2(n555), .ZN(n513) );
  XNOR2_X1 U634 ( .A(n512), .B(n513), .ZN(n520) );
  XNOR2_X1 U635 ( .A(n514), .B(KEYINPUT97), .ZN(n518) );
  XOR2_X1 U636 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n516) );
  XNOR2_X1 U637 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U638 ( .A(n518), .B(n517), .Z(n519) );
  XNOR2_X1 U639 ( .A(n520), .B(n519), .ZN(n648) );
  AND2_X1 U640 ( .A1(n648), .A2(n544), .ZN(n522) );
  XNOR2_X1 U641 ( .A(KEYINPUT98), .B(KEYINPUT99), .ZN(n521) );
  XNOR2_X1 U642 ( .A(G478), .B(n572), .ZN(n523) );
  XNOR2_X1 U643 ( .A(G134), .B(G131), .ZN(n524) );
  XNOR2_X2 U644 ( .A(n525), .B(n524), .ZN(n542) );
  NAND2_X1 U645 ( .A1(n739), .A2(G227), .ZN(n526) );
  XNOR2_X1 U646 ( .A(n526), .B(G104), .ZN(n528) );
  XNOR2_X1 U647 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U648 ( .A(G469), .B(KEYINPUT72), .ZN(n531) );
  XNOR2_X1 U649 ( .A(n578), .B(KEYINPUT103), .ZN(n562) );
  XOR2_X1 U650 ( .A(G101), .B(KEYINPUT5), .Z(n534) );
  NAND2_X1 U651 ( .A1(n532), .A2(G210), .ZN(n533) );
  XNOR2_X1 U652 ( .A(n534), .B(n533), .ZN(n538) );
  BUF_X1 U653 ( .A(n539), .Z(n540) );
  XNOR2_X1 U654 ( .A(n541), .B(n540), .ZN(n543) );
  NAND2_X1 U655 ( .A1(n545), .A2(G217), .ZN(n546) );
  XNOR2_X1 U656 ( .A(G110), .B(KEYINPUT82), .ZN(n547) );
  XNOR2_X1 U657 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U658 ( .A(n550), .B(n549), .ZN(n559) );
  XOR2_X1 U659 ( .A(KEYINPUT24), .B(KEYINPUT78), .Z(n552) );
  XNOR2_X1 U660 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U661 ( .A(n554), .B(n553), .ZN(n557) );
  NAND2_X1 U662 ( .A1(G221), .A2(n555), .ZN(n556) );
  XNOR2_X1 U663 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U664 ( .A(n559), .B(n558), .ZN(n727) );
  NOR2_X1 U665 ( .A1(n727), .A2(G902), .ZN(n560) );
  NAND2_X1 U666 ( .A1(n601), .A2(n676), .ZN(n561) );
  NOR2_X1 U667 ( .A1(n609), .A2(n419), .ZN(n563) );
  NAND2_X1 U668 ( .A1(n563), .A2(n625), .ZN(n564) );
  XNOR2_X1 U669 ( .A(n564), .B(KEYINPUT80), .ZN(n565) );
  XNOR2_X1 U670 ( .A(KEYINPUT75), .B(KEYINPUT34), .ZN(n571) );
  INV_X1 U671 ( .A(n585), .ZN(n573) );
  NOR2_X1 U672 ( .A1(n573), .A2(n584), .ZN(n597) );
  XOR2_X1 U673 ( .A(KEYINPUT79), .B(n597), .Z(n574) );
  XNOR2_X1 U674 ( .A(KEYINPUT85), .B(KEYINPUT35), .ZN(n575) );
  NOR2_X1 U675 ( .A1(n609), .A2(n676), .ZN(n577) );
  NAND2_X1 U676 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U677 ( .A(n579), .B(KEYINPUT102), .ZN(n754) );
  NAND2_X1 U678 ( .A1(n581), .A2(n588), .ZN(n582) );
  XOR2_X1 U679 ( .A(n582), .B(KEYINPUT91), .Z(n583) );
  NAND2_X1 U680 ( .A1(n585), .A2(n584), .ZN(n605) );
  NOR2_X1 U681 ( .A1(n585), .A2(n584), .ZN(n670) );
  NOR2_X1 U682 ( .A1(n668), .A2(n670), .ZN(n700) );
  XOR2_X1 U683 ( .A(KEYINPUT84), .B(KEYINPUT45), .Z(n586) );
  INV_X1 U684 ( .A(n612), .ZN(n628) );
  XNOR2_X1 U685 ( .A(n588), .B(KEYINPUT106), .ZN(n596) );
  XNOR2_X1 U686 ( .A(KEYINPUT104), .B(n589), .ZN(n590) );
  NOR2_X1 U687 ( .A1(G900), .A2(n590), .ZN(n591) );
  NOR2_X1 U688 ( .A1(n592), .A2(n591), .ZN(n599) );
  XNOR2_X1 U689 ( .A(KEYINPUT30), .B(n593), .ZN(n594) );
  NOR2_X1 U690 ( .A1(n599), .A2(n594), .ZN(n595) );
  NAND2_X1 U691 ( .A1(n596), .A2(n595), .ZN(n613) );
  XNOR2_X1 U692 ( .A(KEYINPUT107), .B(n598), .ZN(n753) );
  NOR2_X1 U693 ( .A1(n599), .A2(n677), .ZN(n600) );
  NAND2_X1 U694 ( .A1(n676), .A2(n600), .ZN(n610) );
  NOR2_X1 U695 ( .A1(n610), .A2(n601), .ZN(n602) );
  XNOR2_X1 U696 ( .A(n602), .B(KEYINPUT28), .ZN(n621) );
  INV_X1 U697 ( .A(n670), .ZN(n607) );
  NOR2_X1 U698 ( .A1(n667), .A2(n664), .ZN(n608) );
  XOR2_X1 U699 ( .A(KEYINPUT108), .B(KEYINPUT40), .Z(n615) );
  XNOR2_X1 U700 ( .A(KEYINPUT38), .B(n612), .ZN(n617) );
  XNOR2_X1 U701 ( .A(KEYINPUT41), .B(KEYINPUT110), .ZN(n618) );
  XNOR2_X1 U702 ( .A(n619), .B(n618), .ZN(n675) );
  AND2_X1 U703 ( .A1(n623), .A2(n670), .ZN(n673) );
  XNOR2_X1 U704 ( .A(KEYINPUT105), .B(n624), .ZN(n626) );
  INV_X1 U705 ( .A(n625), .ZN(n682) );
  NAND2_X1 U706 ( .A1(n626), .A2(n682), .ZN(n627) );
  XNOR2_X1 U707 ( .A(n627), .B(KEYINPUT43), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n629), .A2(n628), .ZN(n674) );
  INV_X1 U709 ( .A(n674), .ZN(n630) );
  NOR2_X1 U710 ( .A1(n673), .A2(n630), .ZN(n631) );
  XNOR2_X1 U711 ( .A(n713), .B(KEYINPUT2), .ZN(n634) );
  NAND2_X1 U712 ( .A1(n347), .A2(G475), .ZN(n637) );
  INV_X1 U713 ( .A(G952), .ZN(n638) );
  AND2_X1 U714 ( .A1(n638), .A2(G953), .ZN(n730) );
  XNOR2_X1 U715 ( .A(KEYINPUT60), .B(KEYINPUT66), .ZN(n639) );
  XOR2_X1 U716 ( .A(G125), .B(KEYINPUT37), .Z(n640) );
  XNOR2_X1 U717 ( .A(n641), .B(n640), .ZN(G27) );
  XNOR2_X1 U718 ( .A(G122), .B(KEYINPUT126), .ZN(n643) );
  XNOR2_X1 U719 ( .A(n644), .B(n643), .ZN(G24) );
  NAND2_X1 U720 ( .A1(n346), .A2(G472), .ZN(n646) );
  XOR2_X1 U721 ( .A(KEYINPUT86), .B(KEYINPUT63), .Z(n647) );
  NAND2_X1 U722 ( .A1(n725), .A2(G478), .ZN(n649) );
  NAND2_X1 U723 ( .A1(n347), .A2(G469), .ZN(n652) );
  XOR2_X1 U724 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n650) );
  NAND2_X1 U725 ( .A1(n725), .A2(G210), .ZN(n656) );
  XOR2_X1 U726 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n654) );
  NAND2_X1 U727 ( .A1(n659), .A2(n668), .ZN(n657) );
  XNOR2_X1 U728 ( .A(n657), .B(KEYINPUT112), .ZN(n658) );
  XNOR2_X1 U729 ( .A(G104), .B(n658), .ZN(G6) );
  XOR2_X1 U730 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n661) );
  NAND2_X1 U731 ( .A1(n659), .A2(n670), .ZN(n660) );
  XNOR2_X1 U732 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U733 ( .A(G107), .B(n662), .ZN(G9) );
  XOR2_X1 U734 ( .A(n663), .B(G110), .Z(G12) );
  XOR2_X1 U735 ( .A(KEYINPUT113), .B(KEYINPUT29), .Z(n666) );
  XNOR2_X1 U736 ( .A(G128), .B(n664), .ZN(n665) );
  XNOR2_X1 U737 ( .A(n666), .B(n665), .ZN(G30) );
  XOR2_X1 U738 ( .A(G146), .B(n667), .Z(G48) );
  NAND2_X1 U739 ( .A1(n671), .A2(n668), .ZN(n669) );
  XNOR2_X1 U740 ( .A(n669), .B(G113), .ZN(G15) );
  NAND2_X1 U741 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U742 ( .A(n672), .B(G116), .ZN(G18) );
  XOR2_X1 U743 ( .A(G134), .B(n673), .Z(G36) );
  XNOR2_X1 U744 ( .A(G140), .B(n674), .ZN(G42) );
  XOR2_X1 U745 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n679) );
  NAND2_X1 U746 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U747 ( .A(n679), .B(n678), .ZN(n680) );
  XOR2_X1 U748 ( .A(KEYINPUT114), .B(n680), .Z(n686) );
  NAND2_X1 U749 ( .A1(n682), .A2(n681), .ZN(n684) );
  XOR2_X1 U750 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n683) );
  XNOR2_X1 U751 ( .A(n684), .B(n683), .ZN(n685) );
  NAND2_X1 U752 ( .A1(n686), .A2(n357), .ZN(n688) );
  NAND2_X1 U753 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U754 ( .A(n689), .B(KEYINPUT117), .Z(n690) );
  XNOR2_X1 U755 ( .A(KEYINPUT51), .B(n690), .ZN(n691) );
  NOR2_X1 U756 ( .A1(n675), .A2(n691), .ZN(n706) );
  NOR2_X1 U757 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U758 ( .A(n695), .B(KEYINPUT118), .ZN(n696) );
  NOR2_X1 U759 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U760 ( .A(KEYINPUT119), .B(n698), .Z(n702) );
  NOR2_X1 U761 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U762 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U763 ( .A1(n381), .A2(n703), .ZN(n704) );
  XNOR2_X1 U764 ( .A(n704), .B(KEYINPUT120), .ZN(n705) );
  NOR2_X1 U765 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U766 ( .A(n707), .B(KEYINPUT52), .ZN(n708) );
  NOR2_X1 U767 ( .A1(n709), .A2(n708), .ZN(n711) );
  NOR2_X1 U768 ( .A1(n675), .A2(n381), .ZN(n710) );
  NOR2_X1 U769 ( .A1(n711), .A2(n710), .ZN(n721) );
  INV_X1 U770 ( .A(KEYINPUT83), .ZN(n712) );
  NAND2_X1 U771 ( .A1(n713), .A2(n712), .ZN(n714) );
  BUF_X1 U772 ( .A(n715), .Z(n716) );
  NAND2_X1 U773 ( .A1(n717), .A2(KEYINPUT83), .ZN(n718) );
  NAND2_X1 U774 ( .A1(n721), .A2(n720), .ZN(n722) );
  BUF_X1 U775 ( .A(n346), .Z(n726) );
  NAND2_X1 U776 ( .A1(n726), .A2(G217), .ZN(n728) );
  XNOR2_X1 U777 ( .A(n728), .B(n727), .ZN(n729) );
  NOR2_X1 U778 ( .A1(n730), .A2(n729), .ZN(G66) );
  NAND2_X1 U779 ( .A1(n716), .A2(n739), .ZN(n734) );
  NAND2_X1 U780 ( .A1(G953), .A2(G224), .ZN(n731) );
  XNOR2_X1 U781 ( .A(KEYINPUT61), .B(n731), .ZN(n732) );
  NAND2_X1 U782 ( .A1(n732), .A2(G898), .ZN(n733) );
  NAND2_X1 U783 ( .A1(n734), .A2(n733), .ZN(n743) );
  BUF_X1 U784 ( .A(n735), .Z(n736) );
  BUF_X1 U785 ( .A(n737), .Z(n738) );
  XOR2_X1 U786 ( .A(n736), .B(n738), .Z(n741) );
  NOR2_X1 U787 ( .A1(G898), .A2(n739), .ZN(n740) );
  NOR2_X1 U788 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U789 ( .A(n743), .B(n742), .ZN(G69) );
  NOR2_X1 U790 ( .A1(G953), .A2(n745), .ZN(n746) );
  XNOR2_X1 U791 ( .A(KEYINPUT125), .B(n746), .ZN(n751) );
  XOR2_X1 U792 ( .A(G227), .B(n747), .Z(n748) );
  NAND2_X1 U793 ( .A1(n748), .A2(G900), .ZN(n749) );
  NAND2_X1 U794 ( .A1(n749), .A2(G953), .ZN(n750) );
  NAND2_X1 U795 ( .A1(n751), .A2(n750), .ZN(G72) );
  XOR2_X1 U796 ( .A(n752), .B(G131), .Z(G33) );
  XOR2_X1 U797 ( .A(n415), .B(n753), .Z(G45) );
  XNOR2_X1 U798 ( .A(G101), .B(n754), .ZN(G3) );
  XNOR2_X1 U799 ( .A(KEYINPUT127), .B(n755), .ZN(G21) );
  XOR2_X1 U800 ( .A(G137), .B(n756), .Z(G39) );
endmodule

