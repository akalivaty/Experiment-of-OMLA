

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798;

  INV_X1 U375 ( .A(n604), .ZN(n354) );
  BUF_X1 U376 ( .A(G113), .Z(n356) );
  XNOR2_X1 U377 ( .A(n373), .B(G116), .ZN(n372) );
  XNOR2_X1 U378 ( .A(G119), .B(KEYINPUT3), .ZN(n465) );
  AND2_X2 U379 ( .A1(n384), .A2(n383), .ZN(n365) );
  XNOR2_X1 U380 ( .A(n580), .B(KEYINPUT41), .ZN(n752) );
  NOR2_X1 U381 ( .A1(n355), .A2(n354), .ZN(n394) );
  INV_X1 U382 ( .A(n395), .ZN(n355) );
  NAND2_X2 U383 ( .A1(n363), .A2(n396), .ZN(n422) );
  BUF_X2 U384 ( .A(n625), .Z(n641) );
  XOR2_X1 U385 ( .A(G140), .B(n356), .Z(n500) );
  BUF_X1 U386 ( .A(n759), .Z(n357) );
  AND2_X2 U387 ( .A1(n447), .A2(n442), .ZN(n441) );
  AND2_X2 U388 ( .A1(n436), .A2(n435), .ZN(n434) );
  INV_X1 U389 ( .A(n723), .ZN(n622) );
  AND2_X2 U390 ( .A1(n393), .A2(n394), .ZN(n363) );
  XNOR2_X2 U391 ( .A(n624), .B(n623), .ZN(n753) );
  NOR2_X2 U392 ( .A1(n716), .A2(n737), .ZN(n522) );
  XNOR2_X2 U393 ( .A(KEYINPUT32), .B(n633), .ZN(n798) );
  XNOR2_X2 U394 ( .A(n375), .B(n475), .ZN(n411) );
  INV_X2 U395 ( .A(G113), .ZN(n373) );
  NOR2_X1 U396 ( .A1(n676), .A2(n796), .ZN(n583) );
  NOR2_X1 U397 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U398 ( .A(n659), .B(n414), .ZN(n660) );
  NOR2_X1 U399 ( .A1(n417), .A2(n362), .ZN(n683) );
  NAND2_X1 U400 ( .A1(n419), .A2(n368), .ZN(n417) );
  XNOR2_X1 U401 ( .A(n422), .B(KEYINPUT35), .ZN(n795) );
  XNOR2_X1 U402 ( .A(n639), .B(n380), .ZN(n711) );
  XNOR2_X1 U403 ( .A(n487), .B(KEYINPUT0), .ZN(n625) );
  NOR2_X1 U404 ( .A1(n389), .A2(n737), .ZN(n580) );
  NAND2_X1 U405 ( .A1(n461), .A2(n622), .ZN(n624) );
  XNOR2_X1 U406 ( .A(n613), .B(n570), .ZN(n735) );
  XNOR2_X1 U407 ( .A(n382), .B(n482), .ZN(n592) );
  XNOR2_X1 U408 ( .A(n524), .B(KEYINPUT22), .ZN(n525) );
  XNOR2_X1 U409 ( .A(G146), .B(G125), .ZN(n494) );
  NAND2_X1 U410 ( .A1(n526), .A2(n525), .ZN(n360) );
  NAND2_X1 U411 ( .A1(n358), .A2(n359), .ZN(n361) );
  NAND2_X1 U412 ( .A1(n360), .A2(n361), .ZN(n627) );
  INV_X1 U413 ( .A(n526), .ZN(n358) );
  INV_X1 U414 ( .A(n525), .ZN(n359) );
  NAND2_X1 U415 ( .A1(n711), .A2(n697), .ZN(n379) );
  AND2_X1 U416 ( .A1(n457), .A2(n794), .ZN(n456) );
  INV_X1 U417 ( .A(KEYINPUT39), .ZN(n454) );
  AND2_X1 U418 ( .A1(n392), .A2(n621), .ZN(n461) );
  INV_X1 U419 ( .A(n576), .ZN(n720) );
  XNOR2_X1 U420 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n516) );
  XNOR2_X1 U421 ( .A(G104), .B(G122), .ZN(n492) );
  INV_X1 U422 ( .A(G140), .ZN(n527) );
  AND2_X1 U423 ( .A1(n378), .A2(n646), .ZN(n647) );
  NAND2_X1 U424 ( .A1(n379), .A2(n645), .ZN(n378) );
  NOR2_X1 U425 ( .A1(n650), .A2(KEYINPUT44), .ZN(n652) );
  INV_X1 U426 ( .A(G472), .ZN(n450) );
  NOR2_X1 U427 ( .A1(G237), .A2(G953), .ZN(n469) );
  XNOR2_X1 U428 ( .A(n399), .B(n464), .ZN(n529) );
  XNOR2_X1 U429 ( .A(G131), .B(G134), .ZN(n464) );
  XNOR2_X1 U430 ( .A(n391), .B(n390), .ZN(n774) );
  INV_X1 U431 ( .A(G104), .ZN(n390) );
  XNOR2_X1 U432 ( .A(G107), .B(G110), .ZN(n391) );
  INV_X2 U433 ( .A(G953), .ZN(n788) );
  XNOR2_X1 U434 ( .A(n494), .B(KEYINPUT10), .ZN(n781) );
  XNOR2_X1 U435 ( .A(G107), .B(G122), .ZN(n511) );
  XOR2_X1 U436 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n512) );
  AND2_X1 U437 ( .A1(n750), .A2(KEYINPUT65), .ZN(n448) );
  NAND2_X1 U438 ( .A1(n445), .A2(n443), .ZN(n442) );
  NAND2_X1 U439 ( .A1(n488), .A2(n446), .ZN(n445) );
  NAND2_X1 U440 ( .A1(n657), .A2(n444), .ZN(n443) );
  NAND2_X1 U441 ( .A1(KEYINPUT2), .A2(n446), .ZN(n444) );
  XNOR2_X1 U442 ( .A(n774), .B(n473), .ZN(n532) );
  INV_X1 U443 ( .A(KEYINPUT75), .ZN(n414) );
  INV_X1 U444 ( .A(n708), .ZN(n451) );
  NAND2_X1 U445 ( .A1(n423), .A2(n452), .ZN(n401) );
  NOR2_X1 U446 ( .A1(n571), .A2(n454), .ZN(n452) );
  NOR2_X1 U447 ( .A1(n641), .A2(KEYINPUT34), .ZN(n397) );
  OR2_X1 U448 ( .A1(n693), .A2(G902), .ZN(n555) );
  NOR2_X1 U449 ( .A1(n428), .A2(KEYINPUT73), .ZN(n387) );
  XNOR2_X1 U450 ( .A(n381), .B(KEYINPUT16), .ZN(n476) );
  INV_X1 U451 ( .A(KEYINPUT71), .ZN(n381) );
  INV_X1 U452 ( .A(KEYINPUT65), .ZN(n446) );
  XNOR2_X1 U453 ( .A(n494), .B(KEYINPUT88), .ZN(n413) );
  XNOR2_X1 U454 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n410) );
  XNOR2_X1 U455 ( .A(n514), .B(n463), .ZN(n399) );
  INV_X1 U456 ( .A(KEYINPUT4), .ZN(n463) );
  NOR2_X1 U457 ( .A1(n576), .A2(n586), .ZN(n557) );
  XNOR2_X1 U458 ( .A(n479), .B(n478), .ZN(n569) );
  NAND2_X1 U459 ( .A1(n416), .A2(n415), .ZN(n487) );
  XOR2_X1 U460 ( .A(G146), .B(G137), .Z(n466) );
  XNOR2_X1 U461 ( .A(KEYINPUT24), .B(KEYINPUT90), .ZN(n543) );
  XNOR2_X1 U462 ( .A(G128), .B(G119), .ZN(n538) );
  XNOR2_X1 U463 ( .A(n504), .B(n503), .ZN(n662) );
  XNOR2_X1 U464 ( .A(n502), .B(n501), .ZN(n503) );
  BUF_X1 U465 ( .A(n753), .Z(n374) );
  NAND2_X1 U466 ( .A1(n720), .A2(KEYINPUT66), .ZN(n418) );
  NOR2_X1 U467 ( .A1(n720), .A2(KEYINPUT66), .ZN(n420) );
  XNOR2_X1 U468 ( .A(G134), .B(G116), .ZN(n510) );
  AND2_X2 U469 ( .A1(n661), .A2(n660), .ZN(n759) );
  NAND2_X1 U470 ( .A1(n440), .A2(n371), .ZN(n439) );
  AND2_X1 U471 ( .A1(n665), .A2(G953), .ZN(n763) );
  XNOR2_X1 U472 ( .A(n532), .B(n366), .ZN(n533) );
  INV_X1 U473 ( .A(G146), .ZN(n530) );
  AND2_X1 U474 ( .A1(n367), .A2(n660), .ZN(n755) );
  XNOR2_X1 U475 ( .A(n455), .B(n572), .ZN(n676) );
  NAND2_X1 U476 ( .A1(n400), .A2(n401), .ZN(n455) );
  AND2_X1 U477 ( .A1(n424), .A2(n364), .ZN(n400) );
  INV_X1 U478 ( .A(KEYINPUT96), .ZN(n380) );
  XNOR2_X1 U479 ( .A(n377), .B(KEYINPUT82), .ZN(n376) );
  NOR2_X1 U480 ( .A1(n626), .A2(n392), .ZN(n377) );
  AND2_X1 U481 ( .A1(n626), .A2(KEYINPUT66), .ZN(n362) );
  AND2_X1 U482 ( .A1(n453), .A2(n451), .ZN(n364) );
  XOR2_X1 U483 ( .A(n531), .B(n530), .Z(n366) );
  XNOR2_X1 U484 ( .A(n481), .B(KEYINPUT76), .ZN(n482) );
  NAND2_X1 U485 ( .A1(n751), .A2(n750), .ZN(n367) );
  AND2_X1 U486 ( .A1(n418), .A2(n717), .ZN(n368) );
  AND2_X1 U487 ( .A1(n424), .A2(n453), .ZN(n369) );
  XNOR2_X1 U488 ( .A(KEYINPUT109), .B(KEYINPUT28), .ZN(n370) );
  XNOR2_X1 U489 ( .A(n555), .B(n554), .ZN(n717) );
  AND2_X1 U490 ( .A1(n657), .A2(n446), .ZN(n371) );
  NOR2_X1 U491 ( .A1(n686), .A2(n657), .ZN(n479) );
  NAND2_X1 U492 ( .A1(n398), .A2(n397), .ZN(n396) );
  XNOR2_X2 U493 ( .A(n372), .B(n465), .ZN(n477) );
  NOR2_X2 U494 ( .A1(n625), .A2(n523), .ZN(n526) );
  AND2_X1 U495 ( .A1(n797), .A2(KEYINPUT81), .ZN(n459) );
  INV_X1 U496 ( .A(n476), .ZN(n375) );
  NAND2_X1 U497 ( .A1(n421), .A2(n420), .ZN(n419) );
  NAND2_X1 U498 ( .A1(n611), .A2(n723), .ZN(n612) );
  AND2_X1 U499 ( .A1(n587), .A2(n460), .ZN(n611) );
  NAND2_X1 U500 ( .A1(n433), .A2(n432), .ZN(n431) );
  XNOR2_X1 U501 ( .A(n577), .B(n370), .ZN(n579) );
  NAND2_X1 U502 ( .A1(n458), .A2(n438), .ZN(n457) );
  NAND2_X1 U503 ( .A1(n376), .A2(n630), .ZN(n646) );
  INV_X1 U504 ( .A(n592), .ZN(n416) );
  NAND2_X1 U505 ( .A1(n569), .A2(n734), .ZN(n382) );
  NOR2_X2 U506 ( .A1(n428), .A2(n437), .ZN(n388) );
  NAND2_X1 U507 ( .A1(n385), .A2(n365), .ZN(n656) );
  NAND2_X1 U508 ( .A1(n437), .A2(KEYINPUT73), .ZN(n383) );
  NAND2_X1 U509 ( .A1(n428), .A2(KEYINPUT73), .ZN(n384) );
  NAND2_X1 U510 ( .A1(n387), .A2(n386), .ZN(n385) );
  INV_X1 U511 ( .A(n437), .ZN(n386) );
  AND2_X1 U512 ( .A1(n388), .A2(KEYINPUT2), .ZN(n658) );
  XNOR2_X1 U513 ( .A(n388), .B(n787), .ZN(n789) );
  NAND2_X1 U514 ( .A1(n749), .A2(n388), .ZN(n751) );
  NOR2_X1 U515 ( .A1(n732), .A2(n389), .ZN(n733) );
  NAND2_X1 U516 ( .A1(n735), .A2(n734), .ZN(n389) );
  NAND2_X1 U517 ( .A1(n392), .A2(n584), .ZN(n585) );
  XNOR2_X1 U518 ( .A(n392), .B(KEYINPUT78), .ZN(n628) );
  XNOR2_X2 U519 ( .A(n576), .B(KEYINPUT6), .ZN(n392) );
  NAND2_X1 U520 ( .A1(n753), .A2(KEYINPUT34), .ZN(n393) );
  NAND2_X1 U521 ( .A1(n641), .A2(KEYINPUT34), .ZN(n395) );
  INV_X1 U522 ( .A(n753), .ZN(n398) );
  XNOR2_X1 U523 ( .A(n399), .B(n532), .ZN(n407) );
  NAND2_X1 U524 ( .A1(n369), .A2(n401), .ZN(n618) );
  XNOR2_X1 U525 ( .A(n529), .B(n467), .ZN(n405) );
  INV_X1 U526 ( .A(n646), .ZN(n635) );
  NAND2_X1 U527 ( .A1(n627), .A2(n723), .ZN(n626) );
  XNOR2_X1 U528 ( .A(n783), .B(n533), .ZN(n671) );
  XNOR2_X1 U529 ( .A(n405), .B(n472), .ZN(n678) );
  OR2_X2 U530 ( .A1(n678), .A2(G902), .ZN(n425) );
  NAND2_X1 U531 ( .A1(n402), .A2(KEYINPUT80), .ZN(n406) );
  NAND2_X1 U532 ( .A1(n404), .A2(n403), .ZN(n402) );
  INV_X1 U533 ( .A(KEYINPUT47), .ZN(n403) );
  INV_X1 U534 ( .A(n706), .ZN(n404) );
  NOR2_X1 U535 ( .A1(n593), .A2(n592), .ZN(n702) );
  NOR2_X1 U536 ( .A1(n609), .A2(KEYINPUT48), .ZN(n432) );
  NAND2_X1 U537 ( .A1(n406), .A2(n645), .ZN(n600) );
  XNOR2_X1 U538 ( .A(n408), .B(n407), .ZN(n686) );
  XNOR2_X1 U539 ( .A(n409), .B(n772), .ZN(n408) );
  XNOR2_X1 U540 ( .A(n412), .B(n413), .ZN(n409) );
  XNOR2_X2 U541 ( .A(n477), .B(n411), .ZN(n772) );
  XNOR2_X1 U542 ( .A(n474), .B(n410), .ZN(n412) );
  NOR2_X1 U543 ( .A1(n745), .A2(n485), .ZN(n415) );
  INV_X1 U544 ( .A(n626), .ZN(n421) );
  NOR2_X1 U545 ( .A1(n795), .A2(n683), .ZN(n634) );
  INV_X1 U546 ( .A(n601), .ZN(n423) );
  NAND2_X1 U547 ( .A1(n568), .A2(n567), .ZN(n601) );
  NAND2_X1 U548 ( .A1(n601), .A2(n454), .ZN(n424) );
  XNOR2_X2 U549 ( .A(n425), .B(n450), .ZN(n576) );
  NAND2_X1 U550 ( .A1(n426), .A2(n438), .ZN(n427) );
  NAND2_X1 U551 ( .A1(n434), .A2(n431), .ZN(n426) );
  NAND2_X2 U552 ( .A1(n427), .A2(n456), .ZN(n428) );
  NOR2_X2 U553 ( .A1(n430), .A2(n429), .ZN(n437) );
  INV_X1 U554 ( .A(n434), .ZN(n429) );
  NAND2_X1 U555 ( .A1(n431), .A2(n459), .ZN(n430) );
  INV_X1 U556 ( .A(n610), .ZN(n433) );
  NAND2_X1 U557 ( .A1(n609), .A2(KEYINPUT48), .ZN(n435) );
  NAND2_X1 U558 ( .A1(n610), .A2(KEYINPUT48), .ZN(n436) );
  INV_X1 U559 ( .A(KEYINPUT81), .ZN(n438) );
  NAND2_X1 U560 ( .A1(n441), .A2(n439), .ZN(n661) );
  INV_X1 U561 ( .A(n449), .ZN(n440) );
  NAND2_X1 U562 ( .A1(n449), .A2(n448), .ZN(n447) );
  NAND2_X1 U563 ( .A1(n656), .A2(n749), .ZN(n449) );
  NAND2_X1 U564 ( .A1(n571), .A2(n454), .ZN(n453) );
  INV_X1 U565 ( .A(n797), .ZN(n458) );
  NOR2_X1 U566 ( .A1(n708), .A2(n586), .ZN(n460) );
  INV_X1 U567 ( .A(KEYINPUT67), .ZN(n524) );
  XNOR2_X1 U568 ( .A(n477), .B(n466), .ZN(n467) );
  XNOR2_X1 U569 ( .A(n471), .B(n470), .ZN(n472) );
  INV_X1 U570 ( .A(KEYINPUT19), .ZN(n481) );
  XNOR2_X1 U571 ( .A(n588), .B(KEYINPUT110), .ZN(n589) );
  XNOR2_X1 U572 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X2 U573 ( .A(G128), .B(KEYINPUT64), .ZN(n462) );
  XNOR2_X2 U574 ( .A(n462), .B(G143), .ZN(n514) );
  XOR2_X1 U575 ( .A(KEYINPUT68), .B(G101), .Z(n473) );
  XNOR2_X1 U576 ( .A(n473), .B(KEYINPUT5), .ZN(n468) );
  XNOR2_X1 U577 ( .A(n468), .B(KEYINPUT95), .ZN(n471) );
  XNOR2_X1 U578 ( .A(n469), .B(KEYINPUT74), .ZN(n498) );
  AND2_X1 U579 ( .A1(G210), .A2(n498), .ZN(n470) );
  AND2_X1 U580 ( .A1(G224), .A2(n788), .ZN(n474) );
  XNOR2_X1 U581 ( .A(KEYINPUT72), .B(G122), .ZN(n475) );
  XNOR2_X1 U582 ( .A(G902), .B(KEYINPUT15), .ZN(n488) );
  INV_X1 U583 ( .A(n488), .ZN(n657) );
  OR2_X1 U584 ( .A1(G237), .A2(G902), .ZN(n480) );
  NAND2_X1 U585 ( .A1(G210), .A2(n480), .ZN(n478) );
  NAND2_X1 U586 ( .A1(G214), .A2(n480), .ZN(n734) );
  NAND2_X1 U587 ( .A1(G952), .A2(n788), .ZN(n562) );
  INV_X1 U588 ( .A(n562), .ZN(n484) );
  NAND2_X1 U589 ( .A1(G953), .A2(G902), .ZN(n558) );
  NOR2_X1 U590 ( .A1(G898), .A2(n558), .ZN(n483) );
  NOR2_X1 U591 ( .A1(n484), .A2(n483), .ZN(n485) );
  NAND2_X1 U592 ( .A1(G234), .A2(G237), .ZN(n486) );
  XOR2_X1 U593 ( .A(KEYINPUT14), .B(n486), .Z(n745) );
  INV_X1 U594 ( .A(n745), .ZN(n560) );
  NAND2_X1 U595 ( .A1(n488), .A2(G234), .ZN(n489) );
  XNOR2_X1 U596 ( .A(n489), .B(KEYINPUT20), .ZN(n548) );
  NAND2_X1 U597 ( .A1(n548), .A2(G221), .ZN(n491) );
  INV_X1 U598 ( .A(KEYINPUT21), .ZN(n490) );
  XNOR2_X1 U599 ( .A(n491), .B(n490), .ZN(n573) );
  INV_X1 U600 ( .A(n573), .ZN(n716) );
  XOR2_X1 U601 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n493) );
  XNOR2_X1 U602 ( .A(n493), .B(n492), .ZN(n497) );
  XNOR2_X1 U603 ( .A(KEYINPUT99), .B(KEYINPUT11), .ZN(n495) );
  XNOR2_X1 U604 ( .A(n781), .B(n495), .ZN(n496) );
  XOR2_X1 U605 ( .A(n497), .B(n496), .Z(n504) );
  NAND2_X1 U606 ( .A1(G214), .A2(n498), .ZN(n502) );
  XNOR2_X1 U607 ( .A(G143), .B(G131), .ZN(n499) );
  XNOR2_X1 U608 ( .A(n500), .B(n499), .ZN(n501) );
  INV_X1 U609 ( .A(G902), .ZN(n505) );
  NAND2_X1 U610 ( .A1(n662), .A2(n505), .ZN(n509) );
  XOR2_X1 U611 ( .A(KEYINPUT101), .B(KEYINPUT13), .Z(n507) );
  XNOR2_X1 U612 ( .A(KEYINPUT100), .B(G475), .ZN(n506) );
  XNOR2_X1 U613 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X2 U614 ( .A(n509), .B(n508), .ZN(n603) );
  XNOR2_X1 U615 ( .A(n510), .B(KEYINPUT102), .ZN(n520) );
  XNOR2_X1 U616 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U617 ( .A(n514), .B(n513), .Z(n518) );
  NAND2_X1 U618 ( .A1(n788), .A2(G234), .ZN(n515) );
  XNOR2_X1 U619 ( .A(n516), .B(n515), .ZN(n537) );
  NAND2_X1 U620 ( .A1(G217), .A2(n537), .ZN(n517) );
  XNOR2_X1 U621 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U622 ( .A(n520), .B(n519), .ZN(n760) );
  NOR2_X1 U623 ( .A1(n760), .A2(G902), .ZN(n521) );
  XNOR2_X1 U624 ( .A(G478), .B(n521), .ZN(n602) );
  NAND2_X1 U625 ( .A1(n603), .A2(n602), .ZN(n737) );
  XNOR2_X1 U626 ( .A(n522), .B(KEYINPUT103), .ZN(n523) );
  XNOR2_X1 U627 ( .A(n527), .B(G137), .ZN(n539) );
  INV_X1 U628 ( .A(n539), .ZN(n528) );
  XNOR2_X1 U629 ( .A(n529), .B(n528), .ZN(n783) );
  NAND2_X1 U630 ( .A1(G227), .A2(n788), .ZN(n531) );
  NOR2_X1 U631 ( .A1(n671), .A2(G902), .ZN(n535) );
  INV_X1 U632 ( .A(G469), .ZN(n534) );
  XNOR2_X2 U633 ( .A(n535), .B(n534), .ZN(n578) );
  INV_X1 U634 ( .A(KEYINPUT1), .ZN(n536) );
  XNOR2_X2 U635 ( .A(n578), .B(n536), .ZN(n723) );
  NAND2_X1 U636 ( .A1(n537), .A2(G221), .ZN(n542) );
  XNOR2_X1 U637 ( .A(n538), .B(KEYINPUT89), .ZN(n540) );
  XNOR2_X1 U638 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U639 ( .A(n542), .B(n541), .ZN(n547) );
  XNOR2_X1 U640 ( .A(G110), .B(KEYINPUT23), .ZN(n544) );
  XNOR2_X1 U641 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U642 ( .A(n781), .B(n545), .ZN(n546) );
  XNOR2_X1 U643 ( .A(n547), .B(n546), .ZN(n693) );
  AND2_X1 U644 ( .A1(n548), .A2(G217), .ZN(n553) );
  XNOR2_X1 U645 ( .A(KEYINPUT93), .B(KEYINPUT25), .ZN(n549) );
  XNOR2_X1 U646 ( .A(n549), .B(KEYINPUT77), .ZN(n551) );
  XNOR2_X1 U647 ( .A(KEYINPUT91), .B(KEYINPUT92), .ZN(n550) );
  XNOR2_X1 U648 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U649 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U650 ( .A(n635), .B(G101), .Z(G3) );
  INV_X1 U651 ( .A(n734), .ZN(n586) );
  XNOR2_X1 U652 ( .A(KEYINPUT108), .B(KEYINPUT30), .ZN(n556) );
  XNOR2_X1 U653 ( .A(n557), .B(n556), .ZN(n566) );
  NOR2_X1 U654 ( .A1(G900), .A2(n558), .ZN(n559) );
  NAND2_X1 U655 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U656 ( .A(KEYINPUT104), .B(n561), .Z(n564) );
  NOR2_X1 U657 ( .A1(n562), .A2(n745), .ZN(n563) );
  NOR2_X1 U658 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U659 ( .A(n565), .B(KEYINPUT79), .ZN(n574) );
  AND2_X1 U660 ( .A1(n566), .A2(n574), .ZN(n568) );
  OR2_X1 U661 ( .A1(n717), .A2(n716), .ZN(n722) );
  INV_X1 U662 ( .A(n722), .ZN(n621) );
  NAND2_X1 U663 ( .A1(n578), .A2(n621), .ZN(n640) );
  XNOR2_X1 U664 ( .A(n640), .B(KEYINPUT107), .ZN(n567) );
  BUF_X2 U665 ( .A(n569), .Z(n613) );
  INV_X1 U666 ( .A(KEYINPUT38), .ZN(n570) );
  INV_X1 U667 ( .A(n735), .ZN(n571) );
  INV_X1 U668 ( .A(n602), .ZN(n594) );
  OR2_X1 U669 ( .A1(n603), .A2(n594), .ZN(n708) );
  INV_X1 U670 ( .A(KEYINPUT40), .ZN(n572) );
  INV_X1 U671 ( .A(n717), .ZN(n630) );
  NAND2_X1 U672 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U673 ( .A1(n630), .A2(n575), .ZN(n584) );
  NAND2_X1 U674 ( .A1(n584), .A2(n720), .ZN(n577) );
  NAND2_X1 U675 ( .A1(n579), .A2(n578), .ZN(n593) );
  NOR2_X1 U676 ( .A1(n593), .A2(n752), .ZN(n581) );
  XNOR2_X1 U677 ( .A(n581), .B(KEYINPUT42), .ZN(n796) );
  INV_X1 U678 ( .A(KEYINPUT46), .ZN(n582) );
  XNOR2_X1 U679 ( .A(n583), .B(n582), .ZN(n610) );
  XNOR2_X1 U680 ( .A(n585), .B(KEYINPUT105), .ZN(n587) );
  AND2_X1 U681 ( .A1(n613), .A2(n611), .ZN(n590) );
  XNOR2_X1 U682 ( .A(KEYINPUT36), .B(KEYINPUT84), .ZN(n588) );
  AND2_X1 U683 ( .A1(n591), .A2(n622), .ZN(n714) );
  INV_X1 U684 ( .A(n714), .ZN(n608) );
  INV_X1 U685 ( .A(n702), .ZN(n706) );
  AND2_X1 U686 ( .A1(n603), .A2(n594), .ZN(n701) );
  INV_X1 U687 ( .A(n701), .ZN(n710) );
  NAND2_X1 U688 ( .A1(n710), .A2(n708), .ZN(n645) );
  INV_X1 U689 ( .A(n645), .ZN(n732) );
  NAND2_X1 U690 ( .A1(n732), .A2(KEYINPUT80), .ZN(n595) );
  NAND2_X1 U691 ( .A1(n595), .A2(n702), .ZN(n596) );
  NAND2_X1 U692 ( .A1(n596), .A2(KEYINPUT47), .ZN(n598) );
  OR2_X1 U693 ( .A1(KEYINPUT80), .A2(KEYINPUT47), .ZN(n597) );
  AND2_X1 U694 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U695 ( .A1(n600), .A2(n599), .ZN(n606) );
  NAND2_X1 U696 ( .A1(n604), .A2(n613), .ZN(n605) );
  NOR2_X1 U697 ( .A1(n601), .A2(n605), .ZN(n705) );
  NOR2_X1 U698 ( .A1(n606), .A2(n705), .ZN(n607) );
  NAND2_X1 U699 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U700 ( .A(n612), .B(KEYINPUT43), .ZN(n615) );
  INV_X1 U701 ( .A(n613), .ZN(n614) );
  AND2_X1 U702 ( .A1(n615), .A2(n614), .ZN(n617) );
  INV_X1 U703 ( .A(KEYINPUT106), .ZN(n616) );
  XNOR2_X1 U704 ( .A(n617), .B(n616), .ZN(n797) );
  OR2_X1 U705 ( .A1(n618), .A2(n710), .ZN(n620) );
  INV_X1 U706 ( .A(KEYINPUT111), .ZN(n619) );
  XNOR2_X1 U707 ( .A(n620), .B(n619), .ZN(n794) );
  XOR2_X1 U708 ( .A(KEYINPUT86), .B(KEYINPUT33), .Z(n623) );
  INV_X1 U709 ( .A(n627), .ZN(n629) );
  NOR2_X1 U710 ( .A1(n629), .A2(n628), .ZN(n632) );
  NOR2_X1 U711 ( .A1(n723), .A2(n630), .ZN(n631) );
  NAND2_X1 U712 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U713 ( .A1(n634), .A2(n798), .ZN(n650) );
  NAND2_X1 U714 ( .A1(n650), .A2(KEYINPUT44), .ZN(n648) );
  INV_X1 U715 ( .A(n720), .ZN(n643) );
  NOR2_X1 U716 ( .A1(n643), .A2(n722), .ZN(n636) );
  NAND2_X1 U717 ( .A1(n622), .A2(n636), .ZN(n728) );
  NOR2_X1 U718 ( .A1(n641), .A2(n728), .ZN(n638) );
  XNOR2_X1 U719 ( .A(KEYINPUT97), .B(KEYINPUT31), .ZN(n637) );
  XNOR2_X1 U720 ( .A(n638), .B(n637), .ZN(n639) );
  NOR2_X1 U721 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U722 ( .A(n642), .B(KEYINPUT94), .ZN(n644) );
  NAND2_X1 U723 ( .A1(n644), .A2(n643), .ZN(n697) );
  NAND2_X1 U724 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U725 ( .A(n649), .B(KEYINPUT83), .ZN(n654) );
  INV_X1 U726 ( .A(KEYINPUT70), .ZN(n651) );
  XNOR2_X1 U727 ( .A(n652), .B(n651), .ZN(n653) );
  NAND2_X1 U728 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X2 U729 ( .A(n655), .B(KEYINPUT45), .ZN(n749) );
  INV_X1 U730 ( .A(KEYINPUT2), .ZN(n750) );
  NAND2_X1 U731 ( .A1(n749), .A2(n658), .ZN(n659) );
  NAND2_X1 U732 ( .A1(n759), .A2(G475), .ZN(n664) );
  XOR2_X1 U733 ( .A(KEYINPUT59), .B(n662), .Z(n663) );
  XNOR2_X1 U734 ( .A(n664), .B(n663), .ZN(n666) );
  INV_X1 U735 ( .A(G952), .ZN(n665) );
  INV_X1 U736 ( .A(n763), .ZN(n689) );
  NAND2_X1 U737 ( .A1(n666), .A2(n689), .ZN(n668) );
  INV_X1 U738 ( .A(KEYINPUT60), .ZN(n667) );
  XNOR2_X1 U739 ( .A(n668), .B(n667), .ZN(G60) );
  NAND2_X1 U740 ( .A1(n759), .A2(G469), .ZN(n673) );
  XNOR2_X1 U741 ( .A(KEYINPUT118), .B(KEYINPUT57), .ZN(n669) );
  XNOR2_X1 U742 ( .A(n669), .B(KEYINPUT58), .ZN(n670) );
  XNOR2_X1 U743 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U744 ( .A(n673), .B(n672), .ZN(n674) );
  NAND2_X1 U745 ( .A1(n674), .A2(n689), .ZN(n675) );
  XNOR2_X1 U746 ( .A(n675), .B(KEYINPUT119), .ZN(G54) );
  XOR2_X1 U747 ( .A(n676), .B(G131), .Z(G33) );
  NAND2_X1 U748 ( .A1(n759), .A2(G472), .ZN(n680) );
  XNOR2_X1 U749 ( .A(KEYINPUT87), .B(KEYINPUT62), .ZN(n677) );
  XNOR2_X1 U750 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U751 ( .A(n680), .B(n679), .ZN(n681) );
  NAND2_X1 U752 ( .A1(n681), .A2(n689), .ZN(n682) );
  XNOR2_X1 U753 ( .A(n682), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U754 ( .A(n683), .B(G110), .Z(G12) );
  NAND2_X1 U755 ( .A1(n759), .A2(G210), .ZN(n688) );
  XNOR2_X1 U756 ( .A(KEYINPUT85), .B(KEYINPUT54), .ZN(n684) );
  XOR2_X1 U757 ( .A(n684), .B(KEYINPUT55), .Z(n685) );
  XNOR2_X1 U758 ( .A(n686), .B(n685), .ZN(n687) );
  XNOR2_X1 U759 ( .A(n688), .B(n687), .ZN(n690) );
  NAND2_X1 U760 ( .A1(n690), .A2(n689), .ZN(n692) );
  INV_X1 U761 ( .A(KEYINPUT56), .ZN(n691) );
  XNOR2_X1 U762 ( .A(n692), .B(n691), .ZN(G51) );
  NAND2_X1 U763 ( .A1(n357), .A2(G217), .ZN(n694) );
  XNOR2_X1 U764 ( .A(n694), .B(n693), .ZN(n695) );
  NOR2_X1 U765 ( .A1(n695), .A2(n763), .ZN(G66) );
  NOR2_X1 U766 ( .A1(n708), .A2(n697), .ZN(n696) );
  XOR2_X1 U767 ( .A(G104), .B(n696), .Z(G6) );
  NOR2_X1 U768 ( .A1(n710), .A2(n697), .ZN(n699) );
  XNOR2_X1 U769 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n698) );
  XNOR2_X1 U770 ( .A(n699), .B(n698), .ZN(n700) );
  XNOR2_X1 U771 ( .A(G107), .B(n700), .ZN(G9) );
  XOR2_X1 U772 ( .A(G128), .B(KEYINPUT29), .Z(n704) );
  NAND2_X1 U773 ( .A1(n404), .A2(n701), .ZN(n703) );
  XNOR2_X1 U774 ( .A(n704), .B(n703), .ZN(G30) );
  XOR2_X1 U775 ( .A(G143), .B(n705), .Z(G45) );
  OR2_X1 U776 ( .A1(n706), .A2(n708), .ZN(n707) );
  XNOR2_X1 U777 ( .A(n707), .B(G146), .ZN(G48) );
  NOR2_X1 U778 ( .A1(n711), .A2(n708), .ZN(n709) );
  XOR2_X1 U779 ( .A(n356), .B(n709), .Z(G15) );
  NOR2_X1 U780 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U781 ( .A(KEYINPUT112), .B(n712), .Z(n713) );
  XNOR2_X1 U782 ( .A(G116), .B(n713), .ZN(G18) );
  XNOR2_X1 U783 ( .A(G125), .B(n714), .ZN(n715) );
  XNOR2_X1 U784 ( .A(n715), .B(KEYINPUT37), .ZN(G27) );
  NAND2_X1 U785 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U786 ( .A(n718), .B(KEYINPUT49), .ZN(n719) );
  NOR2_X1 U787 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U788 ( .A(n721), .B(KEYINPUT114), .ZN(n727) );
  NAND2_X1 U789 ( .A1(n723), .A2(n722), .ZN(n725) );
  XOR2_X1 U790 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n724) );
  XNOR2_X1 U791 ( .A(n725), .B(n724), .ZN(n726) );
  NAND2_X1 U792 ( .A1(n727), .A2(n726), .ZN(n729) );
  NAND2_X1 U793 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U794 ( .A(KEYINPUT51), .B(n730), .ZN(n731) );
  NOR2_X1 U795 ( .A1(n752), .A2(n731), .ZN(n742) );
  XNOR2_X1 U796 ( .A(KEYINPUT116), .B(n733), .ZN(n739) );
  NOR2_X1 U797 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U798 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U799 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U800 ( .A1(n374), .A2(n740), .ZN(n741) );
  NOR2_X1 U801 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U802 ( .A(n743), .B(KEYINPUT52), .ZN(n744) );
  NOR2_X1 U803 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U804 ( .A1(n746), .A2(G952), .ZN(n747) );
  XNOR2_X1 U805 ( .A(KEYINPUT117), .B(n747), .ZN(n748) );
  NOR2_X1 U806 ( .A1(G953), .A2(n748), .ZN(n757) );
  NOR2_X1 U807 ( .A1(n374), .A2(n752), .ZN(n754) );
  NOR2_X1 U808 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U809 ( .A1(n757), .A2(n756), .ZN(n758) );
  XOR2_X1 U810 ( .A(KEYINPUT53), .B(n758), .Z(G75) );
  NAND2_X1 U811 ( .A1(n357), .A2(G478), .ZN(n761) );
  XNOR2_X1 U812 ( .A(n761), .B(n760), .ZN(n762) );
  NOR2_X1 U813 ( .A1(n763), .A2(n762), .ZN(G63) );
  INV_X1 U814 ( .A(n749), .ZN(n764) );
  NOR2_X1 U815 ( .A1(G953), .A2(n764), .ZN(n765) );
  XNOR2_X1 U816 ( .A(KEYINPUT121), .B(n765), .ZN(n770) );
  NAND2_X1 U817 ( .A1(G953), .A2(G224), .ZN(n766) );
  XNOR2_X1 U818 ( .A(KEYINPUT61), .B(n766), .ZN(n767) );
  NAND2_X1 U819 ( .A1(n767), .A2(G898), .ZN(n768) );
  XNOR2_X1 U820 ( .A(KEYINPUT120), .B(n768), .ZN(n769) );
  NAND2_X1 U821 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U822 ( .A(n771), .B(KEYINPUT124), .ZN(n780) );
  XOR2_X1 U823 ( .A(n772), .B(KEYINPUT122), .Z(n773) );
  XNOR2_X1 U824 ( .A(n774), .B(n773), .ZN(n775) );
  XNOR2_X1 U825 ( .A(n775), .B(G101), .ZN(n777) );
  NOR2_X1 U826 ( .A1(n788), .A2(G898), .ZN(n776) );
  NOR2_X1 U827 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U828 ( .A(n778), .B(KEYINPUT123), .Z(n779) );
  XNOR2_X1 U829 ( .A(n780), .B(n779), .ZN(G69) );
  XNOR2_X1 U830 ( .A(n781), .B(KEYINPUT125), .ZN(n782) );
  XNOR2_X1 U831 ( .A(n783), .B(n782), .ZN(n787) );
  XNOR2_X1 U832 ( .A(n787), .B(KEYINPUT127), .ZN(n784) );
  XNOR2_X1 U833 ( .A(G227), .B(n784), .ZN(n785) );
  NAND2_X1 U834 ( .A1(n785), .A2(G900), .ZN(n786) );
  NAND2_X1 U835 ( .A1(n786), .A2(G953), .ZN(n792) );
  NAND2_X1 U836 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U837 ( .A(KEYINPUT126), .B(n790), .ZN(n791) );
  NAND2_X1 U838 ( .A1(n792), .A2(n791), .ZN(G72) );
  XOR2_X1 U839 ( .A(G134), .B(KEYINPUT113), .Z(n793) );
  XNOR2_X1 U840 ( .A(n794), .B(n793), .ZN(G36) );
  XOR2_X1 U841 ( .A(n795), .B(G122), .Z(G24) );
  XOR2_X1 U842 ( .A(n796), .B(G137), .Z(G39) );
  XNOR2_X1 U843 ( .A(n797), .B(G140), .ZN(G42) );
  XNOR2_X1 U844 ( .A(G119), .B(n798), .ZN(G21) );
endmodule

