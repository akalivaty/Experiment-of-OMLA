//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 1 1 0 0 0 1 0 0 1 1 0 0 1 0 0 1 0 0 1 0 1 1 1 1 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT67), .B1(new_n188), .B2(G116), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT67), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G119), .ZN(new_n192));
  AND2_X1   g006(.A1(new_n189), .A2(new_n192), .ZN(new_n193));
  XOR2_X1   g007(.A(KEYINPUT2), .B(G113), .Z(new_n194));
  OAI21_X1  g008(.A(KEYINPUT66), .B1(new_n191), .B2(G119), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT66), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(new_n188), .A3(G116), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n193), .A2(new_n194), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n194), .B1(new_n193), .B2(new_n198), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT30), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT64), .B1(new_n205), .B2(G137), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT11), .ZN(new_n207));
  AND2_X1   g021(.A1(KEYINPUT65), .A2(G131), .ZN(new_n208));
  NOR2_X1   g022(.A1(KEYINPUT65), .A2(G131), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT11), .ZN(new_n211));
  OAI211_X1 g025(.A(KEYINPUT64), .B(new_n211), .C1(new_n205), .C2(G137), .ZN(new_n212));
  INV_X1    g026(.A(G137), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(G134), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n207), .A2(new_n210), .A3(new_n212), .A4(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n205), .A2(G137), .ZN(new_n217));
  OAI21_X1  g031(.A(G131), .B1(new_n217), .B2(new_n214), .ZN(new_n218));
  INV_X1    g032(.A(G143), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT1), .B1(new_n219), .B2(G146), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n219), .A2(G146), .ZN(new_n221));
  INV_X1    g035(.A(G146), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n222), .A2(G143), .ZN(new_n223));
  OAI211_X1 g037(.A(G128), .B(new_n220), .C1(new_n221), .C2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(G143), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n219), .A2(G146), .ZN(new_n226));
  INV_X1    g040(.A(G128), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n225), .B(new_n226), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n224), .A2(KEYINPUT68), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(KEYINPUT68), .B1(new_n224), .B2(new_n228), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n216), .B(new_n218), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  AND2_X1   g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n225), .A2(new_n226), .A3(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(G143), .B(G146), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT0), .B(G128), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n216), .ZN(new_n238));
  INV_X1    g052(.A(G131), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n214), .B1(new_n206), .B2(KEYINPUT11), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n239), .B1(new_n240), .B2(new_n212), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n237), .B1(new_n238), .B2(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n204), .B1(new_n231), .B2(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n216), .A2(new_n218), .A3(new_n228), .A4(new_n224), .ZN(new_n244));
  AND3_X1   g058(.A1(new_n242), .A2(new_n244), .A3(new_n204), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n203), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n229), .A2(new_n230), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n216), .A2(new_n218), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n202), .B(new_n242), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(G237), .A2(G953), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G210), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n252), .B(KEYINPUT27), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT26), .B(G101), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n253), .B(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n250), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT29), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n249), .A2(KEYINPUT28), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT28), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n231), .A2(new_n260), .A3(new_n202), .A4(new_n242), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n242), .A2(new_n244), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n203), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n257), .B(new_n258), .C1(new_n256), .C2(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT71), .B(G902), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n224), .A2(new_n228), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT68), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n224), .A2(KEYINPUT68), .A3(new_n228), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n248), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n240), .A2(new_n212), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G131), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n236), .B1(new_n275), .B2(new_n216), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n203), .B1(new_n273), .B2(new_n276), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n262), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n256), .A2(new_n258), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n268), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n187), .B1(new_n266), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n281), .B(KEYINPUT72), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT32), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT69), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n249), .A2(new_n255), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT30), .B1(new_n273), .B2(new_n276), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n242), .A2(new_n204), .A3(new_n244), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n285), .B1(new_n288), .B2(new_n203), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT31), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n284), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n249), .A2(new_n255), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n246), .A2(new_n292), .A3(new_n284), .A4(new_n290), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n259), .A2(new_n261), .B1(new_n203), .B2(new_n263), .ZN(new_n296));
  OAI22_X1  g110(.A1(new_n289), .A2(new_n290), .B1(new_n296), .B2(new_n255), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT70), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n246), .A2(new_n292), .A3(new_n290), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT69), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n293), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT70), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n246), .A2(new_n292), .ZN(new_n303));
  AOI22_X1  g117(.A1(new_n256), .A2(new_n265), .B1(new_n303), .B2(KEYINPUT31), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n301), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n298), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(G472), .A2(G902), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n283), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n307), .ZN(new_n309));
  AOI211_X1 g123(.A(KEYINPUT32), .B(new_n309), .C1(new_n298), .C2(new_n305), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n282), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G953), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(G221), .A3(G234), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n313), .B(KEYINPUT77), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT22), .B(G137), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n314), .B(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT73), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n317), .B1(new_n227), .B2(G119), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n227), .A2(G119), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n188), .A2(KEYINPUT73), .A3(G128), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT24), .B(G110), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G140), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G125), .ZN(new_n325));
  INV_X1    g139(.A(G125), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G140), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n327), .A3(KEYINPUT16), .ZN(new_n328));
  OR3_X1    g142(.A1(new_n326), .A2(KEYINPUT16), .A3(G140), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n222), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n328), .A2(new_n329), .A3(G146), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n323), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT74), .B1(new_n188), .B2(G128), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT23), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT23), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n319), .A2(KEYINPUT74), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n188), .A2(G128), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n335), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n339), .A2(KEYINPUT75), .A3(G110), .ZN(new_n340));
  AOI21_X1  g154(.A(KEYINPUT75), .B1(new_n339), .B2(G110), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n333), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT78), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n321), .A2(new_n322), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n344), .B1(new_n339), .B2(G110), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n325), .A2(new_n327), .A3(new_n222), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(KEYINPUT76), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n345), .A2(new_n332), .A3(new_n347), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n342), .A2(new_n343), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n343), .B1(new_n342), .B2(new_n348), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n316), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n342), .A2(new_n343), .A3(new_n348), .ZN(new_n352));
  INV_X1    g166(.A(new_n316), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n351), .A2(new_n267), .A3(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT79), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n356), .A2(KEYINPUT25), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n357), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n351), .A2(new_n267), .A3(new_n354), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G217), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n362), .B1(new_n267), .B2(G234), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n351), .A2(new_n354), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n363), .A2(G902), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n366), .B(KEYINPUT80), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n364), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(G214), .B1(G237), .B2(G902), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT91), .ZN(new_n374));
  INV_X1    g188(.A(G224), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT7), .B1(new_n375), .B2(G953), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n236), .A2(G125), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n269), .A2(new_n326), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n377), .B1(new_n378), .B2(KEYINPUT90), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT90), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n380), .B1(new_n269), .B2(new_n326), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n376), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n377), .A2(KEYINPUT87), .ZN(new_n383));
  INV_X1    g197(.A(new_n376), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT87), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n236), .A2(new_n385), .A3(G125), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n383), .A2(new_n384), .A3(new_n378), .A4(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n382), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(G110), .B(G122), .ZN(new_n389));
  XOR2_X1   g203(.A(new_n389), .B(KEYINPUT8), .Z(new_n390));
  NAND4_X1  g204(.A1(new_n198), .A2(KEYINPUT5), .A3(new_n189), .A4(new_n192), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT88), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT88), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n193), .A2(new_n393), .A3(KEYINPUT5), .A4(new_n198), .ZN(new_n394));
  NOR3_X1   g208(.A1(new_n191), .A2(KEYINPUT5), .A3(G119), .ZN(new_n395));
  INV_X1    g209(.A(G113), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT89), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT89), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n188), .A2(G116), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n398), .B(G113), .C1(new_n399), .C2(KEYINPUT5), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n392), .A2(new_n394), .A3(new_n397), .A4(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(G104), .ZN(new_n402));
  OAI21_X1  g216(.A(KEYINPUT3), .B1(new_n402), .B2(G107), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT3), .ZN(new_n404));
  INV_X1    g218(.A(G107), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(new_n405), .A3(G104), .ZN(new_n406));
  INV_X1    g220(.A(G101), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n402), .A2(G107), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n403), .A2(new_n406), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n402), .A2(G107), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n405), .A2(G104), .ZN(new_n411));
  OAI21_X1  g225(.A(G101), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AND2_X1   g226(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n199), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n401), .A2(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n395), .A2(new_n396), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n391), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n413), .B1(new_n418), .B2(new_n199), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n390), .B1(new_n416), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n374), .B1(new_n388), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n403), .A2(new_n406), .A3(new_n408), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G101), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(KEYINPUT4), .A3(new_n409), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n423), .A2(G101), .A3(new_n426), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n425), .B(new_n427), .C1(new_n200), .C2(new_n201), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n418), .A2(new_n199), .A3(new_n413), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n428), .A2(new_n389), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n390), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n397), .A2(new_n400), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n432), .B1(KEYINPUT88), .B2(new_n391), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n414), .B1(new_n433), .B2(new_n394), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n431), .B1(new_n434), .B2(new_n419), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n435), .A2(KEYINPUT91), .A3(new_n382), .A4(new_n387), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n422), .A2(new_n430), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n383), .A2(new_n378), .A3(new_n386), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n375), .A2(G953), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n438), .B(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n389), .B1(new_n428), .B2(new_n429), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT86), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT6), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n441), .B1(new_n430), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n441), .A2(new_n444), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n440), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(G902), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n437), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(G210), .B1(G237), .B2(G902), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n430), .A2(new_n444), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n446), .B1(new_n454), .B2(new_n441), .ZN(new_n455));
  AOI21_X1  g269(.A(G902), .B1(new_n455), .B2(new_n440), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n456), .A2(new_n437), .A3(new_n451), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n373), .B1(new_n453), .B2(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT9), .B(G234), .ZN(new_n459));
  OAI21_X1  g273(.A(G221), .B1(new_n459), .B2(G902), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n238), .A2(new_n241), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  AND2_X1   g276(.A1(new_n423), .A2(G101), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n409), .A2(KEYINPUT4), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n237), .B(new_n427), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT82), .B(KEYINPUT10), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n409), .A2(new_n412), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n466), .B1(new_n269), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n409), .A2(new_n412), .A3(KEYINPUT10), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n470), .B1(new_n271), .B2(new_n272), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n462), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  OAI211_X1 g286(.A(KEYINPUT10), .B(new_n413), .C1(new_n229), .C2(new_n230), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n473), .A2(new_n461), .A3(new_n465), .A4(new_n468), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(G110), .B(G140), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n312), .A2(G227), .ZN(new_n477));
  XOR2_X1   g291(.A(new_n476), .B(new_n477), .Z(new_n478));
  NAND2_X1  g292(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT85), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT83), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n482), .B1(new_n269), .B2(new_n467), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n269), .A2(new_n467), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n269), .A2(new_n467), .A3(new_n482), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n462), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT12), .ZN(new_n489));
  OR2_X1    g303(.A1(new_n489), .A2(KEYINPUT84), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(KEYINPUT84), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n488), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n478), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n487), .A2(KEYINPUT84), .A3(new_n489), .A4(new_n462), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n492), .A2(new_n493), .A3(new_n494), .A4(new_n474), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n475), .A2(KEYINPUT85), .A3(new_n478), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n481), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G469), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(new_n498), .A3(new_n267), .ZN(new_n499));
  NAND2_X1  g313(.A1(G469), .A2(G902), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n475), .A2(new_n478), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n492), .A2(new_n494), .A3(new_n474), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n501), .B1(new_n502), .B2(new_n478), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(G469), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n499), .A2(new_n500), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n458), .A2(new_n460), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT96), .ZN(new_n507));
  NOR2_X1   g321(.A1(G475), .A2(G902), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  XOR2_X1   g323(.A(G113), .B(G122), .Z(new_n510));
  XOR2_X1   g324(.A(KEYINPUT93), .B(G104), .Z(new_n511));
  XOR2_X1   g325(.A(new_n510), .B(new_n511), .Z(new_n512));
  NAND2_X1  g326(.A1(new_n325), .A2(new_n327), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(G146), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n346), .A2(KEYINPUT76), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT76), .ZN(new_n516));
  XNOR2_X1  g330(.A(G125), .B(G140), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n516), .B1(new_n517), .B2(new_n222), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n514), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(G237), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n312), .A3(G214), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n219), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n251), .A2(G143), .A3(G214), .ZN(new_n523));
  NAND3_X1  g337(.A1(KEYINPUT92), .A2(KEYINPUT18), .A3(G131), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n524), .ZN(new_n526));
  AND4_X1   g340(.A1(G143), .A2(new_n520), .A3(new_n312), .A4(G214), .ZN(new_n527));
  AOI21_X1  g341(.A(G143), .B1(new_n251), .B2(G214), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n519), .A2(new_n525), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT94), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n328), .A2(G146), .A3(new_n329), .ZN(new_n532));
  AOI21_X1  g346(.A(G146), .B1(new_n328), .B2(new_n329), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n331), .A2(KEYINPUT94), .A3(new_n332), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OR2_X1    g350(.A1(new_n208), .A2(new_n209), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n537), .B(KEYINPUT17), .C1(new_n527), .C2(new_n528), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n537), .B1(new_n527), .B2(new_n528), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n522), .A2(new_n210), .A3(new_n523), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n538), .B1(new_n541), .B2(KEYINPUT17), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n512), .B(new_n530), .C1(new_n536), .C2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n512), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n325), .A2(new_n327), .A3(KEYINPUT19), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT19), .B1(new_n325), .B2(new_n327), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n222), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n541), .A2(new_n547), .A3(new_n332), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n529), .A2(new_n525), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n549), .B1(new_n347), .B2(new_n514), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n544), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n543), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT95), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n543), .A2(new_n551), .A3(KEYINPUT95), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n509), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT20), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n507), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n555), .ZN(new_n559));
  AOI21_X1  g373(.A(KEYINPUT95), .B1(new_n543), .B2(new_n551), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n508), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n561), .A2(KEYINPUT96), .A3(KEYINPUT20), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n509), .A2(KEYINPUT20), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n552), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n558), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  OR2_X1    g379(.A1(new_n536), .A2(new_n542), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n512), .B1(new_n566), .B2(new_n530), .ZN(new_n567));
  INV_X1    g381(.A(new_n543), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n449), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(G475), .ZN(new_n570));
  INV_X1    g384(.A(G952), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(G953), .ZN(new_n572));
  INV_X1    g386(.A(G234), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n572), .B1(new_n573), .B2(new_n520), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  AOI211_X1 g389(.A(new_n312), .B(new_n267), .C1(G234), .C2(G237), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT21), .B(G898), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n219), .A2(G128), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n227), .A2(G143), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(new_n205), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n191), .A2(KEYINPUT14), .A3(G122), .ZN(new_n584));
  XNOR2_X1  g398(.A(G116), .B(G122), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  OAI211_X1 g400(.A(G107), .B(new_n584), .C1(new_n586), .C2(KEYINPUT14), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n583), .B(new_n587), .C1(G107), .C2(new_n586), .ZN(new_n588));
  INV_X1    g402(.A(new_n580), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n589), .A2(KEYINPUT13), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n581), .B1(new_n589), .B2(KEYINPUT13), .ZN(new_n591));
  OAI21_X1  g405(.A(G134), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n582), .A2(new_n205), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n585), .B(new_n405), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n459), .A2(new_n362), .A3(G953), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n588), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n596), .B1(new_n588), .B2(new_n595), .ZN(new_n598));
  OR2_X1    g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(G478), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n599), .B(new_n267), .C1(KEYINPUT15), .C2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n267), .B1(new_n597), .B2(new_n598), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT15), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n602), .A2(new_n603), .A3(G478), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n565), .A2(new_n570), .A3(new_n579), .A4(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n506), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n311), .A2(new_n371), .A3(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G101), .ZN(G3));
  NAND2_X1  g424(.A1(new_n565), .A2(new_n570), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT33), .ZN(new_n613));
  OAI22_X1  g427(.A1(new_n597), .A2(new_n598), .B1(KEYINPUT97), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n268), .A2(new_n600), .ZN(new_n615));
  XNOR2_X1  g429(.A(KEYINPUT97), .B(KEYINPUT33), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n614), .B(new_n615), .C1(new_n599), .C2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n602), .A2(new_n600), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n612), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n453), .A2(new_n457), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n623), .A2(new_n372), .A3(new_n579), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n301), .A2(new_n302), .A3(new_n304), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n302), .B1(new_n301), .B2(new_n304), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n267), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AOI22_X1  g442(.A1(new_n628), .A2(G472), .B1(new_n306), .B2(new_n307), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n505), .A2(new_n460), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(new_n370), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n625), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT34), .B(G104), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G6));
  INV_X1    g449(.A(new_n624), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n554), .A2(new_n555), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n563), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n558), .A2(new_n562), .A3(new_n638), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n639), .A2(new_n570), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n636), .A2(new_n605), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n632), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT35), .B(G107), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  NOR2_X1   g458(.A1(new_n353), .A2(KEYINPUT36), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n342), .A2(new_n348), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n368), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n364), .A2(KEYINPUT98), .A3(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT98), .ZN(new_n650));
  INV_X1    g464(.A(new_n363), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n651), .B1(new_n358), .B2(new_n360), .ZN(new_n652));
  INV_X1    g466(.A(new_n648), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n650), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n649), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n608), .A2(new_n629), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT37), .B(G110), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G12));
  INV_X1    g472(.A(new_n655), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n307), .B1(new_n626), .B2(new_n627), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(KEYINPUT32), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n306), .A2(new_n283), .A3(new_n307), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n659), .B1(new_n663), .B2(new_n282), .ZN(new_n664));
  INV_X1    g478(.A(new_n506), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n640), .A2(new_n605), .ZN(new_n666));
  INV_X1    g480(.A(G900), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n575), .B1(new_n576), .B2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n664), .A2(new_n665), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G128), .ZN(G30));
  NOR2_X1   g485(.A1(new_n612), .A2(new_n606), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n659), .A2(new_n672), .A3(new_n372), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n673), .B(KEYINPUT99), .Z(new_n674));
  AOI21_X1  g488(.A(new_n255), .B1(new_n277), .B2(new_n249), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n449), .B1(new_n289), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(G472), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n663), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n623), .B(KEYINPUT38), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT100), .B(KEYINPUT39), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n668), .B(new_n680), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n630), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(new_n682), .B(KEYINPUT40), .Z(new_n683));
  NAND4_X1  g497(.A1(new_n674), .A2(new_n678), .A3(new_n679), .A4(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT101), .B(G143), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G45));
  AOI211_X1 g500(.A(new_n668), .B(new_n620), .C1(new_n565), .C2(new_n570), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n664), .A2(new_n665), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G146), .ZN(G48));
  AOI21_X1  g503(.A(new_n370), .B1(new_n663), .B2(new_n282), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n497), .A2(new_n267), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(G469), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n692), .A2(new_n460), .A3(new_n499), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n690), .A2(new_n625), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT41), .B(G113), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G15));
  NAND3_X1  g511(.A1(new_n690), .A2(new_n641), .A3(new_n694), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G116), .ZN(G18));
  INV_X1    g513(.A(KEYINPUT102), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n450), .A2(new_n452), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n451), .B1(new_n456), .B2(new_n437), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n372), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n700), .B1(new_n693), .B2(new_n703), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n497), .A2(new_n498), .A3(new_n267), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n498), .B1(new_n497), .B2(new_n267), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n707), .A2(new_n458), .A3(KEYINPUT102), .A4(new_n460), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n607), .B1(new_n704), .B2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n709), .A2(new_n311), .A3(new_n655), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G119), .ZN(G21));
  OAI221_X1 g525(.A(new_n301), .B1(new_n290), .B2(new_n289), .C1(new_n255), .C2(new_n278), .ZN(new_n712));
  AOI22_X1  g526(.A1(new_n628), .A2(G472), .B1(new_n307), .B2(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n624), .A2(new_n693), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n713), .A2(new_n672), .A3(new_n714), .A4(new_n371), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G122), .ZN(G24));
  AND2_X1   g530(.A1(new_n704), .A2(new_n708), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n713), .A2(new_n655), .A3(new_n687), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(new_n326), .ZN(G27));
  INV_X1    g534(.A(KEYINPUT104), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n502), .A2(new_n478), .ZN(new_n722));
  OAI21_X1  g536(.A(KEYINPUT103), .B1(new_n475), .B2(new_n478), .ZN(new_n723));
  OR3_X1    g537(.A1(new_n475), .A2(KEYINPUT103), .A3(new_n478), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n722), .A2(G469), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n499), .A2(new_n500), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n460), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n453), .A2(new_n372), .A3(new_n457), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n721), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n728), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n730), .A2(KEYINPUT104), .A3(new_n460), .A4(new_n726), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n311), .A2(new_n732), .A3(new_n371), .A4(new_n687), .ZN(new_n733));
  XOR2_X1   g547(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n736), .B1(new_n308), .B2(new_n310), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n661), .A2(new_n662), .A3(KEYINPUT106), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n282), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n687), .A2(KEYINPUT42), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n740), .B1(new_n729), .B2(new_n731), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n739), .A2(new_n371), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n735), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G131), .ZN(G33));
  NAND4_X1  g558(.A1(new_n311), .A2(new_n732), .A3(new_n371), .A4(new_n669), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G134), .ZN(G36));
  NOR2_X1   g560(.A1(new_n611), .A2(new_n620), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(KEYINPUT43), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n629), .A2(new_n659), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n730), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT44), .B1(new_n748), .B2(new_n749), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n752), .B1(KEYINPUT108), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n754), .B1(KEYINPUT108), .B2(new_n753), .ZN(new_n755));
  OR2_X1    g569(.A1(new_n755), .A2(KEYINPUT109), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(KEYINPUT109), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n722), .A2(KEYINPUT45), .A3(new_n723), .A4(new_n724), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n758), .B(G469), .C1(KEYINPUT45), .C2(new_n503), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n759), .A2(new_n500), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(KEYINPUT46), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n759), .A2(KEYINPUT46), .A3(new_n500), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n499), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n761), .B1(KEYINPUT107), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n764), .B1(KEYINPUT107), .B2(new_n763), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n460), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n681), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n756), .A2(new_n757), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G137), .ZN(G39));
  INV_X1    g583(.A(KEYINPUT47), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n765), .A2(KEYINPUT47), .A3(new_n460), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n687), .A2(new_n370), .A3(new_n730), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n311), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G140), .ZN(G42));
  XOR2_X1   g591(.A(new_n707), .B(KEYINPUT49), .Z(new_n778));
  NAND3_X1  g592(.A1(new_n371), .A2(new_n372), .A3(new_n460), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n778), .A2(new_n679), .A3(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n678), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(new_n781), .A3(new_n747), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n783));
  INV_X1    g597(.A(new_n719), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n672), .A2(new_n372), .A3(new_n623), .ZN(new_n785));
  NOR4_X1   g599(.A1(new_n727), .A2(new_n652), .A3(new_n653), .A4(new_n668), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(new_n678), .A3(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n784), .A2(new_n670), .A3(new_n688), .A4(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n788), .B(new_n789), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n690), .B(new_n694), .C1(new_n625), .C2(new_n641), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n619), .B1(new_n565), .B2(new_n570), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n792), .B1(new_n612), .B2(new_n606), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n629), .A2(new_n793), .A3(new_n636), .A4(new_n631), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n794), .A2(new_n715), .A3(new_n656), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n791), .A2(new_n795), .A3(new_n609), .A4(new_n710), .ZN(new_n796));
  XOR2_X1   g610(.A(new_n281), .B(KEYINPUT72), .Z(new_n797));
  AOI21_X1  g611(.A(new_n797), .B1(new_n663), .B2(new_n736), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n370), .B1(new_n798), .B2(new_n738), .ZN(new_n799));
  AOI22_X1  g613(.A1(new_n799), .A2(new_n741), .B1(new_n733), .B2(new_n734), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n505), .A2(new_n460), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n605), .A2(new_n668), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n639), .A2(new_n570), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT110), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n639), .A2(new_n570), .A3(KEYINPUT110), .A4(new_n803), .ZN(new_n807));
  AND4_X1   g621(.A1(new_n802), .A2(new_n806), .A3(new_n730), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n628), .A2(G472), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n712), .A2(new_n307), .ZN(new_n810));
  AND4_X1   g624(.A1(new_n809), .A2(new_n687), .A3(new_n655), .A4(new_n810), .ZN(new_n811));
  AOI22_X1  g625(.A1(new_n664), .A2(new_n808), .B1(new_n811), .B2(new_n732), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT111), .B1(new_n812), .B2(new_n745), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n808), .A2(new_n311), .A3(new_n655), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n811), .A2(new_n732), .ZN(new_n815));
  AND4_X1   g629(.A1(KEYINPUT111), .A2(new_n745), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT112), .B1(new_n801), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n710), .A2(new_n609), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n794), .A2(new_n715), .A3(new_n656), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n743), .A2(new_n821), .A3(new_n791), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n745), .A2(new_n814), .A3(new_n815), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT111), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n812), .A2(KEYINPUT111), .A3(new_n745), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT112), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n822), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n790), .B1(new_n818), .B2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n788), .B(KEYINPUT52), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n801), .A2(new_n817), .A3(KEYINPUT112), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n828), .B1(new_n822), .B2(new_n827), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n784), .A2(new_n670), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT53), .B1(new_n837), .B2(KEYINPUT52), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n783), .B1(new_n832), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n822), .A2(new_n827), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n837), .A2(KEYINPUT52), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n790), .A2(new_n842), .A3(KEYINPUT53), .A4(new_n843), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n783), .B(new_n844), .C1(new_n836), .C2(KEYINPUT53), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT113), .B1(new_n841), .B2(new_n846), .ZN(new_n847));
  AOI211_X1 g661(.A(new_n838), .B(new_n833), .C1(new_n835), .C2(new_n834), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n834), .A2(new_n835), .ZN(new_n849));
  AOI21_X1  g663(.A(KEYINPUT53), .B1(new_n849), .B2(new_n790), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT54), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT113), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n851), .A2(new_n852), .A3(new_n845), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n693), .A2(new_n728), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n781), .A2(new_n371), .A3(new_n575), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n748), .A2(new_n575), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n713), .A2(new_n371), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  OAI221_X1 g673(.A(new_n572), .B1(new_n622), .B2(new_n855), .C1(new_n859), .C2(new_n717), .ZN(new_n860));
  INV_X1    g674(.A(new_n799), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n748), .A2(new_n575), .A3(new_n854), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n864), .A2(KEYINPUT48), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(KEYINPUT48), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n860), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n705), .A2(new_n706), .A3(new_n460), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n730), .B(new_n858), .C1(new_n773), .C2(new_n868), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n855), .A2(new_n611), .A3(new_n619), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n713), .A2(new_n655), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n862), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n694), .A2(new_n373), .ZN(new_n875));
  OR2_X1    g689(.A1(new_n875), .A2(KEYINPUT114), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT50), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n679), .B1(KEYINPUT115), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n875), .A2(KEYINPUT114), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n858), .A2(new_n876), .A3(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n877), .A2(KEYINPUT115), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n881), .A2(new_n882), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n883), .A2(KEYINPUT51), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n867), .B1(new_n874), .B2(new_n885), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n881), .A2(new_n882), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n881), .A2(new_n882), .ZN(new_n888));
  OAI21_X1  g702(.A(KEYINPUT116), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT116), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n883), .A2(new_n890), .A3(new_n884), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n869), .A2(new_n889), .A3(new_n891), .A4(new_n873), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT51), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(KEYINPUT117), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT117), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n892), .A2(new_n896), .A3(new_n893), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n886), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n847), .A2(new_n853), .A3(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT118), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n847), .A2(new_n898), .A3(KEYINPUT118), .A4(new_n853), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n571), .A2(new_n312), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n782), .B1(new_n901), .B2(new_n904), .ZN(G75));
  AOI21_X1  g719(.A(new_n267), .B1(new_n832), .B2(new_n844), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n452), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT120), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT56), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n455), .B(new_n440), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT55), .Z(new_n911));
  INV_X1    g725(.A(KEYINPUT120), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n906), .A2(new_n912), .A3(new_n452), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n908), .A2(new_n909), .A3(new_n911), .A4(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n312), .A2(G952), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT119), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT56), .B1(new_n907), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n906), .A2(KEYINPUT119), .A3(new_n452), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n911), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n917), .A2(new_n921), .ZN(G51));
  INV_X1    g736(.A(new_n844), .ZN(new_n923));
  OAI21_X1  g737(.A(KEYINPUT54), .B1(new_n850), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n924), .A2(KEYINPUT121), .A3(new_n845), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT121), .ZN(new_n926));
  OAI211_X1 g740(.A(new_n926), .B(KEYINPUT54), .C1(new_n850), .C2(new_n923), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n500), .B(KEYINPUT57), .Z(new_n928));
  NAND3_X1  g742(.A1(new_n925), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT122), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n925), .A2(KEYINPUT122), .A3(new_n927), .A4(new_n928), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n931), .A2(new_n497), .A3(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n759), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n906), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n915), .B1(new_n933), .B2(new_n935), .ZN(G54));
  NAND3_X1  g750(.A1(new_n906), .A2(KEYINPUT58), .A3(G475), .ZN(new_n937));
  INV_X1    g751(.A(new_n637), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n937), .A2(new_n938), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n939), .A2(new_n940), .A3(new_n915), .ZN(G60));
  OAI21_X1  g755(.A(new_n614), .B1(new_n599), .B2(new_n616), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n847), .A2(new_n853), .ZN(new_n944));
  NAND2_X1  g758(.A1(G478), .A2(G902), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT59), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n943), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  AND4_X1   g761(.A1(new_n943), .A2(new_n925), .A3(new_n927), .A4(new_n946), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n947), .A2(new_n915), .A3(new_n948), .ZN(G63));
  NAND2_X1  g763(.A1(G217), .A2(G902), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT60), .Z(new_n951));
  OAI211_X1 g765(.A(new_n647), .B(new_n951), .C1(new_n850), .C2(new_n923), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n916), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT123), .ZN(new_n954));
  OAI21_X1  g768(.A(KEYINPUT61), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n832), .A2(new_n844), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n365), .B1(new_n956), .B2(new_n951), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n957), .A2(new_n953), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n955), .B(new_n958), .Z(G66));
  OAI21_X1  g773(.A(G953), .B1(new_n577), .B2(new_n375), .ZN(new_n960));
  INV_X1    g774(.A(new_n796), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n960), .B1(new_n961), .B2(G953), .ZN(new_n962));
  INV_X1    g776(.A(G898), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n455), .B1(new_n963), .B2(G953), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n962), .B(new_n964), .Z(G69));
  NOR2_X1   g779(.A1(new_n545), .A2(new_n546), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n288), .B(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  OAI211_X1 g782(.A(G900), .B(G953), .C1(new_n968), .C2(G227), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(G227), .B2(new_n968), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n670), .A2(new_n784), .A3(new_n688), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n684), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n776), .B1(KEYINPUT62), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(KEYINPUT62), .ZN(new_n974));
  OR2_X1    g788(.A1(new_n974), .A2(KEYINPUT124), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(KEYINPUT124), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n682), .A2(new_n728), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n690), .A2(new_n793), .A3(new_n978), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n768), .A2(KEYINPUT125), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(KEYINPUT125), .B1(new_n768), .B2(new_n979), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n977), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n967), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n767), .A2(new_n799), .A3(new_n785), .ZN(new_n984));
  AND4_X1   g798(.A1(new_n743), .A2(new_n984), .A3(new_n745), .A4(new_n971), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n768), .A2(new_n985), .A3(new_n776), .ZN(new_n986));
  AOI21_X1  g800(.A(G953), .B1(new_n986), .B2(new_n968), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n970), .B1(new_n983), .B2(new_n987), .ZN(G72));
  OAI211_X1 g802(.A(new_n961), .B(new_n977), .C1(new_n980), .C2(new_n981), .ZN(new_n989));
  NAND2_X1  g803(.A1(G472), .A2(G902), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT63), .Z(new_n991));
  NAND2_X1  g805(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n250), .B(KEYINPUT126), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n992), .A2(new_n255), .A3(new_n993), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n768), .A2(new_n985), .A3(new_n776), .A4(new_n961), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n995), .A2(new_n991), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n993), .A2(new_n255), .ZN(new_n997));
  INV_X1    g811(.A(new_n997), .ZN(new_n998));
  OAI211_X1 g812(.A(KEYINPUT127), .B(new_n916), .C1(new_n996), .C2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT127), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n998), .B1(new_n995), .B2(new_n991), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n1000), .B1(new_n1001), .B2(new_n915), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n257), .A2(new_n303), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n991), .B(new_n1004), .C1(new_n848), .C2(new_n850), .ZN(new_n1005));
  AND3_X1   g819(.A1(new_n994), .A2(new_n1003), .A3(new_n1005), .ZN(G57));
endmodule


