

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717;

  NAND2_X1 U368 ( .A1(n537), .A2(n538), .ZN(n540) );
  NOR2_X1 U369 ( .A1(n717), .A2(n716), .ZN(n568) );
  AND2_X1 U370 ( .A1(n533), .A2(n375), .ZN(n534) );
  XNOR2_X1 U371 ( .A(n376), .B(KEYINPUT35), .ZN(n533) );
  XNOR2_X1 U372 ( .A(n362), .B(n515), .ZN(n535) );
  NAND2_X1 U373 ( .A1(n610), .A2(n378), .ZN(n362) );
  NOR2_X1 U374 ( .A1(n570), .A2(n560), .ZN(n551) );
  XNOR2_X1 U375 ( .A(n504), .B(n505), .ZN(n506) );
  NOR2_X1 U376 ( .A1(n531), .A2(n556), .ZN(n513) );
  OR2_X1 U377 ( .A1(n674), .A2(G902), .ZN(n374) );
  XNOR2_X1 U378 ( .A(n377), .B(G128), .ZN(n372) );
  XNOR2_X1 U379 ( .A(n365), .B(G104), .ZN(n458) );
  INV_X1 U380 ( .A(G122), .ZN(n365) );
  INV_X1 U381 ( .A(G953), .ZN(n706) );
  OR2_X2 U382 ( .A1(n667), .A2(n353), .ZN(n672) );
  XNOR2_X1 U383 ( .A(n546), .B(KEYINPUT80), .ZN(n549) );
  XNOR2_X1 U384 ( .A(n462), .B(n424), .ZN(n704) );
  XNOR2_X1 U385 ( .A(n567), .B(KEYINPUT40), .ZN(n716) );
  AND2_X2 U386 ( .A1(n385), .A2(n666), .ZN(n371) );
  XOR2_X2 U387 ( .A(KEYINPUT68), .B(G131), .Z(n441) );
  XNOR2_X2 U388 ( .A(n540), .B(n539), .ZN(n698) );
  NOR2_X1 U389 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U390 ( .A(n691), .B(n358), .ZN(n668) );
  XNOR2_X1 U391 ( .A(n416), .B(n461), .ZN(n691) );
  XNOR2_X1 U392 ( .A(n403), .B(n427), .ZN(n461) );
  XNOR2_X1 U393 ( .A(n428), .B(KEYINPUT73), .ZN(n403) );
  XNOR2_X1 U394 ( .A(n372), .B(n422), .ZN(n462) );
  XNOR2_X1 U395 ( .A(n393), .B(KEYINPUT15), .ZN(n666) );
  XNOR2_X1 U396 ( .A(G146), .B(G125), .ZN(n463) );
  INV_X2 U397 ( .A(n410), .ZN(n686) );
  XNOR2_X2 U398 ( .A(n469), .B(KEYINPUT19), .ZN(n581) );
  NOR2_X1 U399 ( .A1(G953), .A2(G237), .ZN(n434) );
  INV_X1 U400 ( .A(G143), .ZN(n377) );
  XNOR2_X1 U401 ( .A(n704), .B(n425), .ZN(n481) );
  INV_X1 U402 ( .A(G146), .ZN(n425) );
  XNOR2_X1 U403 ( .A(n464), .B(KEYINPUT84), .ZN(n465) );
  INV_X1 U404 ( .A(n426), .ZN(n428) );
  INV_X1 U405 ( .A(KEYINPUT1), .ZN(n373) );
  OR2_X1 U406 ( .A1(n543), .A2(n352), .ZN(n544) );
  AND2_X1 U407 ( .A1(n603), .A2(n529), .ZN(n360) );
  AND2_X1 U408 ( .A1(n392), .A2(n647), .ZN(n593) );
  XNOR2_X1 U409 ( .A(n461), .B(n402), .ZN(n433) );
  XNOR2_X1 U410 ( .A(n431), .B(n432), .ZN(n402) );
  INV_X1 U411 ( .A(G110), .ZN(n364) );
  XNOR2_X1 U412 ( .A(n481), .B(n482), .ZN(n674) );
  XNOR2_X1 U413 ( .A(n414), .B(n462), .ZN(n358) );
  XNOR2_X1 U414 ( .A(n415), .B(n421), .ZN(n414) );
  NAND2_X1 U415 ( .A1(n367), .A2(n366), .ZN(n385) );
  AND2_X1 U416 ( .A1(n350), .A2(n398), .ZN(n366) );
  XNOR2_X1 U417 ( .A(n380), .B(n379), .ZN(n413) );
  INV_X1 U418 ( .A(KEYINPUT82), .ZN(n379) );
  XNOR2_X1 U419 ( .A(n632), .B(n404), .ZN(n556) );
  INV_X1 U420 ( .A(KEYINPUT106), .ZN(n404) );
  NAND2_X2 U421 ( .A1(n371), .A2(n386), .ZN(n410) );
  NOR2_X1 U422 ( .A1(n410), .A2(n409), .ZN(n408) );
  INV_X1 U423 ( .A(G475), .ZN(n409) );
  XNOR2_X1 U424 ( .A(n679), .B(n407), .ZN(n406) );
  INV_X1 U425 ( .A(KEYINPUT59), .ZN(n407) );
  INV_X1 U426 ( .A(KEYINPUT44), .ZN(n375) );
  OR2_X1 U427 ( .A1(G237), .A2(G902), .ZN(n467) );
  XNOR2_X1 U428 ( .A(G137), .B(G116), .ZN(n429) );
  XOR2_X1 U429 ( .A(KEYINPUT5), .B(KEYINPUT79), .Z(n430) );
  XNOR2_X1 U430 ( .A(G119), .B(G113), .ZN(n426) );
  XNOR2_X1 U431 ( .A(G113), .B(G143), .ZN(n437) );
  XOR2_X1 U432 ( .A(KEYINPUT11), .B(G140), .Z(n438) );
  XOR2_X1 U433 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n436) );
  XNOR2_X1 U434 ( .A(n463), .B(KEYINPUT10), .ZN(n495) );
  XNOR2_X1 U435 ( .A(G101), .B(G104), .ZN(n476) );
  XOR2_X1 U436 ( .A(G110), .B(G107), .Z(n477) );
  XOR2_X1 U437 ( .A(G137), .B(G140), .Z(n496) );
  XNOR2_X1 U438 ( .A(n471), .B(n370), .ZN(n473) );
  XOR2_X1 U439 ( .A(KEYINPUT93), .B(KEYINPUT14), .Z(n471) );
  XNOR2_X1 U440 ( .A(n470), .B(KEYINPUT78), .ZN(n370) );
  NAND2_X1 U441 ( .A1(G234), .A2(G237), .ZN(n470) );
  XNOR2_X1 U442 ( .A(n355), .B(n592), .ZN(n398) );
  INV_X1 U443 ( .A(KEYINPUT70), .ZN(n368) );
  AND2_X1 U444 ( .A1(n530), .A2(n360), .ZN(n538) );
  XNOR2_X1 U445 ( .A(KEYINPUT67), .B(KEYINPUT8), .ZN(n450) );
  XNOR2_X1 U446 ( .A(G122), .B(KEYINPUT7), .ZN(n447) );
  XNOR2_X1 U447 ( .A(KEYINPUT91), .B(G902), .ZN(n393) );
  AND2_X1 U448 ( .A1(n556), .A2(n647), .ZN(n547) );
  XNOR2_X1 U449 ( .A(n457), .B(n456), .ZN(n525) );
  XNOR2_X1 U450 ( .A(G478), .B(KEYINPUT102), .ZN(n456) );
  OR2_X1 U451 ( .A1(n500), .A2(G902), .ZN(n405) );
  OR2_X1 U452 ( .A1(n688), .A2(G902), .ZN(n384) );
  XNOR2_X1 U453 ( .A(n460), .B(n459), .ZN(n416) );
  XNOR2_X1 U454 ( .A(n458), .B(n363), .ZN(n460) );
  XNOR2_X1 U455 ( .A(n364), .B(KEYINPUT16), .ZN(n363) );
  INV_X1 U456 ( .A(G478), .ZN(n396) );
  XNOR2_X1 U457 ( .A(n595), .B(n369), .ZN(n597) );
  XNOR2_X1 U458 ( .A(KEYINPUT43), .B(KEYINPUT110), .ZN(n369) );
  NAND2_X1 U459 ( .A1(n579), .A2(n578), .ZN(n625) );
  XNOR2_X1 U460 ( .A(n391), .B(n577), .ZN(n578) );
  XNOR2_X1 U461 ( .A(n412), .B(n411), .ZN(n378) );
  XNOR2_X1 U462 ( .A(n511), .B(KEYINPUT81), .ZN(n411) );
  XNOR2_X1 U463 ( .A(n395), .B(n394), .ZN(n685) );
  XNOR2_X1 U464 ( .A(n684), .B(KEYINPUT123), .ZN(n394) );
  NOR2_X1 U465 ( .A1(n410), .A2(n396), .ZN(n395) );
  XNOR2_X1 U466 ( .A(n408), .B(n406), .ZN(n681) );
  XNOR2_X1 U467 ( .A(n675), .B(n676), .ZN(n418) );
  INV_X1 U468 ( .A(KEYINPUT56), .ZN(n356) );
  NAND2_X1 U469 ( .A1(n673), .A2(n680), .ZN(n357) );
  XNOR2_X1 U470 ( .A(n672), .B(n671), .ZN(n673) );
  XOR2_X1 U471 ( .A(n499), .B(KEYINPUT25), .Z(n346) );
  INV_X1 U472 ( .A(n628), .ZN(n514) );
  XOR2_X1 U473 ( .A(G472), .B(KEYINPUT76), .Z(n347) );
  XOR2_X1 U474 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n348) );
  XOR2_X1 U475 ( .A(KEYINPUT87), .B(n535), .Z(n349) );
  AND2_X1 U476 ( .A1(n390), .A2(KEYINPUT2), .ZN(n350) );
  XOR2_X1 U477 ( .A(n483), .B(G469), .Z(n351) );
  AND2_X1 U478 ( .A1(n542), .A2(G953), .ZN(n352) );
  NAND2_X1 U479 ( .A1(n666), .A2(G210), .ZN(n353) );
  NAND2_X1 U480 ( .A1(n354), .A2(n680), .ZN(n361) );
  XNOR2_X1 U481 ( .A(n599), .B(n600), .ZN(n354) );
  XNOR2_X1 U482 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U483 ( .A(n555), .B(n368), .ZN(n573) );
  NAND2_X1 U484 ( .A1(n399), .A2(n400), .ZN(n355) );
  NAND2_X1 U485 ( .A1(n705), .A2(n389), .ZN(n387) );
  XNOR2_X1 U486 ( .A(n492), .B(n491), .ZN(n494) );
  XNOR2_X1 U487 ( .A(n357), .B(n356), .ZN(G51) );
  NAND2_X1 U488 ( .A1(n628), .A2(n629), .ZN(n633) );
  XNOR2_X2 U489 ( .A(n384), .B(n346), .ZN(n628) );
  XNOR2_X1 U490 ( .A(n534), .B(KEYINPUT66), .ZN(n536) );
  XNOR2_X1 U491 ( .A(n348), .B(n463), .ZN(n415) );
  NAND2_X1 U492 ( .A1(n417), .A2(n680), .ZN(n677) );
  XNOR2_X2 U493 ( .A(n359), .B(KEYINPUT0), .ZN(n519) );
  NOR2_X2 U494 ( .A1(n581), .A2(n475), .ZN(n359) );
  AND2_X2 U495 ( .A1(n550), .A2(n647), .ZN(n469) );
  AND2_X2 U496 ( .A1(n509), .A2(n519), .ZN(n510) );
  XNOR2_X1 U497 ( .A(n361), .B(n602), .ZN(G57) );
  INV_X1 U498 ( .A(n698), .ZN(n367) );
  XNOR2_X1 U499 ( .A(n419), .B(n418), .ZN(n417) );
  NAND2_X1 U500 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U501 ( .A1(n657), .A2(G953), .ZN(n543) );
  XNOR2_X1 U502 ( .A(n372), .B(n447), .ZN(n448) );
  XNOR2_X2 U503 ( .A(n558), .B(n373), .ZN(n634) );
  XNOR2_X2 U504 ( .A(n374), .B(n351), .ZN(n558) );
  INV_X1 U505 ( .A(n533), .ZN(n715) );
  NOR2_X2 U506 ( .A1(n506), .A2(n569), .ZN(n376) );
  XNOR2_X1 U507 ( .A(n378), .B(G119), .ZN(G21) );
  NAND2_X1 U508 ( .A1(n386), .A2(n385), .ZN(n667) );
  NAND2_X1 U509 ( .A1(n382), .A2(n381), .ZN(n380) );
  NOR2_X1 U510 ( .A1(n634), .A2(n628), .ZN(n381) );
  XNOR2_X1 U511 ( .A(n572), .B(KEYINPUT83), .ZN(n382) );
  AND2_X1 U512 ( .A1(n383), .A2(n514), .ZN(n554) );
  INV_X1 U513 ( .A(n553), .ZN(n383) );
  NAND2_X1 U514 ( .A1(n698), .A2(n389), .ZN(n388) );
  AND2_X2 U515 ( .A1(n388), .A2(n387), .ZN(n386) );
  NAND2_X1 U516 ( .A1(n398), .A2(n390), .ZN(n705) );
  INV_X1 U517 ( .A(KEYINPUT2), .ZN(n389) );
  AND2_X1 U518 ( .A1(n627), .A2(n397), .ZN(n390) );
  NAND2_X1 U519 ( .A1(n593), .A2(n576), .ZN(n391) );
  XNOR2_X1 U520 ( .A(n575), .B(KEYINPUT108), .ZN(n392) );
  NAND2_X1 U521 ( .A1(n512), .A2(n413), .ZN(n412) );
  INV_X1 U522 ( .A(n626), .ZN(n397) );
  XNOR2_X1 U523 ( .A(n568), .B(KEYINPUT46), .ZN(n399) );
  XNOR2_X1 U524 ( .A(n591), .B(n401), .ZN(n400) );
  INV_X1 U525 ( .A(KEYINPUT69), .ZN(n401) );
  XNOR2_X2 U526 ( .A(n405), .B(n347), .ZN(n632) );
  XNOR2_X2 U527 ( .A(n510), .B(KEYINPUT22), .ZN(n512) );
  NAND2_X1 U528 ( .A1(n686), .A2(G469), .ZN(n419) );
  XNOR2_X1 U529 ( .A(n632), .B(KEYINPUT6), .ZN(n572) );
  AND2_X1 U530 ( .A1(G221), .A2(n493), .ZN(n420) );
  AND2_X1 U531 ( .A1(G224), .A2(n706), .ZN(n421) );
  INV_X1 U532 ( .A(KEYINPUT48), .ZN(n592) );
  XNOR2_X1 U533 ( .A(n501), .B(KEYINPUT107), .ZN(n502) );
  INV_X1 U534 ( .A(KEYINPUT74), .ZN(n489) );
  XNOR2_X1 U535 ( .A(n503), .B(n502), .ZN(n658) );
  NOR2_X1 U536 ( .A1(n526), .A2(n507), .ZN(n645) );
  XNOR2_X1 U537 ( .A(n494), .B(n420), .ZN(n497) );
  XNOR2_X1 U538 ( .A(n670), .B(n669), .ZN(n671) );
  INV_X1 U539 ( .A(KEYINPUT32), .ZN(n511) );
  XOR2_X1 U540 ( .A(KEYINPUT63), .B(KEYINPUT89), .Z(n602) );
  XNOR2_X1 U541 ( .A(KEYINPUT4), .B(KEYINPUT64), .ZN(n422) );
  XNOR2_X1 U542 ( .A(n441), .B(G134), .ZN(n423) );
  INV_X1 U543 ( .A(n423), .ZN(n424) );
  XNOR2_X1 U544 ( .A(KEYINPUT3), .B(G101), .ZN(n427) );
  XNOR2_X1 U545 ( .A(n430), .B(n429), .ZN(n431) );
  NAND2_X1 U546 ( .A1(n434), .A2(G210), .ZN(n432) );
  XNOR2_X1 U547 ( .A(n481), .B(n433), .ZN(n500) );
  XOR2_X1 U548 ( .A(n500), .B(KEYINPUT62), .Z(n600) );
  INV_X1 U549 ( .A(n666), .ZN(n598) );
  NAND2_X1 U550 ( .A1(G214), .A2(n434), .ZN(n435) );
  XNOR2_X1 U551 ( .A(n436), .B(n435), .ZN(n440) );
  XNOR2_X1 U552 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U553 ( .A(n440), .B(n439), .Z(n443) );
  XNOR2_X1 U554 ( .A(n441), .B(n458), .ZN(n442) );
  XNOR2_X1 U555 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U556 ( .A(n495), .B(n444), .ZN(n678) );
  NOR2_X1 U557 ( .A1(G902), .A2(n678), .ZN(n446) );
  XNOR2_X1 U558 ( .A(KEYINPUT13), .B(G475), .ZN(n445) );
  XNOR2_X1 U559 ( .A(n446), .B(n445), .ZN(n526) );
  XOR2_X1 U560 ( .A(G116), .B(G107), .Z(n459) );
  XNOR2_X1 U561 ( .A(G134), .B(n459), .ZN(n449) );
  XNOR2_X1 U562 ( .A(n449), .B(n448), .ZN(n455) );
  XOR2_X1 U563 ( .A(KEYINPUT9), .B(KEYINPUT101), .Z(n453) );
  NAND2_X1 U564 ( .A1(n706), .A2(G234), .ZN(n451) );
  XNOR2_X1 U565 ( .A(n451), .B(n450), .ZN(n493) );
  NAND2_X1 U566 ( .A1(G217), .A2(n493), .ZN(n452) );
  XNOR2_X1 U567 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U568 ( .A(n455), .B(n454), .ZN(n684) );
  NOR2_X1 U569 ( .A1(G902), .A2(n684), .ZN(n457) );
  INV_X1 U570 ( .A(n525), .ZN(n507) );
  NAND2_X1 U571 ( .A1(n526), .A2(n507), .ZN(n569) );
  INV_X1 U572 ( .A(KEYINPUT34), .ZN(n505) );
  NOR2_X1 U573 ( .A1(n668), .A2(n666), .ZN(n466) );
  NAND2_X1 U574 ( .A1(G210), .A2(n467), .ZN(n464) );
  XNOR2_X1 U575 ( .A(n466), .B(n465), .ZN(n550) );
  NAND2_X1 U576 ( .A1(G214), .A2(n467), .ZN(n468) );
  XNOR2_X1 U577 ( .A(KEYINPUT92), .B(n468), .ZN(n647) );
  NAND2_X1 U578 ( .A1(n473), .A2(G952), .ZN(n472) );
  XNOR2_X1 U579 ( .A(n472), .B(KEYINPUT94), .ZN(n657) );
  NAND2_X1 U580 ( .A1(G902), .A2(n473), .ZN(n541) );
  XNOR2_X1 U581 ( .A(G898), .B(KEYINPUT95), .ZN(n696) );
  NAND2_X1 U582 ( .A1(G953), .A2(n696), .ZN(n693) );
  NOR2_X1 U583 ( .A1(n541), .A2(n693), .ZN(n474) );
  NOR2_X1 U584 ( .A1(n543), .A2(n474), .ZN(n475) );
  XOR2_X1 U585 ( .A(n519), .B(KEYINPUT96), .Z(n523) );
  XNOR2_X1 U586 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U587 ( .A(n496), .B(n478), .Z(n480) );
  NAND2_X1 U588 ( .A1(G227), .A2(n706), .ZN(n479) );
  XNOR2_X1 U589 ( .A(n480), .B(n479), .ZN(n482) );
  XNOR2_X1 U590 ( .A(KEYINPUT72), .B(KEYINPUT71), .ZN(n483) );
  XOR2_X1 U591 ( .A(KEYINPUT98), .B(KEYINPUT21), .Z(n486) );
  NAND2_X1 U592 ( .A1(G234), .A2(n598), .ZN(n484) );
  XNOR2_X1 U593 ( .A(KEYINPUT20), .B(n484), .ZN(n498) );
  NAND2_X1 U594 ( .A1(n498), .A2(G221), .ZN(n485) );
  XNOR2_X1 U595 ( .A(n486), .B(n485), .ZN(n629) );
  XOR2_X1 U596 ( .A(KEYINPUT24), .B(KEYINPUT97), .Z(n488) );
  XNOR2_X1 U597 ( .A(G110), .B(KEYINPUT23), .ZN(n487) );
  XNOR2_X1 U598 ( .A(n488), .B(n487), .ZN(n492) );
  XNOR2_X1 U599 ( .A(G119), .B(G128), .ZN(n490) );
  XOR2_X1 U600 ( .A(n496), .B(n495), .Z(n703) );
  XNOR2_X1 U601 ( .A(n497), .B(n703), .ZN(n688) );
  NAND2_X1 U602 ( .A1(n498), .A2(G217), .ZN(n499) );
  NOR2_X1 U603 ( .A1(n634), .A2(n633), .ZN(n517) );
  NAND2_X1 U604 ( .A1(n517), .A2(n572), .ZN(n503) );
  XOR2_X1 U605 ( .A(KEYINPUT33), .B(KEYINPUT75), .Z(n501) );
  NOR2_X1 U606 ( .A1(n523), .A2(n658), .ZN(n504) );
  NAND2_X1 U607 ( .A1(n629), .A2(n645), .ZN(n508) );
  XNOR2_X1 U608 ( .A(KEYINPUT105), .B(n508), .ZN(n509) );
  NAND2_X1 U609 ( .A1(n634), .A2(n512), .ZN(n531) );
  NAND2_X1 U610 ( .A1(n514), .A2(n513), .ZN(n610) );
  INV_X1 U611 ( .A(KEYINPUT88), .ZN(n515) );
  NAND2_X1 U612 ( .A1(n533), .A2(n535), .ZN(n516) );
  NAND2_X1 U613 ( .A1(n516), .A2(KEYINPUT44), .ZN(n530) );
  INV_X1 U614 ( .A(n517), .ZN(n518) );
  NOR2_X1 U615 ( .A1(n632), .A2(n518), .ZN(n639) );
  NAND2_X1 U616 ( .A1(n519), .A2(n639), .ZN(n520) );
  XOR2_X1 U617 ( .A(KEYINPUT31), .B(n520), .Z(n621) );
  INV_X1 U618 ( .A(n558), .ZN(n521) );
  NOR2_X1 U619 ( .A1(n521), .A2(n633), .ZN(n522) );
  XNOR2_X1 U620 ( .A(n522), .B(KEYINPUT99), .ZN(n545) );
  NOR2_X1 U621 ( .A1(n545), .A2(n523), .ZN(n524) );
  NAND2_X1 U622 ( .A1(n632), .A2(n524), .ZN(n605) );
  NAND2_X1 U623 ( .A1(n621), .A2(n605), .ZN(n527) );
  NAND2_X1 U624 ( .A1(n526), .A2(n525), .ZN(n619) );
  NOR2_X1 U625 ( .A1(n526), .A2(n525), .ZN(n611) );
  INV_X1 U626 ( .A(n611), .ZN(n622) );
  XOR2_X1 U627 ( .A(KEYINPUT103), .B(n622), .Z(n552) );
  NAND2_X1 U628 ( .A1(n619), .A2(n552), .ZN(n642) );
  NAND2_X1 U629 ( .A1(n527), .A2(n642), .ZN(n528) );
  XNOR2_X1 U630 ( .A(n528), .B(KEYINPUT104), .ZN(n529) );
  NOR2_X1 U631 ( .A1(n572), .A2(n531), .ZN(n532) );
  NAND2_X1 U632 ( .A1(n532), .A2(n628), .ZN(n603) );
  NAND2_X1 U633 ( .A1(n536), .A2(n349), .ZN(n537) );
  XOR2_X1 U634 ( .A(KEYINPUT45), .B(KEYINPUT86), .Z(n539) );
  NOR2_X1 U635 ( .A1(G900), .A2(n541), .ZN(n542) );
  XNOR2_X1 U636 ( .A(n544), .B(KEYINPUT85), .ZN(n553) );
  NOR2_X1 U637 ( .A1(n545), .A2(n553), .ZN(n546) );
  XNOR2_X1 U638 ( .A(KEYINPUT30), .B(n547), .ZN(n548) );
  NAND2_X1 U639 ( .A1(n549), .A2(n548), .ZN(n570) );
  BUF_X1 U640 ( .A(n550), .Z(n576) );
  INV_X1 U641 ( .A(n576), .ZN(n596) );
  XOR2_X1 U642 ( .A(KEYINPUT38), .B(n596), .Z(n560) );
  XNOR2_X1 U643 ( .A(n551), .B(KEYINPUT39), .ZN(n566) );
  NOR2_X1 U644 ( .A1(n566), .A2(n552), .ZN(n626) );
  NAND2_X1 U645 ( .A1(n629), .A2(n554), .ZN(n555) );
  AND2_X1 U646 ( .A1(n573), .A2(n556), .ZN(n557) );
  XNOR2_X1 U647 ( .A(n557), .B(KEYINPUT28), .ZN(n559) );
  NAND2_X1 U648 ( .A1(n559), .A2(n558), .ZN(n582) );
  INV_X1 U649 ( .A(n560), .ZN(n646) );
  NAND2_X1 U650 ( .A1(n646), .A2(n647), .ZN(n561) );
  XNOR2_X1 U651 ( .A(n561), .B(KEYINPUT111), .ZN(n643) );
  NAND2_X1 U652 ( .A1(n643), .A2(n645), .ZN(n564) );
  XNOR2_X1 U653 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n562) );
  XNOR2_X1 U654 ( .A(n562), .B(KEYINPUT41), .ZN(n563) );
  XNOR2_X1 U655 ( .A(n564), .B(n563), .ZN(n659) );
  NOR2_X1 U656 ( .A1(n582), .A2(n659), .ZN(n565) );
  XNOR2_X1 U657 ( .A(n565), .B(KEYINPUT42), .ZN(n717) );
  NOR2_X1 U658 ( .A1(n566), .A2(n619), .ZN(n567) );
  NOR2_X1 U659 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U660 ( .A1(n571), .A2(n576), .ZN(n615) );
  INV_X1 U661 ( .A(n634), .ZN(n579) );
  XOR2_X1 U662 ( .A(KEYINPUT114), .B(KEYINPUT36), .Z(n577) );
  NOR2_X1 U663 ( .A1(n619), .A2(n574), .ZN(n575) );
  NAND2_X1 U664 ( .A1(n615), .A2(n625), .ZN(n590) );
  INV_X1 U665 ( .A(n642), .ZN(n580) );
  NOR2_X1 U666 ( .A1(n580), .A2(KEYINPUT77), .ZN(n583) );
  NOR2_X1 U667 ( .A1(n582), .A2(n581), .ZN(n616) );
  NAND2_X1 U668 ( .A1(n583), .A2(n616), .ZN(n584) );
  NAND2_X1 U669 ( .A1(n584), .A2(KEYINPUT47), .ZN(n588) );
  XNOR2_X1 U670 ( .A(KEYINPUT77), .B(n642), .ZN(n585) );
  NOR2_X1 U671 ( .A1(KEYINPUT47), .A2(n585), .ZN(n586) );
  NAND2_X1 U672 ( .A1(n586), .A2(n616), .ZN(n587) );
  NAND2_X1 U673 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U674 ( .A(n593), .B(KEYINPUT109), .Z(n594) );
  NAND2_X1 U675 ( .A1(n594), .A2(n634), .ZN(n595) );
  NAND2_X1 U676 ( .A1(n597), .A2(n596), .ZN(n627) );
  NAND2_X1 U677 ( .A1(G472), .A2(n686), .ZN(n599) );
  NOR2_X1 U678 ( .A1(G952), .A2(n706), .ZN(n601) );
  XNOR2_X1 U679 ( .A(KEYINPUT90), .B(n601), .ZN(n690) );
  INV_X1 U680 ( .A(n690), .ZN(n680) );
  XNOR2_X1 U681 ( .A(G101), .B(n603), .ZN(G3) );
  NOR2_X1 U682 ( .A1(n619), .A2(n605), .ZN(n604) );
  XOR2_X1 U683 ( .A(G104), .B(n604), .Z(G6) );
  NOR2_X1 U684 ( .A1(n622), .A2(n605), .ZN(n607) );
  XNOR2_X1 U685 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n606) );
  XNOR2_X1 U686 ( .A(n607), .B(n606), .ZN(n608) );
  XNOR2_X1 U687 ( .A(G107), .B(n608), .ZN(G9) );
  XOR2_X1 U688 ( .A(G110), .B(KEYINPUT115), .Z(n609) );
  XNOR2_X1 U689 ( .A(n610), .B(n609), .ZN(G12) );
  XOR2_X1 U690 ( .A(KEYINPUT29), .B(KEYINPUT116), .Z(n613) );
  NAND2_X1 U691 ( .A1(n616), .A2(n611), .ZN(n612) );
  XNOR2_X1 U692 ( .A(n613), .B(n612), .ZN(n614) );
  XNOR2_X1 U693 ( .A(G128), .B(n614), .ZN(G30) );
  XNOR2_X1 U694 ( .A(G143), .B(n615), .ZN(G45) );
  INV_X1 U695 ( .A(n619), .ZN(n617) );
  NAND2_X1 U696 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U697 ( .A(G146), .B(n618), .ZN(G48) );
  NOR2_X1 U698 ( .A1(n619), .A2(n621), .ZN(n620) );
  XOR2_X1 U699 ( .A(G113), .B(n620), .Z(G15) );
  NOR2_X1 U700 ( .A1(n622), .A2(n621), .ZN(n623) );
  XOR2_X1 U701 ( .A(G116), .B(n623), .Z(G18) );
  XOR2_X1 U702 ( .A(G125), .B(KEYINPUT37), .Z(n624) );
  XNOR2_X1 U703 ( .A(n625), .B(n624), .ZN(G27) );
  XOR2_X1 U704 ( .A(G134), .B(n626), .Z(G36) );
  XNOR2_X1 U705 ( .A(G140), .B(n627), .ZN(G42) );
  NOR2_X1 U706 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U707 ( .A(n630), .B(KEYINPUT49), .ZN(n631) );
  NAND2_X1 U708 ( .A1(n632), .A2(n631), .ZN(n637) );
  NAND2_X1 U709 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U710 ( .A(KEYINPUT50), .B(n635), .Z(n636) );
  NOR2_X1 U711 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U712 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U713 ( .A(KEYINPUT51), .B(n640), .Z(n641) );
  NOR2_X1 U714 ( .A1(n659), .A2(n641), .ZN(n654) );
  NAND2_X1 U715 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U716 ( .A(KEYINPUT117), .B(n644), .ZN(n651) );
  INV_X1 U717 ( .A(n645), .ZN(n649) );
  NOR2_X1 U718 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U719 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U720 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U721 ( .A1(n652), .A2(n658), .ZN(n653) );
  NOR2_X1 U722 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U723 ( .A(n655), .B(KEYINPUT52), .ZN(n656) );
  NOR2_X1 U724 ( .A1(n657), .A2(n656), .ZN(n662) );
  NOR2_X1 U725 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U726 ( .A(KEYINPUT118), .B(n660), .ZN(n661) );
  NOR2_X1 U727 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U728 ( .A1(n663), .A2(n667), .ZN(n664) );
  NOR2_X1 U729 ( .A1(n664), .A2(G953), .ZN(n665) );
  XNOR2_X1 U730 ( .A(n665), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U731 ( .A(n668), .B(KEYINPUT55), .ZN(n670) );
  XOR2_X1 U732 ( .A(KEYINPUT54), .B(KEYINPUT119), .Z(n669) );
  XOR2_X1 U733 ( .A(n674), .B(KEYINPUT120), .Z(n675) );
  XOR2_X1 U734 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n676) );
  XNOR2_X1 U735 ( .A(n677), .B(KEYINPUT121), .ZN(G54) );
  XNOR2_X1 U736 ( .A(n678), .B(KEYINPUT122), .ZN(n679) );
  NAND2_X1 U737 ( .A1(n681), .A2(n680), .ZN(n683) );
  XNOR2_X1 U738 ( .A(KEYINPUT65), .B(KEYINPUT60), .ZN(n682) );
  XNOR2_X1 U739 ( .A(n683), .B(n682), .ZN(G60) );
  NOR2_X1 U740 ( .A1(n690), .A2(n685), .ZN(G63) );
  NAND2_X1 U741 ( .A1(G217), .A2(n686), .ZN(n687) );
  XNOR2_X1 U742 ( .A(n688), .B(n687), .ZN(n689) );
  NOR2_X1 U743 ( .A1(n690), .A2(n689), .ZN(G66) );
  XOR2_X1 U744 ( .A(n691), .B(KEYINPUT125), .Z(n692) );
  NAND2_X1 U745 ( .A1(n693), .A2(n692), .ZN(n702) );
  XOR2_X1 U746 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n695) );
  NAND2_X1 U747 ( .A1(G224), .A2(G953), .ZN(n694) );
  XNOR2_X1 U748 ( .A(n695), .B(n694), .ZN(n697) );
  NOR2_X1 U749 ( .A1(n697), .A2(n696), .ZN(n700) );
  NOR2_X1 U750 ( .A1(G953), .A2(n698), .ZN(n699) );
  NOR2_X1 U751 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U752 ( .A(n702), .B(n701), .ZN(G69) );
  XOR2_X1 U753 ( .A(n704), .B(n703), .Z(n709) );
  XOR2_X1 U754 ( .A(n709), .B(n705), .Z(n707) );
  NAND2_X1 U755 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U756 ( .A(n708), .B(KEYINPUT126), .ZN(n714) );
  XNOR2_X1 U757 ( .A(n709), .B(G227), .ZN(n710) );
  XNOR2_X1 U758 ( .A(n710), .B(KEYINPUT127), .ZN(n711) );
  NAND2_X1 U759 ( .A1(n711), .A2(G900), .ZN(n712) );
  NAND2_X1 U760 ( .A1(G953), .A2(n712), .ZN(n713) );
  NAND2_X1 U761 ( .A1(n714), .A2(n713), .ZN(G72) );
  XOR2_X1 U762 ( .A(G122), .B(n715), .Z(G24) );
  XOR2_X1 U763 ( .A(n716), .B(G131), .Z(G33) );
  XOR2_X1 U764 ( .A(G137), .B(n717), .Z(G39) );
endmodule

