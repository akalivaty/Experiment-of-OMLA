//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1 0 1 1 1 0 1 0 0 0 1 0 0 1 1 0 1 1 1 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  OR2_X1    g003(.A1(KEYINPUT72), .A2(G125), .ZN(new_n190));
  NAND2_X1  g004(.A1(KEYINPUT72), .A2(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  OR3_X1    g006(.A1(new_n192), .A2(KEYINPUT16), .A3(G140), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT73), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n190), .A2(G140), .A3(new_n191), .ZN(new_n195));
  OR2_X1    g009(.A1(G125), .A2(G140), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n194), .B1(new_n197), .B2(KEYINPUT16), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT16), .ZN(new_n199));
  AOI211_X1 g013(.A(KEYINPUT73), .B(new_n199), .C1(new_n195), .C2(new_n196), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n193), .B1(new_n198), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  OAI211_X1 g017(.A(G146), .B(new_n193), .C1(new_n198), .C2(new_n200), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G119), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(G128), .ZN(new_n207));
  OR2_X1    g021(.A1(new_n207), .A2(KEYINPUT23), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(KEYINPUT23), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n208), .B(new_n209), .C1(G119), .C2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G110), .ZN(new_n212));
  XOR2_X1   g026(.A(KEYINPUT24), .B(G110), .Z(new_n213));
  XNOR2_X1  g027(.A(G119), .B(G128), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n205), .A2(new_n212), .A3(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(G125), .B(G140), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(new_n202), .ZN(new_n218));
  OAI22_X1  g032(.A1(new_n211), .A2(G110), .B1(new_n214), .B2(new_n213), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n204), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G953), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(G221), .A3(G234), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n222), .B(KEYINPUT22), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n223), .B(G137), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n216), .A2(new_n220), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n224), .B1(new_n216), .B2(new_n220), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(KEYINPUT25), .B1(new_n227), .B2(new_n188), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT25), .ZN(new_n229));
  NOR4_X1   g043(.A1(new_n225), .A2(new_n226), .A3(new_n229), .A4(G902), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n189), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT74), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI211_X1 g047(.A(KEYINPUT74), .B(new_n189), .C1(new_n228), .C2(new_n230), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n189), .A2(G902), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n227), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n233), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G472), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT66), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n202), .A2(G143), .ZN(new_n240));
  AND2_X1   g054(.A1(KEYINPUT64), .A2(G143), .ZN(new_n241));
  NOR2_X1   g055(.A1(KEYINPUT64), .A2(G143), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n240), .B1(new_n243), .B2(new_n202), .ZN(new_n244));
  INV_X1    g058(.A(G143), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT1), .B1(new_n245), .B2(G146), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G128), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n239), .B1(new_n244), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(G146), .B1(new_n241), .B2(new_n242), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT1), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n202), .A2(G143), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n250), .A2(new_n251), .A3(G128), .A4(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT64), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(new_n245), .ZN(new_n255));
  NAND2_X1  g069(.A1(KEYINPUT64), .A2(G143), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n255), .A2(new_n202), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n240), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(KEYINPUT66), .A3(new_n247), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n249), .A2(new_n253), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G137), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT65), .B1(new_n262), .B2(G134), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT65), .ZN(new_n264));
  INV_X1    g078(.A(G134), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n264), .A2(new_n265), .A3(G137), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT11), .B1(new_n265), .B2(G137), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT11), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(new_n262), .A3(G134), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G131), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n267), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n265), .A2(G137), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n262), .A2(G134), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n272), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n261), .A2(new_n277), .ZN(new_n278));
  AND4_X1   g092(.A1(KEYINPUT0), .A2(new_n250), .A3(G128), .A4(new_n252), .ZN(new_n279));
  XNOR2_X1  g093(.A(KEYINPUT0), .B(G128), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n280), .B1(new_n257), .B2(new_n258), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n267), .A2(new_n271), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G131), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n267), .A2(new_n271), .A3(new_n272), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT30), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n278), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n278), .A2(KEYINPUT68), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT67), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n272), .B1(new_n267), .B2(new_n271), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n291), .B1(new_n273), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n284), .A2(KEYINPUT67), .A3(new_n285), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(new_n294), .A3(new_n282), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT68), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n261), .A2(new_n296), .A3(new_n277), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n290), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n289), .B1(new_n298), .B2(KEYINPUT30), .ZN(new_n299));
  XNOR2_X1  g113(.A(G116), .B(G119), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT2), .B(G113), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n300), .B(new_n301), .ZN(new_n302));
  OR2_X1    g116(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n290), .A2(new_n302), .A3(new_n295), .A4(new_n297), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G237), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n306), .A2(new_n221), .A3(G210), .ZN(new_n307));
  XOR2_X1   g121(.A(new_n307), .B(KEYINPUT27), .Z(new_n308));
  XNOR2_X1  g122(.A(new_n308), .B(KEYINPUT26), .ZN(new_n309));
  INV_X1    g123(.A(G101), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n309), .B(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n305), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT29), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n278), .A2(new_n295), .A3(new_n302), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT28), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT69), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n315), .A2(KEYINPUT69), .A3(new_n316), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n278), .A2(new_n287), .ZN(new_n322));
  INV_X1    g136(.A(new_n302), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n316), .B1(new_n304), .B2(new_n324), .ZN(new_n325));
  OR3_X1    g139(.A1(new_n321), .A2(new_n325), .A3(new_n312), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n313), .A2(new_n314), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n298), .A2(new_n323), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n304), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n321), .B1(KEYINPUT28), .B2(new_n329), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n312), .A2(new_n314), .ZN(new_n331));
  AOI21_X1  g145(.A(G902), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n238), .B1(new_n327), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(G472), .A2(G902), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n312), .B1(new_n321), .B2(new_n325), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n304), .B(new_n311), .C1(new_n299), .C2(new_n302), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n336), .B1(new_n337), .B2(KEYINPUT31), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n337), .A2(KEYINPUT31), .ZN(new_n339));
  OAI211_X1 g153(.A(KEYINPUT32), .B(new_n335), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT70), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT31), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n303), .A2(new_n342), .A3(new_n304), .A4(new_n311), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n337), .A2(KEYINPUT31), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n344), .A3(new_n336), .ZN(new_n345));
  AOI21_X1  g159(.A(KEYINPUT32), .B1(new_n345), .B2(new_n335), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n341), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n335), .B1(new_n338), .B2(new_n339), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT70), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT32), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n334), .B1(new_n347), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT71), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n348), .A2(new_n350), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(KEYINPUT70), .A3(new_n340), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n351), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT71), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n358), .A3(new_n334), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n237), .B1(new_n354), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(KEYINPUT75), .A2(G104), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT3), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n364));
  NOR2_X1   g178(.A1(KEYINPUT76), .A2(G107), .ZN(new_n365));
  AND2_X1   g179(.A1(KEYINPUT76), .A2(G107), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n363), .B(new_n364), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G107), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(G104), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(G104), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n369), .B1(KEYINPUT3), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n310), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT78), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT4), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n373), .B1(new_n372), .B2(new_n374), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT77), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n367), .A2(new_n371), .A3(new_n310), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n379), .A2(new_n372), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n378), .B1(new_n380), .B2(KEYINPUT4), .ZN(new_n381));
  NOR4_X1   g195(.A1(new_n379), .A2(new_n372), .A3(KEYINPUT77), .A4(new_n374), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n282), .B(new_n377), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT79), .ZN(new_n384));
  INV_X1    g198(.A(new_n370), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n366), .A2(new_n365), .ZN(new_n386));
  INV_X1    g200(.A(G104), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT80), .B1(new_n388), .B2(new_n310), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n367), .A2(new_n371), .A3(new_n310), .ZN(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT76), .B(G107), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n370), .B1(new_n391), .B2(G104), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT80), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n393), .A3(G101), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n389), .A2(new_n390), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT81), .ZN(new_n397));
  OR2_X1    g211(.A1(new_n253), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n250), .A2(new_n252), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n251), .B1(new_n243), .B2(new_n202), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n399), .B1(new_n400), .B2(new_n210), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n253), .A2(new_n397), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n398), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n396), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT10), .ZN(new_n405));
  AOI221_X4 g219(.A(new_n239), .B1(new_n246), .B2(G128), .C1(new_n257), .C2(new_n258), .ZN(new_n406));
  AOI21_X1  g220(.A(KEYINPUT66), .B1(new_n259), .B2(new_n247), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n405), .B1(new_n408), .B2(new_n253), .ZN(new_n409));
  AOI22_X1  g223(.A1(new_n404), .A2(new_n405), .B1(new_n409), .B2(new_n396), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n380), .A2(new_n378), .A3(KEYINPUT4), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n367), .A2(new_n371), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G101), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(KEYINPUT4), .A3(new_n390), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT77), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT79), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n416), .A2(new_n417), .A3(new_n282), .A4(new_n377), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n384), .A2(new_n410), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n293), .A2(new_n294), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  AND2_X1   g236(.A1(new_n384), .A2(new_n418), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n423), .A2(KEYINPUT82), .A3(new_n420), .A4(new_n410), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n384), .A2(new_n420), .A3(new_n410), .A4(new_n418), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT82), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n422), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(G110), .B(G140), .ZN(new_n429));
  INV_X1    g243(.A(G227), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(G953), .ZN(new_n431));
  XOR2_X1   g245(.A(new_n429), .B(new_n431), .Z(new_n432));
  OAI21_X1  g246(.A(KEYINPUT83), .B1(new_n428), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n424), .A2(new_n427), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n404), .B1(new_n261), .B2(new_n396), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT12), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n436), .A3(new_n421), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n435), .A2(new_n286), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT12), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n434), .A2(new_n432), .A3(new_n437), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n419), .A2(new_n421), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n425), .A2(new_n426), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n425), .A2(new_n426), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT83), .ZN(new_n445));
  INV_X1    g259(.A(new_n432), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n433), .A2(new_n440), .A3(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(G469), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(new_n449), .A3(new_n188), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n449), .A2(new_n188), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n437), .B(new_n439), .C1(new_n442), .C2(new_n443), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n446), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n428), .A2(new_n432), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(G469), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n450), .A2(new_n452), .A3(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(G210), .B1(G237), .B2(G902), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(G110), .B(G122), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(KEYINPUT8), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT5), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(new_n206), .A3(G116), .ZN(new_n463));
  INV_X1    g277(.A(new_n300), .ZN(new_n464));
  OAI211_X1 g278(.A(G113), .B(new_n463), .C1(new_n464), .C2(new_n462), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n465), .B1(new_n464), .B2(new_n301), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n395), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n395), .A2(new_n466), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n461), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT86), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI211_X1 g285(.A(KEYINPUT86), .B(new_n461), .C1(new_n467), .C2(new_n468), .ZN(new_n472));
  INV_X1    g286(.A(new_n192), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n473), .B1(new_n279), .B2(new_n281), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT84), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g290(.A(KEYINPUT84), .B(new_n473), .C1(new_n279), .C2(new_n281), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT85), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n408), .A2(new_n479), .A3(new_n253), .A4(new_n192), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n249), .A2(new_n253), .A3(new_n260), .A4(new_n192), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT85), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n478), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n221), .A2(G224), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT7), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n471), .A2(new_n472), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT87), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n481), .B(new_n479), .ZN(new_n489));
  INV_X1    g303(.A(new_n474), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n488), .B(new_n485), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n490), .B1(new_n480), .B2(new_n482), .ZN(new_n492));
  OAI21_X1  g306(.A(KEYINPUT87), .B1(new_n492), .B2(new_n486), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT88), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n487), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n495), .B1(new_n487), .B2(new_n494), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n416), .A2(new_n323), .A3(new_n377), .ZN(new_n498));
  INV_X1    g312(.A(new_n468), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n460), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NOR3_X1   g315(.A1(new_n496), .A2(new_n497), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n498), .A2(new_n499), .ZN(new_n503));
  INV_X1    g317(.A(new_n460), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n505), .A2(KEYINPUT6), .A3(new_n500), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n483), .B(new_n484), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT6), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n503), .A2(new_n508), .A3(new_n504), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n506), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n188), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n459), .B1(new_n502), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n487), .A2(new_n494), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT88), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n487), .A2(new_n494), .A3(new_n495), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n500), .A3(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n516), .A2(new_n188), .A3(new_n458), .A4(new_n510), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n512), .A2(KEYINPUT89), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT89), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n519), .B(new_n459), .C1(new_n502), .C2(new_n511), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n221), .A2(G952), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n521), .B1(G234), .B2(G237), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  XOR2_X1   g337(.A(KEYINPUT21), .B(G898), .Z(new_n524));
  NAND2_X1  g338(.A1(G234), .A2(G237), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(G902), .A3(G953), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n523), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(G214), .B1(G237), .B2(G902), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n518), .A2(new_n520), .A3(new_n531), .ZN(new_n532));
  XOR2_X1   g346(.A(KEYINPUT9), .B(G234), .Z(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(G221), .B1(new_n534), .B2(G902), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n245), .A2(new_n306), .A3(new_n221), .A4(G214), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n255), .A2(new_n256), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n306), .A2(new_n221), .A3(G214), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT18), .ZN(new_n540));
  NOR3_X1   g354(.A1(new_n539), .A2(new_n540), .A3(new_n272), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n541), .B1(new_n272), .B2(new_n539), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n539), .A2(new_n540), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT90), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n544), .B(new_n218), .C1(new_n197), .C2(new_n202), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n195), .A2(KEYINPUT90), .A3(G146), .A4(new_n196), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n542), .A2(new_n543), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(G113), .B(G122), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(new_n387), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT92), .B1(new_n539), .B2(new_n272), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n306), .A2(new_n221), .A3(G214), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n243), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT92), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n552), .A2(new_n553), .A3(G131), .A4(new_n536), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT17), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n539), .A2(new_n272), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT91), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT91), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n539), .A2(new_n559), .A3(new_n272), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n558), .A2(new_n550), .A3(new_n554), .A4(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n556), .B1(new_n561), .B2(KEYINPUT17), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n547), .B(new_n549), .C1(new_n562), .C2(new_n205), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT94), .ZN(new_n564));
  INV_X1    g378(.A(new_n555), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT17), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n565), .A2(new_n566), .A3(new_n558), .A4(new_n560), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n567), .A2(new_n203), .A3(new_n204), .A4(new_n556), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT94), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n568), .A2(new_n569), .A3(new_n549), .A4(new_n547), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n564), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT19), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n217), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n573), .B1(new_n197), .B2(new_n572), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n574), .A2(G146), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT93), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n577), .A2(new_n204), .A3(new_n561), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n547), .ZN(new_n579));
  INV_X1    g393(.A(new_n549), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n571), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(G475), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n583), .A3(new_n188), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT20), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n549), .B1(new_n568), .B2(new_n547), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n587), .B1(new_n564), .B2(new_n570), .ZN(new_n588));
  OAI21_X1  g402(.A(G475), .B1(new_n588), .B2(G902), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n582), .A2(KEYINPUT20), .A3(new_n583), .A4(new_n188), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n586), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT15), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(G478), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT96), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT13), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n537), .A2(new_n595), .A3(G128), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n245), .A2(G128), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n598), .B1(new_n243), .B2(new_n210), .ZN(new_n599));
  OAI211_X1 g413(.A(G134), .B(new_n596), .C1(new_n599), .C2(new_n595), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n265), .B(new_n598), .C1(new_n243), .C2(new_n210), .ZN(new_n601));
  INV_X1    g415(.A(G116), .ZN(new_n602));
  OR2_X1    g416(.A1(new_n602), .A2(G122), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(G122), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n386), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n391), .A2(new_n604), .A3(new_n603), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n600), .A2(new_n601), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT95), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n600), .A2(KEYINPUT95), .A3(new_n601), .A4(new_n608), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n607), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n599), .A2(G134), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n614), .B1(new_n615), .B2(new_n601), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n604), .A2(KEYINPUT14), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n603), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n604), .A2(KEYINPUT14), .ZN(new_n619));
  OAI21_X1  g433(.A(G107), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n613), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n533), .A2(G217), .A3(new_n221), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n623), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n613), .A2(new_n621), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n594), .B1(new_n627), .B2(new_n188), .ZN(new_n628));
  AOI221_X4 g442(.A(new_n623), .B1(new_n620), .B2(new_n616), .C1(new_n611), .C2(new_n612), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n625), .B1(new_n613), .B2(new_n621), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n594), .B(new_n188), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n593), .B1(new_n628), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n631), .A2(new_n592), .A3(G478), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n591), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n457), .A2(new_n532), .A3(new_n535), .A4(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n360), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G101), .ZN(G3));
  INV_X1    g454(.A(new_n237), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n345), .A2(new_n188), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(G472), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n348), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n457), .A2(new_n641), .A3(new_n535), .A4(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n512), .A2(new_n517), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(new_n527), .A3(new_n529), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n627), .B(KEYINPUT33), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n650), .A2(G478), .A3(new_n188), .ZN(new_n651));
  INV_X1    g465(.A(G478), .ZN(new_n652));
  INV_X1    g466(.A(new_n627), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n652), .B1(new_n653), .B2(G902), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n591), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n649), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n647), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT34), .B(G104), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G6));
  AND4_X1   g474(.A1(new_n589), .A2(new_n586), .A3(new_n590), .A4(new_n635), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n649), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n647), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT35), .B(G107), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G9));
  NAND2_X1  g480(.A1(new_n216), .A2(new_n220), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT97), .ZN(new_n668));
  INV_X1    g482(.A(new_n224), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(KEYINPUT36), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n668), .A2(new_n671), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n235), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n233), .A2(new_n234), .A3(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(new_n644), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n637), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT37), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G110), .ZN(G12));
  NAND2_X1  g495(.A1(new_n354), .A2(new_n359), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n457), .A2(new_n535), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n522), .B(KEYINPUT98), .Z(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n686), .B1(G900), .B2(new_n526), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n661), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT99), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n648), .A2(new_n675), .A3(new_n529), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n682), .A2(new_n684), .A3(new_n690), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G128), .ZN(G30));
  NAND2_X1  g507(.A1(new_n518), .A2(new_n520), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(KEYINPUT100), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT38), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n696), .A2(new_n675), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n329), .A2(new_n312), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT101), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n329), .A2(KEYINPUT101), .A3(new_n312), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n700), .A2(new_n337), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n238), .B1(new_n702), .B2(new_n188), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n703), .B1(new_n356), .B2(new_n351), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT102), .ZN(new_n705));
  AND4_X1   g519(.A1(new_n591), .A2(new_n705), .A3(new_n635), .A4(new_n529), .ZN(new_n706));
  XOR2_X1   g520(.A(new_n687), .B(KEYINPUT39), .Z(new_n707));
  NOR2_X1   g521(.A1(new_n683), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n697), .A2(new_n706), .A3(new_n710), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(new_n243), .ZN(G45));
  INV_X1    g527(.A(new_n687), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n656), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n682), .A2(new_n684), .A3(new_n691), .A4(new_n715), .ZN(new_n716));
  XOR2_X1   g530(.A(KEYINPUT104), .B(G146), .Z(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G48));
  NAND2_X1  g532(.A1(new_n448), .A2(new_n188), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(G469), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n720), .A2(new_n535), .A3(new_n450), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n682), .A2(new_n641), .A3(new_n657), .A4(new_n721), .ZN(new_n722));
  XOR2_X1   g536(.A(KEYINPUT41), .B(G113), .Z(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(KEYINPUT105), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n722), .B(new_n724), .ZN(G15));
  NAND4_X1  g539(.A1(new_n682), .A2(new_n641), .A3(new_n663), .A4(new_n721), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G116), .ZN(G18));
  NAND2_X1  g541(.A1(new_n721), .A2(new_n691), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n591), .A2(new_n635), .A3(new_n528), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n358), .B1(new_n357), .B2(new_n334), .ZN(new_n730));
  AOI211_X1 g544(.A(KEYINPUT71), .B(new_n333), .C1(new_n356), .C2(new_n351), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g546(.A(KEYINPUT106), .B1(new_n728), .B2(new_n732), .ZN(new_n733));
  AND4_X1   g547(.A1(new_n535), .A2(new_n691), .A3(new_n450), .A4(new_n720), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT106), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n734), .A2(new_n682), .A3(new_n735), .A4(new_n729), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(KEYINPUT107), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G119), .ZN(G21));
  NAND2_X1  g553(.A1(new_n237), .A2(KEYINPUT109), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n233), .A2(new_n741), .A3(new_n234), .A4(new_n236), .ZN(new_n742));
  XOR2_X1   g556(.A(KEYINPUT108), .B(G472), .Z(new_n743));
  OAI211_X1 g557(.A(new_n343), .B(new_n344), .C1(new_n311), .C2(new_n330), .ZN(new_n744));
  AOI22_X1  g558(.A1(new_n642), .A2(new_n743), .B1(new_n335), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n740), .A2(new_n742), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(KEYINPUT110), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT110), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n740), .A2(new_n748), .A3(new_n742), .A4(new_n745), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n648), .A2(new_n591), .A3(new_n635), .A4(new_n529), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  AND4_X1   g566(.A1(new_n535), .A2(new_n720), .A3(new_n450), .A4(new_n527), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n750), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G122), .ZN(G24));
  INV_X1    g569(.A(new_n656), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n687), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n715), .A2(KEYINPUT111), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n734), .A2(new_n745), .A3(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G125), .ZN(G27));
  NAND2_X1  g577(.A1(new_n454), .A2(KEYINPUT112), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT112), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n453), .A2(new_n765), .A3(new_n446), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n764), .A2(G469), .A3(new_n455), .A4(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n450), .A2(new_n452), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(KEYINPUT113), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n450), .A2(new_n770), .A3(new_n767), .A4(new_n452), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n769), .A2(new_n535), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n530), .B1(new_n518), .B2(new_n520), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT42), .B1(new_n759), .B2(new_n760), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n772), .A2(new_n360), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n769), .A2(new_n535), .A3(new_n773), .A4(new_n771), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n759), .A2(new_n760), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n740), .A2(new_n742), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n334), .A2(new_n355), .A3(new_n340), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n776), .A2(new_n777), .A3(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT42), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n775), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(new_n272), .ZN(G33));
  NAND4_X1  g598(.A1(new_n772), .A2(new_n360), .A3(new_n690), .A4(new_n773), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G134), .ZN(G36));
  INV_X1    g600(.A(new_n773), .ZN(new_n787));
  INV_X1    g601(.A(new_n655), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n788), .A2(new_n591), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(KEYINPUT116), .ZN(new_n790));
  XOR2_X1   g604(.A(new_n790), .B(KEYINPUT43), .Z(new_n791));
  NOR3_X1   g605(.A1(new_n791), .A2(new_n645), .A3(new_n676), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n787), .B1(new_n792), .B2(KEYINPUT44), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n792), .A2(KEYINPUT44), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT45), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n456), .B1(new_n796), .B2(new_n449), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT114), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n764), .A2(KEYINPUT45), .A3(new_n455), .A4(new_n766), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n456), .B(new_n800), .C1(new_n796), .C2(new_n449), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n798), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT46), .B1(new_n802), .B2(new_n452), .ZN(new_n803));
  INV_X1    g617(.A(new_n450), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n802), .A2(KEYINPUT46), .A3(new_n452), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n535), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n707), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n795), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NOR4_X1   g625(.A1(new_n807), .A2(KEYINPUT115), .A3(new_n808), .A4(new_n707), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n793), .B(new_n794), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G137), .ZN(G39));
  OAI21_X1  g628(.A(KEYINPUT47), .B1(new_n807), .B2(new_n808), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n805), .A2(new_n806), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT47), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(new_n817), .A3(new_n535), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n682), .A2(new_n641), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n820), .A2(new_n715), .A3(new_n773), .A4(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(G140), .ZN(G42));
  NOR2_X1   g637(.A1(new_n791), .A2(new_n686), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n824), .A2(new_n721), .A3(new_n750), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(new_n648), .A3(new_n529), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n721), .A2(new_n773), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(new_n780), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT48), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n705), .A2(new_n523), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n831), .A2(new_n641), .A3(new_n827), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n656), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n830), .A2(new_n521), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT51), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n745), .A2(new_n675), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n828), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n832), .A2(new_n591), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n837), .B1(new_n838), .B2(new_n788), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n720), .A2(new_n450), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n808), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n787), .B1(new_n819), .B2(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n824), .A2(new_n750), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n840), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n825), .A2(new_n530), .A3(new_n696), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT50), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n846), .B(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n835), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n819), .A2(new_n842), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n850), .A2(new_n773), .A3(new_n844), .ZN(new_n851));
  AND4_X1   g665(.A1(new_n835), .A2(new_n851), .A3(new_n848), .A4(new_n839), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n826), .B(new_n834), .C1(new_n849), .C2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT123), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n845), .A2(new_n848), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT51), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n845), .A2(new_n835), .A3(new_n848), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n859), .A2(KEYINPUT123), .A3(new_n826), .A4(new_n834), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  XOR2_X1   g675(.A(KEYINPUT120), .B(KEYINPUT53), .Z(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n687), .B(KEYINPUT119), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n676), .A2(new_n864), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n704), .A2(new_n865), .A3(new_n751), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n866), .A2(new_n535), .A3(new_n769), .A4(new_n771), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n692), .A2(new_n716), .A3(new_n762), .A4(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT52), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n683), .B1(new_n359), .B2(new_n354), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n871), .B(new_n691), .C1(new_n690), .C2(new_n715), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n872), .A2(KEYINPUT52), .A3(new_n762), .A4(new_n867), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n775), .B(new_n785), .C1(new_n781), .C2(new_n782), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n722), .A2(new_n726), .A3(new_n754), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n878), .B1(new_n736), .B2(new_n733), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT118), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n641), .B1(new_n730), .B2(new_n731), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n637), .B1(new_n881), .B2(new_n678), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n518), .A2(new_n520), .A3(new_n531), .A4(new_n661), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT117), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n532), .A2(new_n756), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n646), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n880), .B1(new_n882), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n638), .B1(new_n360), .B2(new_n677), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n532), .A2(KEYINPUT117), .A3(new_n661), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT117), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n883), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n889), .A2(new_n885), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n647), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n888), .A2(KEYINPUT118), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n887), .A2(new_n894), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n776), .A2(new_n777), .A3(new_n836), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n636), .A2(new_n675), .A3(new_n687), .ZN(new_n897));
  AND4_X1   g711(.A1(new_n682), .A2(new_n684), .A3(new_n773), .A4(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n879), .A2(new_n895), .A3(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n863), .B1(new_n877), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT121), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n882), .A2(new_n886), .A3(new_n880), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT118), .B1(new_n888), .B2(new_n893), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n722), .A2(new_n726), .A3(new_n754), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n899), .A2(new_n906), .A3(new_n737), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n875), .B1(new_n870), .B2(new_n873), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n908), .A2(KEYINPUT53), .A3(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT54), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n899), .A2(new_n906), .A3(new_n737), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n912), .A2(new_n874), .A3(new_n895), .A4(new_n876), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT121), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n913), .A2(new_n914), .A3(new_n863), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n902), .A2(new_n910), .A3(new_n911), .A4(new_n915), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT122), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n913), .A2(new_n862), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n918), .B1(KEYINPUT53), .B2(new_n913), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(KEYINPUT54), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  OAI22_X1  g735(.A1(new_n861), .A2(new_n921), .B1(G952), .B2(G953), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT49), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n778), .B1(new_n841), .B2(new_n923), .ZN(new_n924));
  AOI211_X1 g738(.A(new_n705), .B(new_n924), .C1(new_n923), .C2(new_n841), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n789), .A2(new_n808), .A3(new_n530), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n925), .A2(new_n696), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n922), .A2(new_n927), .ZN(G75));
  AOI211_X1 g742(.A(KEYINPUT121), .B(new_n862), .C1(new_n908), .C2(new_n909), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n914), .B1(new_n913), .B2(new_n863), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n188), .B1(new_n931), .B2(new_n910), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT56), .B1(new_n932), .B2(G210), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n506), .A2(new_n509), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(new_n507), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT55), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n933), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n933), .A2(new_n937), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n221), .A2(G952), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(G51));
  XNOR2_X1  g755(.A(new_n451), .B(KEYINPUT57), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n911), .B1(new_n931), .B2(new_n910), .ZN(new_n943));
  INV_X1    g757(.A(new_n916), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n945), .A2(KEYINPUT124), .A3(new_n448), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT124), .ZN(new_n947));
  INV_X1    g761(.A(new_n942), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n902), .A2(new_n910), .A3(new_n915), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(KEYINPUT54), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n948), .B1(new_n950), .B2(new_n916), .ZN(new_n951));
  INV_X1    g765(.A(new_n448), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n947), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n802), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n932), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n946), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n940), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n956), .A2(new_n957), .ZN(G54));
  INV_X1    g772(.A(KEYINPUT58), .ZN(new_n959));
  OAI21_X1  g773(.A(KEYINPUT125), .B1(new_n959), .B2(new_n583), .ZN(new_n960));
  OR3_X1    g774(.A1(new_n959), .A2(new_n583), .A3(KEYINPUT125), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n932), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(new_n582), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n963), .A2(new_n957), .ZN(G60));
  NAND2_X1  g778(.A1(G478), .A2(G902), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT59), .Z(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n650), .B1(new_n921), .B2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n650), .ZN(new_n969));
  AOI211_X1 g783(.A(new_n969), .B(new_n966), .C1(new_n950), .C2(new_n916), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n968), .A2(new_n940), .A3(new_n970), .ZN(G63));
  NAND2_X1  g785(.A1(G217), .A2(G902), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT60), .Z(new_n973));
  OAI211_X1 g787(.A(new_n949), .B(new_n973), .C1(new_n673), .C2(new_n672), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n949), .A2(new_n973), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n974), .B(new_n957), .C1(new_n975), .C2(new_n227), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT61), .Z(G66));
  AOI21_X1  g791(.A(new_n221), .B1(new_n524), .B2(G224), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n879), .A2(new_n895), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n978), .B1(new_n979), .B2(new_n221), .ZN(new_n980));
  INV_X1    g794(.A(G898), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n934), .B1(new_n981), .B2(G953), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n980), .B(new_n982), .ZN(G69));
  AND2_X1   g797(.A1(new_n872), .A2(new_n762), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n712), .A2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT62), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n712), .A2(KEYINPUT62), .A3(new_n984), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n662), .A2(new_n656), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n360), .A2(new_n708), .A3(new_n773), .A4(new_n990), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n989), .A2(new_n822), .A3(new_n813), .A4(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n221), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n299), .B(new_n574), .Z(new_n994));
  AOI21_X1  g808(.A(KEYINPUT126), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT126), .ZN(new_n996));
  INV_X1    g810(.A(new_n994), .ZN(new_n997));
  AOI211_X1 g811(.A(new_n996), .B(new_n997), .C1(new_n992), .C2(new_n221), .ZN(new_n998));
  OR2_X1    g812(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(G900), .ZN(new_n1000));
  OAI21_X1  g814(.A(G953), .B1(new_n430), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT127), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OR2_X1    g817(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n822), .A2(new_n813), .ZN(new_n1005));
  INV_X1    g819(.A(new_n780), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n752), .B(new_n1006), .C1(new_n811), .C2(new_n812), .ZN(new_n1007));
  AND2_X1   g821(.A1(new_n1007), .A2(new_n876), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n1005), .A2(new_n1008), .A3(new_n221), .A4(new_n984), .ZN(new_n1009));
  OAI211_X1 g823(.A(new_n1009), .B(new_n997), .C1(new_n1000), .C2(new_n221), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n999), .A2(new_n1003), .A3(new_n1004), .A4(new_n1010), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1010), .B1(new_n995), .B2(new_n998), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1012), .A2(new_n1002), .A3(new_n1001), .ZN(new_n1013));
  AND2_X1   g827(.A1(new_n1011), .A2(new_n1013), .ZN(G72));
  NAND2_X1  g828(.A1(G472), .A2(G902), .ZN(new_n1015));
  XOR2_X1   g829(.A(new_n1015), .B(KEYINPUT63), .Z(new_n1016));
  NAND3_X1  g830(.A1(new_n1005), .A2(new_n1008), .A3(new_n984), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1016), .B1(new_n1017), .B2(new_n979), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n1018), .A2(new_n303), .A3(new_n304), .A4(new_n312), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1016), .B1(new_n992), .B2(new_n979), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n1020), .A2(new_n305), .A3(new_n311), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n313), .A2(new_n337), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n919), .A2(new_n1016), .A3(new_n1022), .ZN(new_n1023));
  AND4_X1   g837(.A1(new_n957), .A2(new_n1019), .A3(new_n1021), .A4(new_n1023), .ZN(G57));
endmodule


