//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 0 0 0 1 0 0 1 0 0 0 1 0 0 0 0 1 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 1 0 1 0 1 1 1 0 0 0 1 1 0 0 1 0 0 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n865, new_n866, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT11), .B(G169gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT12), .ZN(new_n206));
  INV_X1    g005(.A(G8gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(G15gat), .B(G22gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT90), .ZN(new_n209));
  AND2_X1   g008(.A1(new_n209), .A2(G1gat), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT16), .B1(new_n209), .B2(G1gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n208), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT91), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n207), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n212), .B1(G1gat), .B2(new_n208), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI221_X1 g015(.A(new_n212), .B1(new_n213), .B2(new_n207), .C1(G1gat), .C2(new_n208), .ZN(new_n217));
  INV_X1    g016(.A(G29gat), .ZN(new_n218));
  INV_X1    g017(.A(G36gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT14), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT14), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(G29gat), .B2(G36gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(G29gat), .A2(G36gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n220), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT15), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n220), .A2(new_n222), .A3(KEYINPUT15), .A4(new_n223), .ZN(new_n227));
  XNOR2_X1  g026(.A(G43gat), .B(G50gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n220), .A2(new_n223), .ZN(new_n230));
  XOR2_X1   g029(.A(G43gat), .B(G50gat), .Z(new_n231));
  NAND4_X1  g030(.A1(new_n230), .A2(KEYINPUT15), .A3(new_n222), .A4(new_n231), .ZN(new_n232));
  AOI22_X1  g031(.A1(new_n216), .A2(new_n217), .B1(new_n229), .B2(new_n232), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n224), .A2(new_n225), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n227), .A2(new_n228), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n232), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT17), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT17), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n232), .B(new_n238), .C1(new_n234), .C2(new_n235), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n216), .A2(new_n217), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n233), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G229gat), .A2(G233gat), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n244), .A2(KEYINPUT18), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n241), .A2(new_n236), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n216), .A2(new_n217), .A3(new_n229), .A4(new_n232), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(new_n244), .B(KEYINPUT13), .Z(new_n249));
  AOI22_X1  g048(.A1(new_n243), .A2(new_n245), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n239), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n238), .B1(new_n229), .B2(new_n232), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n244), .B(new_n246), .C1(new_n253), .C2(new_n241), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n206), .B1(new_n250), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n250), .A2(new_n256), .A3(new_n206), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT93), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n250), .A2(new_n256), .A3(KEYINPUT93), .A4(new_n206), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n257), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(G183gat), .A2(G190gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT24), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT24), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n265), .A2(G183gat), .A3(G190gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n268));
  OR3_X1    g067(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  AND3_X1   g069(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT65), .ZN(new_n273));
  OR3_X1    g072(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT25), .ZN(new_n275));
  NOR2_X1   g074(.A1(G169gat), .A2(G176gat), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT23), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n275), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n273), .B1(new_n271), .B2(new_n272), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n270), .A2(new_n274), .A3(new_n280), .A4(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n279), .ZN(new_n283));
  NOR3_X1   g082(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n284));
  OAI22_X1  g083(.A1(new_n283), .A2(new_n284), .B1(new_n271), .B2(new_n272), .ZN(new_n285));
  INV_X1    g084(.A(G183gat), .ZN(new_n286));
  INV_X1    g085(.A(G190gat), .ZN(new_n287));
  AOI22_X1  g086(.A1(new_n264), .A2(new_n266), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n275), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n282), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT26), .ZN(new_n291));
  OAI22_X1  g090(.A1(new_n271), .A2(new_n272), .B1(new_n291), .B2(new_n276), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT67), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI221_X1 g093(.A(KEYINPUT67), .B1(new_n276), .B2(new_n291), .C1(new_n271), .C2(new_n272), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n276), .A2(new_n291), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n263), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n286), .A2(KEYINPUT27), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT27), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(G183gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n301), .A3(new_n287), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT28), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(KEYINPUT27), .B(G183gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n305), .A2(KEYINPUT28), .A3(new_n287), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n298), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n297), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G113gat), .ZN(new_n309));
  INV_X1    g108(.A(G120gat), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT1), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n311), .B1(new_n309), .B2(new_n310), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT69), .ZN(new_n313));
  INV_X1    g112(.A(G134gat), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n313), .B1(new_n314), .B2(G127gat), .ZN(new_n315));
  INV_X1    g114(.A(G127gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n316), .A2(KEYINPUT69), .A3(G134gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n314), .A2(KEYINPUT68), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT68), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G134gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n315), .B(new_n317), .C1(new_n321), .C2(new_n316), .ZN(new_n322));
  XNOR2_X1  g121(.A(KEYINPUT70), .B(G120gat), .ZN(new_n323));
  OR2_X1    g122(.A1(new_n323), .A2(new_n309), .ZN(new_n324));
  XNOR2_X1  g123(.A(G127gat), .B(G134gat), .ZN(new_n325));
  AND2_X1   g124(.A1(new_n325), .A2(new_n311), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n312), .A2(new_n322), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n290), .A2(new_n308), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT71), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT71), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n290), .A2(new_n308), .A3(new_n330), .A4(new_n327), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n290), .A2(new_n308), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n322), .A2(new_n312), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n324), .A2(new_n326), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n329), .A2(new_n331), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(G227gat), .A2(G233gat), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G15gat), .B(G43gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(G71gat), .B(G99gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT33), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n340), .A2(KEYINPUT32), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT73), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n340), .A2(KEYINPUT73), .A3(KEYINPUT32), .A4(new_n345), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n327), .B1(new_n290), .B2(new_n308), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n351), .B1(KEYINPUT71), .B2(new_n328), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n338), .B1(new_n352), .B2(new_n331), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n344), .B1(new_n353), .B2(KEYINPUT33), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT32), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT72), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT33), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n343), .B1(new_n340), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT72), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n359), .B(new_n360), .C1(new_n355), .C2(new_n353), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n350), .A2(new_n357), .A3(new_n361), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n329), .A2(new_n336), .A3(new_n338), .A4(new_n331), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT74), .ZN(new_n364));
  OR3_X1    g163(.A1(new_n363), .A2(new_n364), .A3(KEYINPUT34), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(KEYINPUT34), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n364), .B1(new_n363), .B2(KEYINPUT34), .ZN(new_n367));
  AND3_X1   g166(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n362), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT76), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n368), .A2(new_n350), .A3(new_n357), .A4(new_n361), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT36), .ZN(new_n374));
  AND2_X1   g173(.A1(new_n357), .A2(new_n361), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n375), .A2(KEYINPUT76), .A3(new_n368), .A4(new_n350), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n373), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n370), .A2(KEYINPUT75), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n372), .A2(KEYINPUT36), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT75), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n362), .A2(new_n380), .A3(new_n369), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n378), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G8gat), .B(G36gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(G64gat), .B(G92gat), .ZN(new_n385));
  XOR2_X1   g184(.A(new_n384), .B(new_n385), .Z(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n332), .A2(KEYINPUT77), .ZN(new_n388));
  INV_X1    g187(.A(G226gat), .ZN(new_n389));
  INV_X1    g188(.A(G233gat), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT77), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n290), .A2(new_n308), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n388), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(G197gat), .B(G204gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(G211gat), .A2(G218gat), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT22), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  OR2_X1    g198(.A1(G211gat), .A2(G218gat), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(new_n396), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n396), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n402), .A2(new_n395), .A3(new_n398), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n391), .A2(KEYINPUT29), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n332), .A2(new_n406), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n394), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n290), .A2(new_n308), .A3(new_n392), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n392), .B1(new_n290), .B2(new_n308), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n406), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n290), .A2(new_n308), .A3(new_n391), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n405), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n387), .B1(new_n408), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT37), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n414), .B1(new_n415), .B2(new_n386), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n394), .A2(new_n407), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n415), .B1(new_n417), .B2(new_n404), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n404), .B1(new_n411), .B2(new_n412), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT38), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT89), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n416), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n406), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n424), .B1(new_n388), .B2(new_n393), .ZN(new_n425));
  INV_X1    g224(.A(new_n412), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n404), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n394), .A2(new_n405), .A3(new_n407), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n386), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n386), .A2(new_n415), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT38), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n394), .A2(new_n407), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT37), .B1(new_n433), .B2(new_n405), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n432), .B1(new_n434), .B2(new_n419), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT89), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n423), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G1gat), .B(G29gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(KEYINPUT0), .ZN(new_n439));
  XNOR2_X1  g238(.A(G57gat), .B(G85gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n439), .B(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G225gat), .A2(G233gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(KEYINPUT80), .B(KEYINPUT2), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(G141gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(G148gat), .ZN(new_n446));
  INV_X1    g245(.A(G148gat), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(G141gat), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT79), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n446), .A2(new_n448), .A3(KEYINPUT79), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n444), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OR2_X1    g251(.A1(G155gat), .A2(G162gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(G155gat), .A2(G162gat), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT81), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n456), .B1(new_n447), .B2(G141gat), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n445), .A2(KEYINPUT81), .A3(G148gat), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(new_n458), .A3(new_n448), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n454), .B1(new_n453), .B2(KEYINPUT2), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n459), .A2(new_n460), .A3(KEYINPUT82), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT82), .B1(new_n459), .B2(new_n460), .ZN(new_n462));
  OAI22_X1  g261(.A1(new_n452), .A2(new_n455), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n335), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n459), .A2(new_n460), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT82), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n459), .A2(new_n460), .A3(KEYINPUT82), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n446), .A2(new_n448), .A3(KEYINPUT79), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n443), .B1(new_n469), .B2(new_n449), .ZN(new_n470));
  INV_X1    g269(.A(new_n455), .ZN(new_n471));
  AOI22_X1  g270(.A1(new_n467), .A2(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n327), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n442), .B1(new_n464), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT5), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT85), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n442), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n463), .A2(new_n335), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n472), .A2(new_n327), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT85), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(new_n481), .A3(KEYINPUT5), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT4), .B1(new_n463), .B2(new_n335), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT83), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT4), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n472), .A2(new_n485), .A3(new_n327), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT84), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT83), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n473), .A2(new_n488), .A3(KEYINPUT4), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT84), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n472), .A2(new_n490), .A3(new_n485), .A4(new_n327), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n484), .A2(new_n487), .A3(new_n489), .A4(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT3), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n472), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(new_n495), .A3(new_n335), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n496), .A2(new_n442), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n476), .A2(new_n482), .B1(new_n492), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n486), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n497), .A2(new_n475), .A3(new_n499), .ZN(new_n500));
  OAI211_X1 g299(.A(KEYINPUT6), .B(new_n441), .C1(new_n498), .C2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n441), .B1(new_n498), .B2(new_n500), .ZN(new_n502));
  INV_X1    g301(.A(new_n441), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n497), .A2(new_n475), .A3(new_n499), .ZN(new_n504));
  AND2_X1   g303(.A1(new_n482), .A2(new_n476), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n496), .A2(new_n442), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n483), .A2(KEYINPUT83), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n488), .B1(new_n473), .B2(KEYINPUT4), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n487), .A2(new_n491), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n503), .B(new_n504), .C1(new_n505), .C2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT6), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n502), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n408), .A2(new_n413), .A3(new_n387), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT37), .B1(new_n408), .B2(new_n413), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(new_n429), .B2(new_n430), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n515), .B1(new_n517), .B2(KEYINPUT38), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n437), .A2(new_n501), .A3(new_n514), .A4(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(G228gat), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n520), .A2(new_n390), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT29), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(new_n405), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT29), .B1(new_n401), .B2(new_n403), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n494), .B1(new_n525), .B2(KEYINPUT86), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT86), .ZN(new_n527));
  AOI211_X1 g326(.A(new_n527), .B(KEYINPUT29), .C1(new_n401), .C2(new_n403), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n463), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n521), .B1(new_n524), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n404), .B1(new_n495), .B2(new_n522), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n463), .A2(new_n525), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n532), .A2(new_n493), .A3(new_n521), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(G22gat), .B1(new_n530), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT87), .ZN(new_n536));
  XOR2_X1   g335(.A(G78gat), .B(G106gat), .Z(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT31), .B(G50gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n521), .ZN(new_n540));
  INV_X1    g339(.A(new_n529), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n540), .B1(new_n541), .B2(new_n531), .ZN(new_n542));
  OR2_X1    g341(.A1(new_n531), .A2(new_n533), .ZN(new_n543));
  INV_X1    g342(.A(G22gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  AOI22_X1  g344(.A1(new_n536), .A2(new_n539), .B1(new_n535), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT87), .ZN(new_n547));
  AND4_X1   g346(.A1(new_n547), .A2(new_n545), .A3(new_n535), .A4(new_n539), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n442), .B1(new_n499), .B2(new_n496), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n464), .A2(new_n473), .A3(new_n442), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT39), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT39), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n441), .B1(new_n550), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT40), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n553), .A2(KEYINPUT40), .A3(new_n555), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n558), .A2(new_n502), .A3(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT30), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n562), .A2(KEYINPUT78), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n563), .B1(new_n515), .B2(new_n429), .ZN(new_n564));
  INV_X1    g363(.A(new_n563), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n427), .A2(new_n428), .A3(new_n386), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n562), .A2(KEYINPUT78), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n565), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT88), .B1(new_n561), .B2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n569), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n565), .B1(new_n414), .B2(new_n566), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT88), .ZN(new_n575));
  NOR3_X1   g374(.A1(new_n574), .A2(new_n560), .A3(new_n575), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n519), .B(new_n549), .C1(new_n571), .C2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n570), .B1(new_n501), .B2(new_n514), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n383), .B(new_n577), .C1(new_n578), .C2(new_n549), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n549), .A2(new_n372), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n580), .A2(new_n378), .A3(new_n578), .A4(new_n381), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT35), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n373), .A2(new_n376), .ZN(new_n583));
  INV_X1    g382(.A(new_n549), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n584), .A2(KEYINPUT35), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n583), .A2(new_n578), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n262), .B1(new_n579), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT21), .ZN(new_n589));
  XNOR2_X1  g388(.A(G57gat), .B(G64gat), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(G71gat), .ZN(new_n592));
  INV_X1    g391(.A(G78gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G71gat), .A2(G78gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT9), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n591), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  OAI211_X1 g398(.A(new_n595), .B(new_n594), .C1(new_n590), .C2(new_n597), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n242), .B1(new_n589), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n589), .ZN(new_n603));
  XOR2_X1   g402(.A(KEYINPUT95), .B(KEYINPUT19), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n602), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G127gat), .B(G155gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT20), .ZN(new_n608));
  NAND2_X1  g407(.A1(G231gat), .A2(G233gat), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n609), .B(KEYINPUT94), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n608), .B(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G183gat), .B(G211gat), .Z(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT96), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n611), .B(new_n613), .ZN(new_n614));
  OR2_X1    g413(.A1(new_n606), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n606), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g416(.A1(G232gat), .A2(G233gat), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n618), .A2(KEYINPUT41), .ZN(new_n619));
  XNOR2_X1  g418(.A(G134gat), .B(G162gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G85gat), .A2(G92gat), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT7), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT97), .ZN(new_n628));
  XNOR2_X1  g427(.A(G99gat), .B(G106gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(G99gat), .A2(G106gat), .ZN(new_n630));
  INV_X1    g429(.A(G85gat), .ZN(new_n631));
  INV_X1    g430(.A(G92gat), .ZN(new_n632));
  AOI22_X1  g431(.A1(KEYINPUT8), .A2(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n627), .A2(new_n628), .A3(new_n629), .A4(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n630), .A2(KEYINPUT8), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n631), .A2(new_n632), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n635), .A2(new_n625), .A3(new_n636), .A4(new_n626), .ZN(new_n637));
  INV_X1    g436(.A(new_n629), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n633), .A2(new_n629), .A3(new_n625), .A4(new_n626), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n639), .A2(KEYINPUT97), .A3(new_n640), .ZN(new_n641));
  OAI211_X1 g440(.A(new_n634), .B(new_n641), .C1(new_n251), .C2(new_n252), .ZN(new_n642));
  XOR2_X1   g441(.A(G190gat), .B(G218gat), .Z(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n641), .A2(new_n634), .ZN(new_n645));
  AOI22_X1  g444(.A1(new_n645), .A2(new_n236), .B1(KEYINPUT41), .B2(new_n618), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n642), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n644), .B1(new_n642), .B2(new_n646), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n622), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n649), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n651), .A2(new_n621), .A3(new_n647), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n617), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT98), .ZN(new_n655));
  XNOR2_X1  g454(.A(G120gat), .B(G148gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(G176gat), .B(G204gat), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n656), .B(new_n657), .Z(new_n658));
  INV_X1    g457(.A(G230gat), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n659), .A2(new_n390), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n641), .A2(new_n601), .A3(new_n634), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT10), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n599), .A2(new_n639), .A3(new_n600), .A4(new_n640), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n601), .A2(new_n662), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n645), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n660), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n660), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n669), .B1(new_n661), .B2(new_n663), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n658), .B1(new_n668), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n658), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n667), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n655), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n588), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n514), .A2(new_n501), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT99), .B(G1gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1324gat));
  INV_X1    g482(.A(new_n678), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT16), .B(G8gat), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n684), .A2(new_n574), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n207), .B1(new_n678), .B2(new_n570), .ZN(new_n687));
  OAI21_X1  g486(.A(KEYINPUT42), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n688), .B1(KEYINPUT42), .B2(new_n686), .ZN(G1325gat));
  OAI21_X1  g488(.A(G15gat), .B1(new_n684), .B2(new_n383), .ZN(new_n690));
  INV_X1    g489(.A(new_n583), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n691), .A2(G15gat), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n690), .B1(new_n684), .B2(new_n692), .ZN(G1326gat));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n584), .ZN(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT43), .B(G22gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1327gat));
  INV_X1    g495(.A(new_n617), .ZN(new_n697));
  INV_X1    g496(.A(new_n653), .ZN(new_n698));
  AND4_X1   g497(.A1(new_n588), .A2(new_n697), .A3(new_n698), .A4(new_n675), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n699), .A2(new_n218), .A3(new_n680), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT45), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT100), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n702), .B1(new_n578), .B2(new_n549), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n679), .A2(new_n574), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n704), .A2(KEYINPUT100), .A3(new_n584), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n383), .A2(new_n706), .A3(new_n577), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n587), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n698), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n579), .A2(new_n587), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n712), .A2(KEYINPUT44), .A3(new_n698), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n262), .A2(new_n617), .A3(new_n676), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(G29gat), .B1(new_n716), .B2(new_n679), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n717), .ZN(G1328gat));
  OAI21_X1  g517(.A(G36gat), .B1(new_n716), .B2(new_n574), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n699), .A2(new_n219), .A3(new_n570), .ZN(new_n720));
  AND2_X1   g519(.A1(KEYINPUT101), .A2(KEYINPUT46), .ZN(new_n721));
  NOR2_X1   g520(.A1(KEYINPUT101), .A2(KEYINPUT46), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n719), .B(new_n723), .C1(new_n721), .C2(new_n720), .ZN(G1329gat));
  INV_X1    g523(.A(G43gat), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n383), .A2(new_n725), .ZN(new_n726));
  AND3_X1   g525(.A1(new_n714), .A2(new_n715), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(G43gat), .B1(new_n699), .B2(new_n583), .ZN(new_n728));
  OAI21_X1  g527(.A(KEYINPUT47), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n728), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT47), .ZN(new_n731));
  INV_X1    g530(.A(new_n726), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n730), .B(new_n731), .C1(new_n716), .C2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n729), .A2(new_n733), .ZN(G1330gat));
  NAND4_X1  g533(.A1(new_n711), .A2(new_n584), .A3(new_n713), .A4(new_n715), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(G50gat), .ZN(new_n736));
  INV_X1    g535(.A(G50gat), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n699), .A2(new_n737), .A3(new_n584), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT48), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n736), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n739), .B1(new_n736), .B2(new_n738), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n740), .A2(new_n741), .ZN(G1331gat));
  NAND2_X1  g541(.A1(new_n260), .A2(new_n261), .ZN(new_n743));
  INV_X1    g542(.A(new_n257), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n655), .A2(new_n745), .A3(new_n675), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n708), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n680), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g549(.A1(new_n747), .A2(new_n574), .ZN(new_n751));
  NOR2_X1   g550(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n752));
  AND2_X1   g551(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n751), .B2(new_n752), .ZN(G1333gat));
  INV_X1    g554(.A(new_n383), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n748), .A2(G71gat), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n583), .B(KEYINPUT102), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n592), .B1(new_n747), .B2(new_n758), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n760), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g560(.A1(new_n747), .A2(new_n549), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(new_n593), .ZN(G1335gat));
  NOR2_X1   g562(.A1(new_n745), .A2(new_n617), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n708), .A2(new_n698), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT51), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n708), .A2(new_n767), .A3(new_n698), .A4(new_n764), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n766), .A2(new_n676), .A3(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n769), .A2(new_n631), .A3(new_n680), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n745), .A2(new_n617), .A3(new_n675), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n714), .A2(new_n680), .A3(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n770), .B1(new_n772), .B2(new_n631), .ZN(G1336gat));
  NOR2_X1   g572(.A1(new_n574), .A2(G92gat), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n766), .A2(new_n676), .A3(new_n768), .A4(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT103), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n675), .B1(new_n765), .B2(KEYINPUT51), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n778), .A2(KEYINPUT103), .A3(new_n768), .A4(new_n774), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n711), .A2(new_n570), .A3(new_n713), .A4(new_n771), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(G92gat), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n777), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT52), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT104), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n769), .A2(new_n784), .A3(new_n774), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n775), .A2(KEYINPUT104), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n785), .A2(new_n786), .A3(new_n781), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n783), .A2(new_n788), .ZN(G1337gat));
  INV_X1    g588(.A(G99gat), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n711), .A2(new_n756), .A3(new_n713), .A4(new_n771), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT105), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n793), .B1(new_n792), .B2(new_n791), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n769), .A2(new_n790), .A3(new_n583), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(G1338gat));
  AND4_X1   g595(.A1(new_n584), .A2(new_n711), .A3(new_n713), .A4(new_n771), .ZN(new_n797));
  INV_X1    g596(.A(G106gat), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n778), .A2(new_n768), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n584), .A2(new_n798), .ZN(new_n800));
  OAI22_X1  g599(.A1(new_n797), .A2(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  XOR2_X1   g600(.A(KEYINPUT106), .B(KEYINPUT53), .Z(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n802), .ZN(new_n804));
  OAI221_X1 g603(.A(new_n804), .B1(new_n799), .B2(new_n800), .C1(new_n797), .C2(new_n798), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(G1339gat));
  NOR3_X1   g605(.A1(new_n655), .A2(new_n745), .A3(new_n676), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT107), .ZN(new_n809));
  AOI211_X1 g608(.A(KEYINPUT54), .B(new_n660), .C1(new_n664), .C2(new_n666), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n809), .B1(new_n810), .B2(new_n658), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n664), .A2(new_n666), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n812), .A2(new_n813), .A3(new_n669), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n814), .A2(KEYINPUT107), .A3(new_n673), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n664), .A2(new_n660), .A3(new_n666), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n668), .A2(KEYINPUT54), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n653), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AOI211_X1 g620(.A(new_n809), .B(new_n658), .C1(new_n667), .C2(new_n813), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT107), .B1(new_n814), .B2(new_n673), .ZN(new_n823));
  OAI211_X1 g622(.A(KEYINPUT55), .B(new_n818), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n674), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n205), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n243), .A2(new_n244), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n248), .A2(new_n249), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n830), .B1(new_n260), .B2(new_n261), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n821), .A2(new_n826), .A3(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT108), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n821), .A2(new_n826), .A3(KEYINPUT108), .A4(new_n831), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT55), .B1(new_n816), .B2(new_n818), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n745), .A2(new_n826), .A3(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT109), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n831), .A2(new_n840), .A3(new_n676), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n831), .B2(new_n676), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n839), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n698), .B1(new_n843), .B2(KEYINPUT110), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT110), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n845), .B(new_n839), .C1(new_n841), .C2(new_n842), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n836), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n808), .B1(new_n847), .B2(new_n617), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n848), .A2(new_n549), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n679), .A2(new_n570), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n691), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n853), .A2(new_n309), .A3(new_n262), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n848), .A2(new_n680), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n580), .A2(new_n378), .A3(new_n381), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n856), .A2(new_n574), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n745), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n854), .B1(new_n309), .B2(new_n860), .ZN(G1340gat));
  OAI21_X1  g660(.A(G120gat), .B1(new_n853), .B2(new_n675), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n676), .A2(new_n323), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n862), .B1(new_n858), .B2(new_n863), .ZN(G1341gat));
  AOI21_X1  g663(.A(G127gat), .B1(new_n859), .B2(new_n617), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n849), .A2(G127gat), .A3(new_n617), .A4(new_n852), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n866), .A2(KEYINPUT111), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n866), .A2(KEYINPUT111), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n865), .A2(new_n867), .A3(new_n868), .ZN(G1342gat));
  OAI21_X1  g668(.A(G134gat), .B1(new_n853), .B2(new_n653), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n653), .A2(new_n321), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(KEYINPUT56), .B1(new_n858), .B2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT56), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n855), .A2(new_n874), .A3(new_n857), .A4(new_n871), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n870), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT112), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n870), .A2(new_n873), .A3(KEYINPUT112), .A4(new_n875), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(G1343gat));
  NOR2_X1   g679(.A1(new_n756), .A2(new_n851), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT57), .B1(new_n848), .B2(new_n584), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n584), .A2(KEYINPUT57), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT113), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n824), .A2(new_n825), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n262), .A2(new_n885), .A3(new_n837), .ZN(new_n886));
  AOI211_X1 g685(.A(new_n830), .B(new_n675), .C1(new_n260), .C2(new_n261), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n884), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n831), .A2(new_n676), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n839), .A2(KEYINPUT113), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n888), .A2(new_n653), .A3(new_n890), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n834), .A2(new_n835), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n617), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n807), .B1(new_n893), .B2(KEYINPUT114), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT114), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n262), .A2(new_n837), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n887), .B1(new_n896), .B2(new_n826), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n698), .B1(new_n897), .B2(KEYINPUT113), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n836), .B1(new_n898), .B2(new_n888), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n895), .B1(new_n899), .B2(new_n617), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n883), .B1(new_n894), .B2(new_n900), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n745), .B(new_n881), .C1(new_n882), .C2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(G141gat), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT115), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n756), .A2(new_n570), .A3(new_n549), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n855), .A2(new_n445), .A3(new_n745), .A4(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n904), .A2(new_n907), .A3(KEYINPUT58), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT58), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n903), .B(new_n906), .C1(KEYINPUT115), .C2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(G1344gat));
  NAND2_X1  g710(.A1(new_n855), .A2(new_n905), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(new_n447), .A3(new_n676), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT59), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(G148gat), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n882), .A2(new_n901), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n917), .A2(new_n756), .A3(new_n851), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n916), .B1(new_n918), .B2(new_n676), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n848), .A2(new_n584), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT57), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n549), .A2(KEYINPUT57), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n617), .B1(new_n891), .B2(new_n832), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n923), .B2(new_n807), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n921), .A2(new_n676), .A3(new_n881), .A4(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n915), .B1(new_n925), .B2(G148gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n914), .B1(new_n919), .B2(new_n926), .ZN(G1345gat));
  INV_X1    g726(.A(G155gat), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n913), .A2(new_n928), .A3(new_n617), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n918), .A2(new_n617), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n929), .B1(new_n930), .B2(new_n928), .ZN(G1346gat));
  AOI21_X1  g730(.A(G162gat), .B1(new_n913), .B2(new_n698), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n698), .A2(G162gat), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n932), .B1(new_n918), .B2(new_n933), .ZN(G1347gat));
  NAND2_X1  g733(.A1(new_n679), .A2(new_n570), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n758), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n849), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(G169gat), .B1(new_n937), .B2(new_n262), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n848), .A2(new_n679), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n856), .A2(new_n570), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n262), .A2(G169gat), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n938), .A2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT116), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n943), .B(new_n944), .ZN(G1348gat));
  NAND2_X1  g744(.A1(new_n676), .A2(G176gat), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n937), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n939), .A2(new_n940), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n948), .A2(new_n675), .ZN(new_n949));
  OAI22_X1  g748(.A1(KEYINPUT117), .A2(new_n947), .B1(new_n949), .B2(G176gat), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n950), .B1(KEYINPUT117), .B2(new_n947), .ZN(G1349gat));
  NAND4_X1  g750(.A1(new_n848), .A2(new_n936), .A3(new_n549), .A4(new_n617), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n286), .B1(new_n952), .B2(KEYINPUT118), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n953), .B1(KEYINPUT118), .B2(new_n952), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n939), .A2(new_n305), .A3(new_n617), .A4(new_n940), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT60), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n957), .A2(KEYINPUT119), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n954), .B(new_n955), .C1(KEYINPUT119), .C2(new_n957), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(G1350gat));
  NOR3_X1   g760(.A1(new_n948), .A2(G190gat), .A3(new_n653), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT61), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n849), .A2(new_n698), .A3(new_n936), .ZN(new_n964));
  AOI21_X1  g763(.A(KEYINPUT120), .B1(new_n964), .B2(G190gat), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n962), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  OR2_X1    g765(.A1(new_n965), .A2(new_n963), .ZN(new_n967));
  AND3_X1   g766(.A1(new_n964), .A2(KEYINPUT120), .A3(G190gat), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(G1351gat));
  NOR3_X1   g768(.A1(new_n756), .A2(new_n574), .A3(new_n549), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n939), .A2(new_n970), .ZN(new_n971));
  INV_X1    g770(.A(new_n971), .ZN(new_n972));
  XNOR2_X1  g771(.A(KEYINPUT121), .B(G197gat), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n972), .A2(new_n745), .A3(new_n973), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n756), .A2(new_n935), .ZN(new_n975));
  NAND4_X1  g774(.A1(new_n921), .A2(new_n745), .A3(new_n924), .A4(new_n975), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT122), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g777(.A(new_n973), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n979), .B1(new_n976), .B2(new_n977), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n974), .B1(new_n978), .B2(new_n980), .ZN(G1352gat));
  NAND2_X1  g780(.A1(new_n921), .A2(new_n924), .ZN(new_n982));
  INV_X1    g781(.A(new_n975), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g783(.A(new_n984), .ZN(new_n985));
  OAI21_X1  g784(.A(G204gat), .B1(new_n985), .B2(new_n675), .ZN(new_n986));
  NOR2_X1   g785(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n987));
  NAND2_X1  g786(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n988));
  OR2_X1    g787(.A1(new_n675), .A2(G204gat), .ZN(new_n989));
  OR3_X1    g788(.A1(new_n971), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n988), .B1(new_n971), .B2(new_n989), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n987), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n986), .A2(new_n992), .ZN(G1353gat));
  NAND4_X1  g792(.A1(new_n921), .A2(new_n617), .A3(new_n924), .A4(new_n975), .ZN(new_n994));
  INV_X1    g793(.A(G211gat), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT63), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n995), .B1(KEYINPUT125), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g797(.A1(new_n996), .A2(KEYINPUT125), .ZN(new_n999));
  OR2_X1    g798(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n998), .A2(new_n999), .ZN(new_n1001));
  NAND4_X1  g800(.A1(new_n939), .A2(new_n995), .A3(new_n617), .A4(new_n970), .ZN(new_n1002));
  XNOR2_X1  g801(.A(new_n1002), .B(KEYINPUT124), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n1000), .A2(new_n1001), .A3(new_n1003), .ZN(G1354gat));
  AOI21_X1  g803(.A(G218gat), .B1(new_n972), .B2(new_n698), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n985), .A2(KEYINPUT126), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n698), .A2(G218gat), .ZN(new_n1007));
  XNOR2_X1  g806(.A(new_n1007), .B(KEYINPUT127), .ZN(new_n1008));
  INV_X1    g807(.A(KEYINPUT126), .ZN(new_n1009));
  AOI21_X1  g808(.A(new_n1008), .B1(new_n984), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g809(.A(new_n1005), .B1(new_n1006), .B2(new_n1010), .ZN(G1355gat));
endmodule


