

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581;

  XNOR2_X1 U322 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U323 ( .A(n331), .B(n330), .ZN(n332) );
  INV_X1 U324 ( .A(KEYINPUT66), .ZN(n345) );
  XNOR2_X1 U325 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U326 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U327 ( .A(KEYINPUT113), .B(KEYINPUT47), .ZN(n373) );
  XOR2_X1 U328 ( .A(G99GAT), .B(G85GAT), .Z(n325) );
  XNOR2_X1 U329 ( .A(n325), .B(n311), .ZN(n313) );
  XNOR2_X1 U330 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U331 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U332 ( .A(n333), .B(n332), .ZN(n337) );
  XNOR2_X1 U333 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U334 ( .A(n343), .B(n342), .Z(n564) );
  XNOR2_X1 U335 ( .A(n461), .B(G204GAT), .ZN(n462) );
  XNOR2_X1 U336 ( .A(n450), .B(KEYINPUT50), .ZN(n451) );
  XNOR2_X1 U337 ( .A(n463), .B(n462), .ZN(G1353GAT) );
  XOR2_X1 U338 ( .A(KEYINPUT85), .B(KEYINPUT83), .Z(n291) );
  XNOR2_X1 U339 ( .A(G64GAT), .B(KEYINPUT84), .ZN(n290) );
  XNOR2_X1 U340 ( .A(n291), .B(n290), .ZN(n295) );
  XOR2_X1 U341 ( .A(G155GAT), .B(G211GAT), .Z(n293) );
  XNOR2_X1 U342 ( .A(G22GAT), .B(G8GAT), .ZN(n292) );
  XNOR2_X1 U343 ( .A(n293), .B(n292), .ZN(n294) );
  XNOR2_X1 U344 ( .A(n295), .B(n294), .ZN(n310) );
  XOR2_X1 U345 ( .A(G78GAT), .B(G71GAT), .Z(n297) );
  XNOR2_X1 U346 ( .A(G183GAT), .B(G127GAT), .ZN(n296) );
  XNOR2_X1 U347 ( .A(n297), .B(n296), .ZN(n302) );
  XNOR2_X1 U348 ( .A(G57GAT), .B(KEYINPUT77), .ZN(n298) );
  XNOR2_X1 U349 ( .A(n298), .B(KEYINPUT13), .ZN(n312) );
  XOR2_X1 U350 ( .A(n312), .B(KEYINPUT15), .Z(n300) );
  NAND2_X1 U351 ( .A1(G231GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U352 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U353 ( .A(n302), .B(n301), .Z(n308) );
  XNOR2_X1 U354 ( .A(G15GAT), .B(G1GAT), .ZN(n303) );
  XNOR2_X1 U355 ( .A(n303), .B(KEYINPUT73), .ZN(n361) );
  XOR2_X1 U356 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n305) );
  XNOR2_X1 U357 ( .A(KEYINPUT82), .B(KEYINPUT86), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U359 ( .A(n361), .B(n306), .ZN(n307) );
  XNOR2_X1 U360 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U361 ( .A(n310), .B(n309), .ZN(n573) );
  AND2_X1 U362 ( .A1(G230GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U363 ( .A(n314), .B(KEYINPUT33), .ZN(n320) );
  XOR2_X1 U364 ( .A(G120GAT), .B(G71GAT), .Z(n427) );
  XOR2_X1 U365 ( .A(n427), .B(G204GAT), .Z(n318) );
  XOR2_X1 U366 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n316) );
  XNOR2_X1 U367 ( .A(KEYINPUT79), .B(KEYINPUT78), .ZN(n315) );
  XOR2_X1 U368 ( .A(n316), .B(n315), .Z(n317) );
  XNOR2_X1 U369 ( .A(G106GAT), .B(G78GAT), .ZN(n321) );
  XNOR2_X1 U370 ( .A(n321), .B(G148GAT), .ZN(n443) );
  XNOR2_X1 U371 ( .A(G176GAT), .B(G92GAT), .ZN(n322) );
  XNOR2_X1 U372 ( .A(n322), .B(G64GAT), .ZN(n400) );
  XNOR2_X1 U373 ( .A(n443), .B(n400), .ZN(n323) );
  XNOR2_X1 U374 ( .A(n324), .B(n323), .ZN(n464) );
  XOR2_X1 U375 ( .A(n325), .B(G162GAT), .Z(n327) );
  XOR2_X1 U376 ( .A(G190GAT), .B(G134GAT), .Z(n430) );
  XNOR2_X1 U377 ( .A(n430), .B(G218GAT), .ZN(n326) );
  XNOR2_X1 U378 ( .A(n327), .B(n326), .ZN(n333) );
  XOR2_X1 U379 ( .A(KEYINPUT81), .B(KEYINPUT9), .Z(n329) );
  XNOR2_X1 U380 ( .A(G106GAT), .B(KEYINPUT80), .ZN(n328) );
  XOR2_X1 U381 ( .A(n329), .B(n328), .Z(n331) );
  NAND2_X1 U382 ( .A1(G232GAT), .A2(G233GAT), .ZN(n330) );
  XOR2_X1 U383 ( .A(KEYINPUT11), .B(KEYINPUT67), .Z(n335) );
  XNOR2_X1 U384 ( .A(G92GAT), .B(KEYINPUT10), .ZN(n334) );
  XNOR2_X1 U385 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U386 ( .A(n337), .B(n336), .ZN(n343) );
  XNOR2_X1 U387 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n338) );
  XNOR2_X1 U388 ( .A(n338), .B(G29GAT), .ZN(n339) );
  XOR2_X1 U389 ( .A(n339), .B(KEYINPUT7), .Z(n341) );
  XNOR2_X1 U390 ( .A(G43GAT), .B(G50GAT), .ZN(n340) );
  XNOR2_X1 U391 ( .A(n341), .B(n340), .ZN(n366) );
  INV_X1 U392 ( .A(n366), .ZN(n342) );
  INV_X1 U393 ( .A(n564), .ZN(n465) );
  XNOR2_X1 U394 ( .A(KEYINPUT36), .B(KEYINPUT103), .ZN(n344) );
  XNOR2_X1 U395 ( .A(n465), .B(n344), .ZN(n579) );
  NOR2_X1 U396 ( .A1(n573), .A2(n579), .ZN(n348) );
  XNOR2_X1 U397 ( .A(KEYINPUT114), .B(KEYINPUT45), .ZN(n346) );
  NOR2_X1 U398 ( .A1(n464), .A2(n349), .ZN(n367) );
  XOR2_X1 U399 ( .A(KEYINPUT68), .B(KEYINPUT29), .Z(n351) );
  XNOR2_X1 U400 ( .A(G113GAT), .B(G197GAT), .ZN(n350) );
  XNOR2_X1 U401 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U402 ( .A(KEYINPUT30), .B(KEYINPUT70), .Z(n353) );
  XNOR2_X1 U403 ( .A(KEYINPUT75), .B(KEYINPUT71), .ZN(n352) );
  XNOR2_X1 U404 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U405 ( .A(n355), .B(n354), .Z(n360) );
  XOR2_X1 U406 ( .A(KEYINPUT74), .B(KEYINPUT69), .Z(n357) );
  NAND2_X1 U407 ( .A1(G229GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U408 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U409 ( .A(KEYINPUT72), .B(n358), .ZN(n359) );
  XNOR2_X1 U410 ( .A(n360), .B(n359), .ZN(n362) );
  XOR2_X1 U411 ( .A(n362), .B(n361), .Z(n364) );
  XOR2_X1 U412 ( .A(G141GAT), .B(G22GAT), .Z(n438) );
  XOR2_X1 U413 ( .A(G169GAT), .B(G8GAT), .Z(n401) );
  XNOR2_X1 U414 ( .A(n438), .B(n401), .ZN(n363) );
  XNOR2_X1 U415 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U416 ( .A(n366), .B(n365), .Z(n503) );
  INV_X1 U417 ( .A(n503), .ZN(n569) );
  XNOR2_X1 U418 ( .A(KEYINPUT76), .B(n569), .ZN(n555) );
  NAND2_X1 U419 ( .A1(n367), .A2(n555), .ZN(n376) );
  XNOR2_X1 U420 ( .A(n464), .B(KEYINPUT64), .ZN(n368) );
  XNOR2_X1 U421 ( .A(n368), .B(KEYINPUT41), .ZN(n559) );
  NOR2_X1 U422 ( .A1(n569), .A2(n559), .ZN(n370) );
  XOR2_X1 U423 ( .A(KEYINPUT112), .B(KEYINPUT46), .Z(n369) );
  XNOR2_X1 U424 ( .A(n370), .B(n369), .ZN(n372) );
  AND2_X1 U425 ( .A1(n564), .A2(n573), .ZN(n371) );
  NAND2_X1 U426 ( .A1(n372), .A2(n371), .ZN(n374) );
  AND2_X1 U427 ( .A1(n376), .A2(n375), .ZN(n377) );
  XNOR2_X1 U428 ( .A(n377), .B(KEYINPUT48), .ZN(n453) );
  XOR2_X1 U429 ( .A(KEYINPUT6), .B(KEYINPUT93), .Z(n379) );
  XNOR2_X1 U430 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n378) );
  XNOR2_X1 U431 ( .A(n379), .B(n378), .ZN(n383) );
  XOR2_X1 U432 ( .A(KEYINPUT95), .B(KEYINPUT5), .Z(n381) );
  XNOR2_X1 U433 ( .A(G57GAT), .B(KEYINPUT96), .ZN(n380) );
  XNOR2_X1 U434 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U435 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U436 ( .A(G148GAT), .B(G120GAT), .Z(n385) );
  XNOR2_X1 U437 ( .A(G29GAT), .B(G141GAT), .ZN(n384) );
  XNOR2_X1 U438 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U439 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U440 ( .A(n388), .B(KEYINPUT1), .Z(n392) );
  XOR2_X1 U441 ( .A(G127GAT), .B(KEYINPUT0), .Z(n390) );
  XNOR2_X1 U442 ( .A(G113GAT), .B(KEYINPUT87), .ZN(n389) );
  XNOR2_X1 U443 ( .A(n390), .B(n389), .ZN(n429) );
  XNOR2_X1 U444 ( .A(n429), .B(KEYINPUT94), .ZN(n391) );
  XNOR2_X1 U445 ( .A(n392), .B(n391), .ZN(n399) );
  XOR2_X1 U446 ( .A(G155GAT), .B(KEYINPUT2), .Z(n394) );
  XNOR2_X1 U447 ( .A(G162GAT), .B(KEYINPUT3), .ZN(n393) );
  XNOR2_X1 U448 ( .A(n394), .B(n393), .ZN(n439) );
  XOR2_X1 U449 ( .A(G85GAT), .B(n439), .Z(n396) );
  NAND2_X1 U450 ( .A1(G225GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U451 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U452 ( .A(G134GAT), .B(n397), .Z(n398) );
  XNOR2_X1 U453 ( .A(n399), .B(n398), .ZN(n506) );
  INV_X1 U454 ( .A(n506), .ZN(n523) );
  XOR2_X1 U455 ( .A(n401), .B(n400), .Z(n403) );
  NAND2_X1 U456 ( .A1(G226GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U457 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U458 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n405) );
  XNOR2_X1 U459 ( .A(G36GAT), .B(G190GAT), .ZN(n404) );
  XNOR2_X1 U460 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U461 ( .A(n407), .B(n406), .Z(n416) );
  XOR2_X1 U462 ( .A(KEYINPUT89), .B(KEYINPUT18), .Z(n409) );
  XNOR2_X1 U463 ( .A(KEYINPUT19), .B(G183GAT), .ZN(n408) );
  XNOR2_X1 U464 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U465 ( .A(KEYINPUT17), .B(n410), .Z(n424) );
  XNOR2_X1 U466 ( .A(G211GAT), .B(G218GAT), .ZN(n411) );
  XNOR2_X1 U467 ( .A(n411), .B(KEYINPUT90), .ZN(n412) );
  XOR2_X1 U468 ( .A(n412), .B(KEYINPUT21), .Z(n414) );
  XNOR2_X1 U469 ( .A(G197GAT), .B(G204GAT), .ZN(n413) );
  XNOR2_X1 U470 ( .A(n414), .B(n413), .ZN(n437) );
  XNOR2_X1 U471 ( .A(n424), .B(n437), .ZN(n415) );
  XNOR2_X1 U472 ( .A(n416), .B(n415), .ZN(n509) );
  XOR2_X1 U473 ( .A(n509), .B(KEYINPUT27), .Z(n469) );
  NAND2_X1 U474 ( .A1(n523), .A2(n469), .ZN(n473) );
  NOR2_X1 U475 ( .A1(n453), .A2(n473), .ZN(n417) );
  XOR2_X1 U476 ( .A(KEYINPUT115), .B(n417), .Z(n541) );
  XOR2_X1 U477 ( .A(G176GAT), .B(KEYINPUT88), .Z(n419) );
  NAND2_X1 U478 ( .A1(G227GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U479 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U480 ( .A(KEYINPUT20), .B(G99GAT), .Z(n421) );
  XNOR2_X1 U481 ( .A(G43GAT), .B(G15GAT), .ZN(n420) );
  XNOR2_X1 U482 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U483 ( .A(n423), .B(n422), .Z(n426) );
  XNOR2_X1 U484 ( .A(G169GAT), .B(n424), .ZN(n425) );
  XNOR2_X1 U485 ( .A(n426), .B(n425), .ZN(n428) );
  XOR2_X1 U486 ( .A(n428), .B(n427), .Z(n432) );
  XNOR2_X1 U487 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U488 ( .A(n432), .B(n431), .ZN(n553) );
  NAND2_X1 U489 ( .A1(n541), .A2(n553), .ZN(n433) );
  XNOR2_X1 U490 ( .A(n433), .B(KEYINPUT116), .ZN(n448) );
  XOR2_X1 U491 ( .A(KEYINPUT23), .B(KEYINPUT92), .Z(n435) );
  XNOR2_X1 U492 ( .A(G50GAT), .B(KEYINPUT91), .ZN(n434) );
  XNOR2_X1 U493 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U494 ( .A(n437), .B(n436), .ZN(n447) );
  XOR2_X1 U495 ( .A(n439), .B(n438), .Z(n441) );
  NAND2_X1 U496 ( .A1(G228GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U497 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U498 ( .A(n442), .B(KEYINPUT24), .Z(n445) );
  XNOR2_X1 U499 ( .A(n443), .B(KEYINPUT22), .ZN(n444) );
  XNOR2_X1 U500 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U501 ( .A(n447), .B(n446), .ZN(n551) );
  XOR2_X1 U502 ( .A(n551), .B(KEYINPUT28), .Z(n529) );
  NOR2_X1 U503 ( .A1(n448), .A2(n529), .ZN(n449) );
  XNOR2_X1 U504 ( .A(n449), .B(KEYINPUT117), .ZN(n536) );
  NOR2_X1 U505 ( .A1(n573), .A2(n536), .ZN(n452) );
  INV_X1 U506 ( .A(G127GAT), .ZN(n450) );
  XNOR2_X1 U507 ( .A(n452), .B(n451), .ZN(G1342GAT) );
  INV_X1 U508 ( .A(KEYINPUT123), .ZN(n459) );
  NOR2_X1 U509 ( .A1(n509), .A2(n453), .ZN(n454) );
  XNOR2_X1 U510 ( .A(n454), .B(KEYINPUT54), .ZN(n455) );
  NAND2_X1 U511 ( .A1(n455), .A2(n506), .ZN(n456) );
  XNOR2_X1 U512 ( .A(n456), .B(KEYINPUT65), .ZN(n550) );
  NOR2_X1 U513 ( .A1(n551), .A2(n553), .ZN(n457) );
  XNOR2_X1 U514 ( .A(n457), .B(KEYINPUT26), .ZN(n540) );
  NAND2_X1 U515 ( .A1(n550), .A2(n540), .ZN(n458) );
  XNOR2_X1 U516 ( .A(n459), .B(n458), .ZN(n578) );
  INV_X1 U517 ( .A(n578), .ZN(n460) );
  NAND2_X1 U518 ( .A1(n460), .A2(n464), .ZN(n463) );
  XOR2_X1 U519 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n461) );
  NOR2_X1 U520 ( .A1(n555), .A2(n464), .ZN(n493) );
  NOR2_X1 U521 ( .A1(n573), .A2(n465), .ZN(n466) );
  XNOR2_X1 U522 ( .A(KEYINPUT16), .B(n466), .ZN(n477) );
  INV_X1 U523 ( .A(n509), .ZN(n525) );
  NAND2_X1 U524 ( .A1(n553), .A2(n525), .ZN(n467) );
  NAND2_X1 U525 ( .A1(n551), .A2(n467), .ZN(n468) );
  XOR2_X1 U526 ( .A(KEYINPUT25), .B(n468), .Z(n471) );
  NAND2_X1 U527 ( .A1(n469), .A2(n540), .ZN(n470) );
  NAND2_X1 U528 ( .A1(n471), .A2(n470), .ZN(n472) );
  NAND2_X1 U529 ( .A1(n472), .A2(n506), .ZN(n476) );
  NOR2_X1 U530 ( .A1(n529), .A2(n473), .ZN(n474) );
  INV_X1 U531 ( .A(n553), .ZN(n513) );
  NAND2_X1 U532 ( .A1(n474), .A2(n513), .ZN(n475) );
  NAND2_X1 U533 ( .A1(n476), .A2(n475), .ZN(n488) );
  AND2_X1 U534 ( .A1(n477), .A2(n488), .ZN(n505) );
  NAND2_X1 U535 ( .A1(n493), .A2(n505), .ZN(n485) );
  NOR2_X1 U536 ( .A1(n506), .A2(n485), .ZN(n479) );
  XNOR2_X1 U537 ( .A(KEYINPUT99), .B(KEYINPUT34), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U539 ( .A(G1GAT), .B(n480), .ZN(G1324GAT) );
  NOR2_X1 U540 ( .A1(n509), .A2(n485), .ZN(n481) );
  XOR2_X1 U541 ( .A(G8GAT), .B(n481), .Z(G1325GAT) );
  NOR2_X1 U542 ( .A1(n513), .A2(n485), .ZN(n483) );
  XNOR2_X1 U543 ( .A(KEYINPUT100), .B(KEYINPUT35), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U545 ( .A(G15GAT), .B(n484), .ZN(G1326GAT) );
  INV_X1 U546 ( .A(n529), .ZN(n517) );
  NOR2_X1 U547 ( .A1(n517), .A2(n485), .ZN(n487) );
  XNOR2_X1 U548 ( .A(G22GAT), .B(KEYINPUT101), .ZN(n486) );
  XNOR2_X1 U549 ( .A(n487), .B(n486), .ZN(G1327GAT) );
  NAND2_X1 U550 ( .A1(n573), .A2(n488), .ZN(n489) );
  XNOR2_X1 U551 ( .A(KEYINPUT104), .B(n489), .ZN(n490) );
  NOR2_X1 U552 ( .A1(n579), .A2(n490), .ZN(n492) );
  XNOR2_X1 U553 ( .A(KEYINPUT37), .B(KEYINPUT105), .ZN(n491) );
  XNOR2_X1 U554 ( .A(n492), .B(n491), .ZN(n520) );
  NAND2_X1 U555 ( .A1(n520), .A2(n493), .ZN(n494) );
  XNOR2_X1 U556 ( .A(KEYINPUT38), .B(n494), .ZN(n501) );
  NOR2_X1 U557 ( .A1(n501), .A2(n506), .ZN(n496) );
  XNOR2_X1 U558 ( .A(KEYINPUT102), .B(KEYINPUT39), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U560 ( .A(G29GAT), .B(n497), .ZN(G1328GAT) );
  NOR2_X1 U561 ( .A1(n509), .A2(n501), .ZN(n498) );
  XOR2_X1 U562 ( .A(G36GAT), .B(n498), .Z(G1329GAT) );
  NOR2_X1 U563 ( .A1(n501), .A2(n513), .ZN(n499) );
  XOR2_X1 U564 ( .A(KEYINPUT40), .B(n499), .Z(n500) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(n500), .ZN(G1330GAT) );
  NOR2_X1 U566 ( .A1(n501), .A2(n517), .ZN(n502) );
  XOR2_X1 U567 ( .A(G50GAT), .B(n502), .Z(G1331GAT) );
  NOR2_X1 U568 ( .A1(n559), .A2(n503), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n504), .B(KEYINPUT106), .ZN(n521) );
  NAND2_X1 U570 ( .A1(n505), .A2(n521), .ZN(n516) );
  NOR2_X1 U571 ( .A1(n506), .A2(n516), .ZN(n507) );
  XOR2_X1 U572 ( .A(G57GAT), .B(n507), .Z(n508) );
  XNOR2_X1 U573 ( .A(KEYINPUT42), .B(n508), .ZN(G1332GAT) );
  NOR2_X1 U574 ( .A1(n509), .A2(n516), .ZN(n511) );
  XNOR2_X1 U575 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U577 ( .A(G64GAT), .B(n512), .ZN(G1333GAT) );
  NOR2_X1 U578 ( .A1(n513), .A2(n516), .ZN(n515) );
  XNOR2_X1 U579 ( .A(G71GAT), .B(KEYINPUT109), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(G1334GAT) );
  NOR2_X1 U581 ( .A1(n517), .A2(n516), .ZN(n519) );
  XNOR2_X1 U582 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  NAND2_X1 U584 ( .A1(n521), .A2(n520), .ZN(n522) );
  XOR2_X1 U585 ( .A(KEYINPUT110), .B(n522), .Z(n530) );
  NAND2_X1 U586 ( .A1(n523), .A2(n530), .ZN(n524) );
  XNOR2_X1 U587 ( .A(G85GAT), .B(n524), .ZN(G1336GAT) );
  NAND2_X1 U588 ( .A1(n530), .A2(n525), .ZN(n526) );
  XNOR2_X1 U589 ( .A(n526), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U590 ( .A(G99GAT), .B(KEYINPUT111), .Z(n528) );
  NAND2_X1 U591 ( .A1(n553), .A2(n530), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n528), .B(n527), .ZN(G1338GAT) );
  NAND2_X1 U593 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U594 ( .A(n531), .B(KEYINPUT44), .ZN(n532) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n532), .ZN(G1339GAT) );
  NOR2_X1 U596 ( .A1(n555), .A2(n536), .ZN(n533) );
  XOR2_X1 U597 ( .A(G113GAT), .B(n533), .Z(G1340GAT) );
  NOR2_X1 U598 ( .A1(n559), .A2(n536), .ZN(n535) );
  XNOR2_X1 U599 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n535), .B(n534), .ZN(G1341GAT) );
  NOR2_X1 U601 ( .A1(n564), .A2(n536), .ZN(n538) );
  XNOR2_X1 U602 ( .A(KEYINPUT118), .B(KEYINPUT51), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U604 ( .A(G134GAT), .B(n539), .ZN(G1343GAT) );
  NAND2_X1 U605 ( .A1(n541), .A2(n540), .ZN(n548) );
  NOR2_X1 U606 ( .A1(n569), .A2(n548), .ZN(n542) );
  XOR2_X1 U607 ( .A(G141GAT), .B(n542), .Z(G1344GAT) );
  NOR2_X1 U608 ( .A1(n548), .A2(n559), .ZN(n546) );
  XOR2_X1 U609 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n544) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT119), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(G1345GAT) );
  NOR2_X1 U613 ( .A1(n573), .A2(n548), .ZN(n547) );
  XOR2_X1 U614 ( .A(G155GAT), .B(n547), .Z(G1346GAT) );
  NOR2_X1 U615 ( .A1(n564), .A2(n548), .ZN(n549) );
  XOR2_X1 U616 ( .A(G162GAT), .B(n549), .Z(G1347GAT) );
  NAND2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n552), .B(KEYINPUT55), .ZN(n554) );
  NAND2_X1 U619 ( .A1(n554), .A2(n553), .ZN(n565) );
  NOR2_X1 U620 ( .A1(n555), .A2(n565), .ZN(n556) );
  XOR2_X1 U621 ( .A(G169GAT), .B(n556), .Z(G1348GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT120), .B(KEYINPUT56), .Z(n558) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(n561) );
  NOR2_X1 U625 ( .A1(n559), .A2(n565), .ZN(n560) );
  XOR2_X1 U626 ( .A(n561), .B(n560), .Z(G1349GAT) );
  NOR2_X1 U627 ( .A1(n573), .A2(n565), .ZN(n563) );
  XNOR2_X1 U628 ( .A(G183GAT), .B(KEYINPUT121), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1350GAT) );
  NOR2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n567) );
  XNOR2_X1 U631 ( .A(KEYINPUT122), .B(KEYINPUT58), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n568) );
  XOR2_X1 U633 ( .A(G190GAT), .B(n568), .Z(G1351GAT) );
  NOR2_X1 U634 ( .A1(n569), .A2(n578), .ZN(n571) );
  XNOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(n572), .ZN(G1352GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n578), .ZN(n575) );
  XNOR2_X1 U639 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1354GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n577) );
  XNOR2_X1 U642 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n581) );
  NOR2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U645 ( .A(n581), .B(n580), .Z(G1355GAT) );
endmodule

