

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752;

  XNOR2_X1 U364 ( .A(n535), .B(n456), .ZN(n545) );
  OR2_X2 U365 ( .A1(n739), .A2(G902), .ZN(n378) );
  BUF_X1 U366 ( .A(n618), .Z(n341) );
  XNOR2_X2 U367 ( .A(n489), .B(n488), .ZN(n542) );
  XNOR2_X2 U368 ( .A(n744), .B(n380), .ZN(n358) );
  XNOR2_X2 U369 ( .A(n491), .B(n448), .ZN(n744) );
  XNOR2_X2 U370 ( .A(n469), .B(n423), .ZN(n743) );
  XNOR2_X2 U371 ( .A(n449), .B(G125), .ZN(n469) );
  XNOR2_X2 U372 ( .A(n631), .B(KEYINPUT38), .ZN(n716) );
  BUF_X2 U373 ( .A(n538), .Z(n631) );
  AND2_X1 U374 ( .A1(n643), .A2(n642), .ZN(n729) );
  NAND2_X1 U375 ( .A1(n401), .A2(n403), .ZN(n385) );
  NAND2_X1 U376 ( .A1(n398), .A2(n397), .ZN(n400) );
  NAND2_X1 U377 ( .A1(n396), .A2(n395), .ZN(n745) );
  XNOR2_X1 U378 ( .A(n557), .B(n556), .ZN(n671) );
  AND2_X1 U379 ( .A1(n612), .A2(n698), .ZN(n693) );
  NAND2_X1 U380 ( .A1(n390), .A2(n349), .ZN(n557) );
  XNOR2_X1 U381 ( .A(n621), .B(n354), .ZN(n622) );
  XNOR2_X1 U382 ( .A(n544), .B(n543), .ZN(n568) );
  NOR2_X1 U383 ( .A1(n608), .A2(n607), .ZN(n627) );
  XNOR2_X1 U384 ( .A(n413), .B(n479), .ZN(n538) );
  OR2_X1 U385 ( .A1(n679), .A2(G902), .ZN(n455) );
  XNOR2_X1 U386 ( .A(n433), .B(n432), .ZN(n490) );
  XNOR2_X1 U387 ( .A(G101), .B(G113), .ZN(n366) );
  NOR2_X1 U388 ( .A1(n527), .A2(n528), .ZN(n529) );
  XNOR2_X1 U389 ( .A(G902), .B(KEYINPUT93), .ZN(n437) );
  XNOR2_X1 U390 ( .A(KEYINPUT73), .B(G131), .ZN(n506) );
  INV_X1 U391 ( .A(G237), .ZN(n478) );
  XOR2_X1 U392 ( .A(KEYINPUT8), .B(KEYINPUT72), .Z(n432) );
  XNOR2_X1 U393 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U394 ( .A(n421), .B(n419), .ZN(n517) );
  NOR2_X1 U395 ( .A1(n752), .A2(n645), .ZN(n394) );
  XNOR2_X1 U396 ( .A(KEYINPUT79), .B(n458), .ZN(n511) );
  NOR2_X1 U397 ( .A1(G953), .A2(G237), .ZN(n457) );
  INV_X1 U398 ( .A(KEYINPUT112), .ZN(n383) );
  XNOR2_X1 U399 ( .A(G143), .B(G128), .ZN(n468) );
  XNOR2_X1 U400 ( .A(KEYINPUT4), .B(G137), .ZN(n447) );
  INV_X1 U401 ( .A(n729), .ZN(n397) );
  NAND2_X1 U402 ( .A1(G234), .A2(G237), .ZN(n482) );
  INV_X1 U403 ( .A(KEYINPUT30), .ZN(n405) );
  AND2_X1 U404 ( .A1(n536), .A2(n697), .ZN(n377) );
  OR2_X1 U405 ( .A1(n657), .A2(n644), .ZN(n413) );
  NOR2_X1 U406 ( .A1(n650), .A2(G902), .ZN(n464) );
  XNOR2_X1 U407 ( .A(n542), .B(KEYINPUT96), .ZN(n554) );
  INV_X1 U408 ( .A(n752), .ZN(n395) );
  XNOR2_X1 U409 ( .A(n365), .B(n363), .ZN(n467) );
  XNOR2_X1 U410 ( .A(n364), .B(KEYINPUT3), .ZN(n363) );
  XNOR2_X1 U411 ( .A(n367), .B(n366), .ZN(n365) );
  XNOR2_X1 U412 ( .A(G119), .B(G116), .ZN(n364) );
  XNOR2_X1 U413 ( .A(n429), .B(n428), .ZN(n427) );
  XNOR2_X1 U414 ( .A(G119), .B(KEYINPUT97), .ZN(n429) );
  XNOR2_X1 U415 ( .A(KEYINPUT23), .B(G110), .ZN(n428) );
  XNOR2_X1 U416 ( .A(n426), .B(KEYINPUT24), .ZN(n425) );
  XNOR2_X1 U417 ( .A(G128), .B(G137), .ZN(n426) );
  XNOR2_X1 U418 ( .A(KEYINPUT10), .B(G140), .ZN(n423) );
  XNOR2_X1 U419 ( .A(G101), .B(KEYINPUT83), .ZN(n368) );
  INV_X1 U420 ( .A(G146), .ZN(n380) );
  XNOR2_X1 U421 ( .A(n362), .B(G104), .ZN(n466) );
  XNOR2_X1 U422 ( .A(G110), .B(G107), .ZN(n362) );
  INV_X1 U423 ( .A(KEYINPUT88), .ZN(n404) );
  XNOR2_X1 U424 ( .A(n372), .B(KEYINPUT33), .ZN(n733) );
  NAND2_X1 U425 ( .A1(n399), .A2(n371), .ZN(n372) );
  NOR2_X1 U426 ( .A1(n565), .A2(n344), .ZN(n399) );
  NAND2_X1 U427 ( .A1(n370), .A2(n369), .ZN(n371) );
  XNOR2_X1 U428 ( .A(n417), .B(KEYINPUT41), .ZN(n732) );
  XNOR2_X1 U429 ( .A(n592), .B(KEYINPUT39), .ZN(n593) );
  NAND2_X1 U430 ( .A1(n591), .A2(n590), .ZN(n592) );
  BUF_X1 U431 ( .A(n526), .Z(n549) );
  XNOR2_X1 U432 ( .A(n519), .B(n518), .ZN(n537) );
  INV_X1 U433 ( .A(KEYINPUT64), .ZN(n431) );
  XNOR2_X1 U434 ( .A(n467), .B(n359), .ZN(n581) );
  XNOR2_X1 U435 ( .A(n466), .B(n360), .ZN(n359) );
  XNOR2_X1 U436 ( .A(n465), .B(n361), .ZN(n360) );
  INV_X1 U437 ( .A(G122), .ZN(n361) );
  NOR2_X1 U438 ( .A1(n693), .A2(n614), .ZN(n615) );
  AND2_X1 U439 ( .A1(n342), .A2(n603), .ZN(n604) );
  XNOR2_X1 U440 ( .A(n533), .B(KEYINPUT86), .ZN(n596) );
  XNOR2_X1 U441 ( .A(KEYINPUT75), .B(KEYINPUT76), .ZN(n367) );
  XNOR2_X1 U442 ( .A(G143), .B(G104), .ZN(n512) );
  XNOR2_X1 U443 ( .A(n743), .B(n422), .ZN(n421) );
  XNOR2_X1 U444 ( .A(n509), .B(n507), .ZN(n422) );
  BUF_X1 U445 ( .A(n506), .Z(n509) );
  XNOR2_X1 U446 ( .A(n508), .B(n420), .ZN(n419) );
  XNOR2_X1 U447 ( .A(n510), .B(KEYINPUT99), .ZN(n420) );
  XNOR2_X1 U448 ( .A(KEYINPUT12), .B(KEYINPUT103), .ZN(n510) );
  NAND2_X1 U449 ( .A1(n393), .A2(n392), .ZN(n398) );
  NAND2_X1 U450 ( .A1(n415), .A2(KEYINPUT2), .ZN(n392) );
  NOR2_X1 U451 ( .A1(n745), .A2(n638), .ZN(n641) );
  XNOR2_X1 U452 ( .A(KEYINPUT4), .B(KEYINPUT18), .ZN(n470) );
  OR2_X1 U453 ( .A1(n545), .A2(n552), .ZN(n370) );
  NAND2_X1 U454 ( .A1(n345), .A2(n545), .ZN(n369) );
  INV_X1 U455 ( .A(G902), .ZN(n501) );
  XNOR2_X1 U456 ( .A(n387), .B(n574), .ZN(n643) );
  INV_X1 U457 ( .A(G134), .ZN(n443) );
  XNOR2_X1 U458 ( .A(G116), .B(G107), .ZN(n495) );
  INV_X1 U459 ( .A(KEYINPUT80), .ZN(n424) );
  XNOR2_X1 U460 ( .A(n406), .B(n405), .ZN(n376) );
  XNOR2_X1 U461 ( .A(n481), .B(n355), .ZN(n486) );
  NOR2_X1 U462 ( .A1(n598), .A2(n703), .ZN(n599) );
  NAND2_X1 U463 ( .A1(n554), .A2(n524), .ZN(n416) );
  BUF_X1 U464 ( .A(n545), .Z(n698) );
  XNOR2_X1 U465 ( .A(n462), .B(n358), .ZN(n650) );
  XNOR2_X1 U466 ( .A(n379), .B(n435), .ZN(n739) );
  XNOR2_X1 U467 ( .A(n434), .B(n743), .ZN(n379) );
  XNOR2_X1 U468 ( .A(n427), .B(n425), .ZN(n434) );
  XNOR2_X1 U469 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U470 ( .A(n452), .B(n374), .ZN(n373) );
  INV_X1 U471 ( .A(n466), .ZN(n374) );
  XNOR2_X1 U472 ( .A(n657), .B(n656), .ZN(n658) );
  OR2_X1 U473 ( .A1(n527), .A2(G952), .ZN(n676) );
  OR2_X1 U474 ( .A1(n734), .A2(n356), .ZN(n389) );
  XNOR2_X1 U475 ( .A(n637), .B(KEYINPUT117), .ZN(n752) );
  XNOR2_X1 U476 ( .A(n391), .B(n353), .ZN(n390) );
  INV_X1 U477 ( .A(n416), .ZN(n683) );
  XNOR2_X1 U478 ( .A(n622), .B(G137), .ZN(G39) );
  AND2_X1 U479 ( .A1(n350), .A2(n486), .ZN(n342) );
  XOR2_X1 U480 ( .A(n439), .B(n346), .Z(n343) );
  NAND2_X1 U481 ( .A1(n381), .A2(n382), .ZN(n403) );
  INV_X1 U482 ( .A(G146), .ZN(n449) );
  NOR2_X1 U483 ( .A1(n697), .A2(KEYINPUT113), .ZN(n344) );
  NAND2_X1 U484 ( .A1(n697), .A2(KEYINPUT113), .ZN(n345) );
  XNOR2_X1 U485 ( .A(KEYINPUT82), .B(KEYINPUT25), .ZN(n346) );
  AND2_X1 U486 ( .A1(n731), .A2(n403), .ZN(n347) );
  XOR2_X1 U487 ( .A(n485), .B(KEYINPUT95), .Z(n348) );
  NOR2_X1 U488 ( .A1(n341), .A2(n619), .ZN(n349) );
  AND2_X1 U489 ( .A1(n745), .A2(n642), .ZN(n728) );
  AND2_X1 U490 ( .A1(n601), .A2(n600), .ZN(n350) );
  NOR2_X1 U491 ( .A1(n341), .A2(n537), .ZN(n351) );
  NAND2_X1 U492 ( .A1(n341), .A2(n714), .ZN(n352) );
  XOR2_X1 U493 ( .A(n555), .B(KEYINPUT34), .Z(n353) );
  XOR2_X1 U494 ( .A(n620), .B(KEYINPUT42), .Z(n354) );
  XOR2_X1 U495 ( .A(KEYINPUT81), .B(KEYINPUT19), .Z(n355) );
  AND2_X1 U496 ( .A1(n733), .A2(n732), .ZN(n356) );
  AND2_X1 U497 ( .A1(n640), .A2(n639), .ZN(n357) );
  INV_X1 U498 ( .A(n645), .ZN(n415) );
  XNOR2_X1 U499 ( .A(n358), .B(n373), .ZN(n679) );
  XNOR2_X1 U500 ( .A(n368), .B(G140), .ZN(n450) );
  XNOR2_X2 U501 ( .A(n375), .B(n424), .ZN(n591) );
  NAND2_X1 U502 ( .A1(n377), .A2(n376), .ZN(n375) );
  XNOR2_X2 U503 ( .A(n378), .B(n343), .ZN(n701) );
  XNOR2_X1 U504 ( .A(n648), .B(n404), .ZN(n381) );
  NAND2_X1 U505 ( .A1(n382), .A2(n640), .ZN(n638) );
  INV_X1 U506 ( .A(n643), .ZN(n382) );
  XNOR2_X1 U507 ( .A(n384), .B(n383), .ZN(n571) );
  NAND2_X1 U508 ( .A1(n569), .A2(n587), .ZN(n384) );
  XNOR2_X2 U509 ( .A(n385), .B(KEYINPUT65), .ZN(n672) );
  XNOR2_X2 U510 ( .A(n386), .B(KEYINPUT31), .ZN(n561) );
  NAND2_X1 U511 ( .A1(n542), .A2(n708), .ZN(n386) );
  NAND2_X1 U512 ( .A1(n572), .A2(n573), .ZN(n387) );
  NAND2_X1 U513 ( .A1(n486), .A2(n348), .ZN(n489) );
  XNOR2_X1 U514 ( .A(n388), .B(n625), .ZN(n634) );
  NAND2_X1 U515 ( .A1(n412), .A2(n624), .ZN(n388) );
  NAND2_X1 U516 ( .A1(n402), .A2(n400), .ZN(n401) );
  NOR2_X1 U517 ( .A1(n347), .A2(n389), .ZN(n735) );
  INV_X1 U518 ( .A(n617), .ZN(n408) );
  XNOR2_X2 U519 ( .A(n595), .B(n594), .ZN(n617) );
  NAND2_X1 U520 ( .A1(n733), .A2(n554), .ZN(n391) );
  NAND2_X1 U521 ( .A1(n396), .A2(n394), .ZN(n393) );
  INV_X1 U522 ( .A(n646), .ZN(n396) );
  NAND2_X1 U523 ( .A1(n545), .A2(n697), .ZN(n553) );
  NOR2_X1 U524 ( .A1(n641), .A2(n357), .ZN(n402) );
  NAND2_X1 U525 ( .A1(n526), .A2(n714), .ZN(n406) );
  NAND2_X1 U526 ( .A1(n407), .A2(n623), .ZN(n411) );
  NAND2_X1 U527 ( .A1(n408), .A2(n622), .ZN(n407) );
  NAND2_X1 U528 ( .A1(n411), .A2(n409), .ZN(n412) );
  NAND2_X1 U529 ( .A1(n410), .A2(n622), .ZN(n409) );
  NOR2_X1 U530 ( .A1(n617), .A2(n623), .ZN(n410) );
  XNOR2_X1 U531 ( .A(n414), .B(n581), .ZN(n657) );
  XNOR2_X1 U532 ( .A(n476), .B(n475), .ZN(n414) );
  NAND2_X1 U533 ( .A1(n562), .A2(n416), .ZN(n563) );
  NAND2_X1 U534 ( .A1(n350), .A2(n732), .ZN(n621) );
  NAND2_X1 U535 ( .A1(n418), .A2(n619), .ZN(n417) );
  NOR2_X1 U536 ( .A1(n716), .A2(n352), .ZN(n418) );
  NAND2_X1 U537 ( .A1(n593), .A2(n351), .ZN(n637) );
  INV_X1 U538 ( .A(n591), .ZN(n589) );
  NOR2_X1 U539 ( .A1(n546), .A2(n606), .ZN(n430) );
  INV_X1 U540 ( .A(n561), .ZN(n562) );
  INV_X1 U541 ( .A(n613), .ZN(n614) );
  AND2_X1 U542 ( .A1(n616), .A2(n615), .ZN(n624) );
  INV_X1 U543 ( .A(G472), .ZN(n463) );
  NAND2_X1 U544 ( .A1(n446), .A2(n445), .ZN(n491) );
  XNOR2_X2 U545 ( .A(n431), .B(G953), .ZN(n527) );
  NAND2_X1 U546 ( .A1(G234), .A2(n527), .ZN(n433) );
  NAND2_X1 U547 ( .A1(G221), .A2(n490), .ZN(n435) );
  INV_X1 U548 ( .A(KEYINPUT15), .ZN(n436) );
  XNOR2_X1 U549 ( .A(n437), .B(n436), .ZN(n477) );
  NAND2_X1 U550 ( .A1(n477), .A2(G234), .ZN(n438) );
  XNOR2_X1 U551 ( .A(n438), .B(KEYINPUT20), .ZN(n440) );
  NAND2_X1 U552 ( .A1(n440), .A2(G217), .ZN(n439) );
  NAND2_X1 U553 ( .A1(G221), .A2(n440), .ZN(n442) );
  INV_X1 U554 ( .A(KEYINPUT21), .ZN(n441) );
  XNOR2_X1 U555 ( .A(n442), .B(n441), .ZN(n700) );
  AND2_X2 U556 ( .A1(n701), .A2(n700), .ZN(n697) );
  NAND2_X1 U557 ( .A1(n468), .A2(n443), .ZN(n446) );
  XOR2_X1 U558 ( .A(G143), .B(G128), .Z(n444) );
  NAND2_X1 U559 ( .A1(n444), .A2(G134), .ZN(n445) );
  XNOR2_X1 U560 ( .A(n506), .B(n447), .ZN(n448) );
  NAND2_X1 U561 ( .A1(n527), .A2(G227), .ZN(n451) );
  XNOR2_X1 U562 ( .A(n451), .B(n450), .ZN(n452) );
  INV_X1 U563 ( .A(KEYINPUT74), .ZN(n453) );
  XNOR2_X1 U564 ( .A(n453), .B(G469), .ZN(n454) );
  XNOR2_X2 U565 ( .A(n455), .B(n454), .ZN(n535) );
  INV_X1 U566 ( .A(KEYINPUT1), .ZN(n456) );
  INV_X1 U567 ( .A(n457), .ZN(n458) );
  NAND2_X1 U568 ( .A1(n511), .A2(G210), .ZN(n460) );
  XNOR2_X1 U569 ( .A(KEYINPUT98), .B(KEYINPUT5), .ZN(n459) );
  XNOR2_X1 U570 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U571 ( .A(n467), .B(n461), .ZN(n462) );
  XNOR2_X1 U572 ( .A(n464), .B(n463), .ZN(n526) );
  INV_X1 U573 ( .A(n549), .ZN(n703) );
  NOR2_X1 U574 ( .A1(n553), .A2(n703), .ZN(n708) );
  XNOR2_X1 U575 ( .A(KEYINPUT78), .B(KEYINPUT16), .ZN(n465) );
  XNOR2_X1 U576 ( .A(n469), .B(n468), .ZN(n472) );
  XNOR2_X1 U577 ( .A(n470), .B(KEYINPUT94), .ZN(n471) );
  XNOR2_X1 U578 ( .A(n472), .B(n471), .ZN(n476) );
  XOR2_X1 U579 ( .A(KEYINPUT17), .B(KEYINPUT84), .Z(n474) );
  NAND2_X1 U580 ( .A1(n527), .A2(G224), .ZN(n473) );
  XNOR2_X1 U581 ( .A(n474), .B(n473), .ZN(n475) );
  INV_X1 U582 ( .A(n477), .ZN(n644) );
  NAND2_X1 U583 ( .A1(n501), .A2(n478), .ZN(n480) );
  AND2_X1 U584 ( .A1(n480), .A2(G210), .ZN(n479) );
  NAND2_X1 U585 ( .A1(n480), .A2(G214), .ZN(n714) );
  NAND2_X1 U586 ( .A1(n538), .A2(n714), .ZN(n481) );
  XNOR2_X1 U587 ( .A(n482), .B(KEYINPUT14), .ZN(n483) );
  NAND2_X1 U588 ( .A1(G952), .A2(n483), .ZN(n727) );
  NOR2_X1 U589 ( .A1(G953), .A2(n727), .ZN(n531) );
  NAND2_X1 U590 ( .A1(G902), .A2(n483), .ZN(n528) );
  INV_X1 U591 ( .A(G898), .ZN(n577) );
  NAND2_X1 U592 ( .A1(G953), .A2(n577), .ZN(n582) );
  NOR2_X1 U593 ( .A1(n528), .A2(n582), .ZN(n484) );
  OR2_X1 U594 ( .A1(n531), .A2(n484), .ZN(n485) );
  XNOR2_X1 U595 ( .A(KEYINPUT91), .B(KEYINPUT0), .ZN(n487) );
  XNOR2_X1 U596 ( .A(n487), .B(KEYINPUT70), .ZN(n488) );
  NAND2_X1 U597 ( .A1(n490), .A2(G217), .ZN(n492) );
  XNOR2_X1 U598 ( .A(n492), .B(n491), .ZN(n500) );
  XOR2_X1 U599 ( .A(KEYINPUT9), .B(KEYINPUT108), .Z(n494) );
  XNOR2_X1 U600 ( .A(G122), .B(KEYINPUT106), .ZN(n493) );
  XNOR2_X1 U601 ( .A(n494), .B(n493), .ZN(n498) );
  XOR2_X1 U602 ( .A(KEYINPUT7), .B(KEYINPUT107), .Z(n496) );
  XNOR2_X1 U603 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U604 ( .A(n498), .B(n497), .Z(n499) );
  XNOR2_X1 U605 ( .A(n500), .B(n499), .ZN(n673) );
  NAND2_X1 U606 ( .A1(n673), .A2(n501), .ZN(n503) );
  INV_X1 U607 ( .A(G478), .ZN(n502) );
  XNOR2_X1 U608 ( .A(n503), .B(n502), .ZN(n618) );
  XOR2_X1 U609 ( .A(KEYINPUT105), .B(KEYINPUT13), .Z(n505) );
  XNOR2_X1 U610 ( .A(KEYINPUT104), .B(G475), .ZN(n504) );
  XNOR2_X1 U611 ( .A(n505), .B(n504), .ZN(n519) );
  XOR2_X1 U612 ( .A(KEYINPUT102), .B(KEYINPUT100), .Z(n508) );
  XNOR2_X1 U613 ( .A(G113), .B(G122), .ZN(n507) );
  NAND2_X1 U614 ( .A1(G214), .A2(n511), .ZN(n515) );
  XOR2_X1 U615 ( .A(KEYINPUT101), .B(KEYINPUT11), .Z(n513) );
  XNOR2_X1 U616 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U617 ( .A(n517), .B(n516), .ZN(n665) );
  NOR2_X1 U618 ( .A1(n665), .A2(G902), .ZN(n518) );
  NAND2_X1 U619 ( .A1(n561), .A2(n351), .ZN(n520) );
  XNOR2_X1 U620 ( .A(n520), .B(G116), .ZN(G18) );
  NAND2_X1 U621 ( .A1(n341), .A2(n537), .ZN(n521) );
  XNOR2_X2 U622 ( .A(n521), .B(KEYINPUT109), .ZN(n690) );
  NAND2_X1 U623 ( .A1(n561), .A2(n690), .ZN(n522) );
  XNOR2_X1 U624 ( .A(n522), .B(G113), .ZN(G15) );
  INV_X1 U625 ( .A(n535), .ZN(n600) );
  NAND2_X1 U626 ( .A1(n697), .A2(n600), .ZN(n523) );
  NOR2_X1 U627 ( .A1(n523), .A2(n549), .ZN(n524) );
  NAND2_X1 U628 ( .A1(n683), .A2(n690), .ZN(n525) );
  XNOR2_X1 U629 ( .A(n525), .B(G104), .ZN(G6) );
  XOR2_X1 U630 ( .A(KEYINPUT114), .B(n529), .Z(n530) );
  NOR2_X1 U631 ( .A1(G900), .A2(n530), .ZN(n532) );
  OR2_X1 U632 ( .A1(n532), .A2(n531), .ZN(n533) );
  INV_X1 U633 ( .A(n596), .ZN(n534) );
  NOR2_X1 U634 ( .A1(n535), .A2(n534), .ZN(n536) );
  INV_X1 U635 ( .A(n537), .ZN(n619) );
  NAND2_X1 U636 ( .A1(n349), .A2(n631), .ZN(n539) );
  OR2_X1 U637 ( .A1(n589), .A2(n539), .ZN(n613) );
  XNOR2_X1 U638 ( .A(n613), .B(G143), .ZN(G45) );
  AND2_X1 U639 ( .A1(n619), .A2(n341), .ZN(n717) );
  NAND2_X1 U640 ( .A1(n717), .A2(n700), .ZN(n540) );
  XNOR2_X1 U641 ( .A(n540), .B(KEYINPUT111), .ZN(n541) );
  NAND2_X1 U642 ( .A1(n542), .A2(n541), .ZN(n544) );
  XNOR2_X1 U643 ( .A(KEYINPUT66), .B(KEYINPUT22), .ZN(n543) );
  INV_X1 U644 ( .A(n568), .ZN(n547) );
  INV_X1 U645 ( .A(n701), .ZN(n626) );
  NAND2_X1 U646 ( .A1(n698), .A2(n626), .ZN(n546) );
  XNOR2_X1 U647 ( .A(n549), .B(KEYINPUT6), .ZN(n565) );
  INV_X1 U648 ( .A(n565), .ZN(n606) );
  NAND2_X1 U649 ( .A1(n547), .A2(n430), .ZN(n548) );
  XNOR2_X1 U650 ( .A(n548), .B(KEYINPUT32), .ZN(n588) );
  INV_X1 U651 ( .A(n698), .ZN(n628) );
  NOR2_X1 U652 ( .A1(n701), .A2(n549), .ZN(n550) );
  NAND2_X1 U653 ( .A1(n628), .A2(n550), .ZN(n551) );
  OR2_X1 U654 ( .A1(n568), .A2(n551), .ZN(n586) );
  AND2_X1 U655 ( .A1(n588), .A2(n586), .ZN(n558) );
  INV_X1 U656 ( .A(KEYINPUT113), .ZN(n552) );
  INV_X1 U657 ( .A(KEYINPUT85), .ZN(n555) );
  INV_X1 U658 ( .A(KEYINPUT35), .ZN(n556) );
  NAND2_X1 U659 ( .A1(n558), .A2(n671), .ZN(n560) );
  NOR2_X1 U660 ( .A1(KEYINPUT77), .A2(KEYINPUT44), .ZN(n559) );
  XNOR2_X1 U661 ( .A(n560), .B(n559), .ZN(n573) );
  OR2_X1 U662 ( .A1(n690), .A2(n351), .ZN(n712) );
  NAND2_X1 U663 ( .A1(n563), .A2(n712), .ZN(n564) );
  XNOR2_X1 U664 ( .A(n564), .B(KEYINPUT110), .ZN(n569) );
  NOR2_X1 U665 ( .A1(n698), .A2(n626), .ZN(n566) );
  NAND2_X1 U666 ( .A1(n566), .A2(n565), .ZN(n567) );
  OR2_X1 U667 ( .A1(n568), .A2(n567), .ZN(n587) );
  NAND2_X1 U668 ( .A1(KEYINPUT77), .A2(KEYINPUT44), .ZN(n570) );
  AND2_X1 U669 ( .A1(n571), .A2(n570), .ZN(n572) );
  INV_X1 U670 ( .A(KEYINPUT45), .ZN(n574) );
  NOR2_X1 U671 ( .A1(n643), .A2(G953), .ZN(n580) );
  XOR2_X1 U672 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n576) );
  NAND2_X1 U673 ( .A1(G224), .A2(G953), .ZN(n575) );
  XNOR2_X1 U674 ( .A(n576), .B(n575), .ZN(n578) );
  NOR2_X1 U675 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U676 ( .A1(n580), .A2(n579), .ZN(n585) );
  INV_X1 U677 ( .A(n581), .ZN(n583) );
  NAND2_X1 U678 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U679 ( .A(n585), .B(n584), .ZN(G69) );
  XNOR2_X1 U680 ( .A(n586), .B(G110), .ZN(G12) );
  XNOR2_X1 U681 ( .A(n587), .B(G101), .ZN(G3) );
  XNOR2_X1 U682 ( .A(n588), .B(G119), .ZN(G21) );
  INV_X1 U683 ( .A(n716), .ZN(n590) );
  NAND2_X1 U684 ( .A1(n593), .A2(n690), .ZN(n595) );
  XNOR2_X1 U685 ( .A(KEYINPUT115), .B(KEYINPUT40), .ZN(n594) );
  XOR2_X1 U686 ( .A(n617), .B(G131), .Z(G33) );
  AND2_X1 U687 ( .A1(n596), .A2(n700), .ZN(n605) );
  INV_X1 U688 ( .A(n605), .ZN(n597) );
  OR2_X1 U689 ( .A1(n701), .A2(n597), .ZN(n598) );
  XNOR2_X1 U690 ( .A(n599), .B(KEYINPUT28), .ZN(n601) );
  INV_X1 U691 ( .A(KEYINPUT71), .ZN(n602) );
  AND2_X1 U692 ( .A1(n712), .A2(n602), .ZN(n603) );
  XNOR2_X1 U693 ( .A(n604), .B(KEYINPUT47), .ZN(n616) );
  AND2_X1 U694 ( .A1(n631), .A2(n626), .ZN(n609) );
  NAND2_X1 U695 ( .A1(n605), .A2(n714), .ZN(n608) );
  NAND2_X1 U696 ( .A1(n606), .A2(n690), .ZN(n607) );
  NAND2_X1 U697 ( .A1(n609), .A2(n627), .ZN(n611) );
  INV_X1 U698 ( .A(KEYINPUT36), .ZN(n610) );
  XNOR2_X1 U699 ( .A(n611), .B(n610), .ZN(n612) );
  INV_X1 U700 ( .A(KEYINPUT116), .ZN(n620) );
  INV_X1 U701 ( .A(KEYINPUT46), .ZN(n623) );
  INV_X1 U702 ( .A(KEYINPUT48), .ZN(n625) );
  AND2_X1 U703 ( .A1(n627), .A2(n626), .ZN(n629) );
  NAND2_X1 U704 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U705 ( .A(n630), .B(KEYINPUT43), .ZN(n633) );
  INV_X1 U706 ( .A(n631), .ZN(n632) );
  NAND2_X1 U707 ( .A1(n633), .A2(n632), .ZN(n695) );
  NAND2_X1 U708 ( .A1(n634), .A2(n695), .ZN(n636) );
  INV_X1 U709 ( .A(KEYINPUT89), .ZN(n635) );
  XNOR2_X1 U710 ( .A(n636), .B(n635), .ZN(n646) );
  INV_X1 U711 ( .A(KEYINPUT68), .ZN(n640) );
  NAND2_X1 U712 ( .A1(n644), .A2(KEYINPUT2), .ZN(n639) );
  INV_X1 U713 ( .A(KEYINPUT2), .ZN(n642) );
  NAND2_X1 U714 ( .A1(n644), .A2(KEYINPUT68), .ZN(n645) );
  NOR2_X1 U715 ( .A1(n646), .A2(n752), .ZN(n647) );
  NAND2_X1 U716 ( .A1(n647), .A2(KEYINPUT2), .ZN(n648) );
  NAND2_X1 U717 ( .A1(n672), .A2(G472), .ZN(n652) );
  XOR2_X1 U718 ( .A(KEYINPUT92), .B(KEYINPUT62), .Z(n649) );
  XNOR2_X1 U719 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U720 ( .A(n652), .B(n651), .ZN(n653) );
  NAND2_X1 U721 ( .A1(n653), .A2(n676), .ZN(n654) );
  XNOR2_X1 U722 ( .A(n654), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U723 ( .A1(n672), .A2(G210), .ZN(n659) );
  XNOR2_X1 U724 ( .A(KEYINPUT123), .B(KEYINPUT54), .ZN(n655) );
  XOR2_X1 U725 ( .A(n655), .B(KEYINPUT55), .Z(n656) );
  XNOR2_X1 U726 ( .A(n659), .B(n658), .ZN(n660) );
  NAND2_X1 U727 ( .A1(n660), .A2(n676), .ZN(n662) );
  XOR2_X1 U728 ( .A(KEYINPUT90), .B(KEYINPUT56), .Z(n661) );
  XNOR2_X1 U729 ( .A(n662), .B(n661), .ZN(G51) );
  NAND2_X1 U730 ( .A1(n672), .A2(G475), .ZN(n667) );
  XNOR2_X1 U731 ( .A(KEYINPUT67), .B(KEYINPUT124), .ZN(n663) );
  XOR2_X1 U732 ( .A(n663), .B(KEYINPUT59), .Z(n664) );
  XNOR2_X1 U733 ( .A(n667), .B(n666), .ZN(n668) );
  NAND2_X1 U734 ( .A1(n668), .A2(n676), .ZN(n670) );
  XNOR2_X1 U735 ( .A(KEYINPUT69), .B(KEYINPUT60), .ZN(n669) );
  XNOR2_X1 U736 ( .A(n670), .B(n669), .ZN(G60) );
  XNOR2_X1 U737 ( .A(n671), .B(G122), .ZN(G24) );
  BUF_X2 U738 ( .A(n672), .Z(n738) );
  NAND2_X1 U739 ( .A1(n738), .A2(G478), .ZN(n675) );
  XNOR2_X1 U740 ( .A(n673), .B(KEYINPUT125), .ZN(n674) );
  XNOR2_X1 U741 ( .A(n675), .B(n674), .ZN(n677) );
  INV_X1 U742 ( .A(n676), .ZN(n742) );
  NOR2_X1 U743 ( .A1(n677), .A2(n742), .ZN(G63) );
  NAND2_X1 U744 ( .A1(n738), .A2(G469), .ZN(n681) );
  XOR2_X1 U745 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n678) );
  XNOR2_X1 U746 ( .A(n679), .B(n678), .ZN(n680) );
  XNOR2_X1 U747 ( .A(n681), .B(n680), .ZN(n682) );
  NOR2_X1 U748 ( .A1(n682), .A2(n742), .ZN(G54) );
  NAND2_X1 U749 ( .A1(n683), .A2(n351), .ZN(n685) );
  XOR2_X1 U750 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n684) );
  XNOR2_X1 U751 ( .A(n685), .B(n684), .ZN(n686) );
  XNOR2_X1 U752 ( .A(G107), .B(n686), .ZN(G9) );
  XOR2_X1 U753 ( .A(KEYINPUT118), .B(KEYINPUT29), .Z(n688) );
  NAND2_X1 U754 ( .A1(n342), .A2(n351), .ZN(n687) );
  XNOR2_X1 U755 ( .A(n688), .B(n687), .ZN(n689) );
  XNOR2_X1 U756 ( .A(G128), .B(n689), .ZN(G30) );
  XOR2_X1 U757 ( .A(G146), .B(KEYINPUT119), .Z(n692) );
  NAND2_X1 U758 ( .A1(n342), .A2(n690), .ZN(n691) );
  XNOR2_X1 U759 ( .A(n692), .B(n691), .ZN(G48) );
  XNOR2_X1 U760 ( .A(G125), .B(n693), .ZN(n694) );
  XNOR2_X1 U761 ( .A(n694), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U762 ( .A(n695), .B(G140), .ZN(n696) );
  XNOR2_X1 U763 ( .A(KEYINPUT120), .B(n696), .ZN(G42) );
  INV_X1 U764 ( .A(G953), .ZN(n736) );
  NOR2_X1 U765 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U766 ( .A(n699), .B(KEYINPUT50), .ZN(n706) );
  NOR2_X1 U767 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U768 ( .A(n702), .B(KEYINPUT49), .ZN(n704) );
  NAND2_X1 U769 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U770 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U771 ( .A(KEYINPUT121), .B(n707), .Z(n709) );
  NOR2_X1 U772 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U773 ( .A(n710), .B(KEYINPUT51), .ZN(n711) );
  NAND2_X1 U774 ( .A1(n711), .A2(n732), .ZN(n723) );
  NAND2_X1 U775 ( .A1(n712), .A2(n714), .ZN(n713) );
  OR2_X1 U776 ( .A1(n713), .A2(n716), .ZN(n720) );
  INV_X1 U777 ( .A(n714), .ZN(n715) );
  NAND2_X1 U778 ( .A1(n716), .A2(n715), .ZN(n718) );
  NAND2_X1 U779 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U780 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U781 ( .A1(n733), .A2(n721), .ZN(n722) );
  NAND2_X1 U782 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U783 ( .A(n724), .B(KEYINPUT52), .ZN(n725) );
  XOR2_X1 U784 ( .A(KEYINPUT122), .B(n725), .Z(n726) );
  NOR2_X1 U785 ( .A1(n727), .A2(n726), .ZN(n734) );
  XOR2_X1 U786 ( .A(KEYINPUT87), .B(n728), .Z(n730) );
  NOR2_X1 U787 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U788 ( .A1(n736), .A2(n735), .ZN(n737) );
  XOR2_X1 U789 ( .A(KEYINPUT53), .B(n737), .Z(G75) );
  NAND2_X1 U790 ( .A1(n738), .A2(G217), .ZN(n740) );
  XNOR2_X1 U791 ( .A(n740), .B(n739), .ZN(n741) );
  NOR2_X1 U792 ( .A1(n742), .A2(n741), .ZN(G66) );
  XNOR2_X1 U793 ( .A(n744), .B(n743), .ZN(n747) );
  XNOR2_X1 U794 ( .A(n745), .B(n747), .ZN(n746) );
  NAND2_X1 U795 ( .A1(n746), .A2(n527), .ZN(n751) );
  XNOR2_X1 U796 ( .A(n747), .B(G227), .ZN(n748) );
  NAND2_X1 U797 ( .A1(n748), .A2(G900), .ZN(n749) );
  NAND2_X1 U798 ( .A1(n749), .A2(G953), .ZN(n750) );
  NAND2_X1 U799 ( .A1(n751), .A2(n750), .ZN(G72) );
  XOR2_X1 U800 ( .A(G134), .B(n752), .Z(G36) );
endmodule

