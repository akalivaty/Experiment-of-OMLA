// Benchmark "locked_c1355" written by ABC on Sat Dec 16 10:33:30 2023

module locked_c1355 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat,
    G22gat, G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat,
    G85gat, G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat,
    G141gat, G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat,
    G197gat, G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat,
    G229gat, G230gat, G231gat, G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat,
    G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat, G57gat, G64gat,
    G71gat, G78gat, G85gat, G92gat, G99gat, G106gat, G113gat, G120gat,
    G127gat, G134gat, G141gat, G148gat, G155gat, G162gat, G169gat, G176gat,
    G183gat, G190gat, G197gat, G204gat, G211gat, G218gat, G225gat, G226gat,
    G227gat, G228gat, G229gat, G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n138, new_n139, new_n140, new_n141, new_n142, new_n143, new_n144,
    new_n145, new_n146, new_n147, new_n148, new_n149, new_n150, new_n151,
    new_n152, new_n153, new_n154, new_n155, new_n156, new_n157, new_n158,
    new_n159, new_n160, new_n161, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n503, new_n504,
    new_n506, new_n507, new_n508, new_n509, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n526, new_n527,
    new_n528, new_n529, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n557, new_n558, new_n560,
    new_n561, new_n562, new_n563, new_n565, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n631,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n675, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703;
  INV_X1    g000(.A(G190gat), .ZN(new_n138));
  AND2_X1   g001(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n139));
  NOR2_X1   g002(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n140));
  OAI21_X1  g003(.A(new_n138), .B1(new_n139), .B2(new_n140), .ZN(new_n141));
  NAND2_X1  g004(.A1(new_n141), .A2(KEYINPUT28), .ZN(new_n142));
  OR3_X1    g005(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n143));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n144));
  OAI21_X1  g007(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n145));
  NAND3_X1  g008(.A1(new_n143), .A2(new_n144), .A3(new_n145), .ZN(new_n146));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n147));
  INV_X1    g010(.A(KEYINPUT28), .ZN(new_n148));
  OAI211_X1 g011(.A(new_n148), .B(new_n138), .C1(new_n139), .C2(new_n140), .ZN(new_n149));
  NAND4_X1  g012(.A1(new_n142), .A2(new_n146), .A3(new_n147), .A4(new_n149), .ZN(new_n150));
  INV_X1    g013(.A(KEYINPUT24), .ZN(new_n151));
  NAND2_X1  g014(.A1(new_n147), .A2(new_n151), .ZN(new_n152));
  OR2_X1    g015(.A1(G183gat), .A2(G190gat), .ZN(new_n153));
  NAND3_X1  g016(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n154));
  NAND3_X1  g017(.A1(new_n152), .A2(new_n153), .A3(new_n154), .ZN(new_n155));
  INV_X1    g018(.A(KEYINPUT23), .ZN(new_n156));
  INV_X1    g019(.A(G169gat), .ZN(new_n157));
  INV_X1    g020(.A(G176gat), .ZN(new_n158));
  NAND3_X1  g021(.A1(new_n156), .A2(new_n157), .A3(new_n158), .ZN(new_n159));
  OAI21_X1  g022(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n160));
  NAND2_X1  g023(.A1(new_n159), .A2(new_n160), .ZN(new_n161));
  NAND3_X1  g024(.A1(new_n155), .A2(new_n161), .A3(new_n144), .ZN(new_n162));
  NAND2_X1  g025(.A1(new_n162), .A2(KEYINPUT25), .ZN(new_n163));
  INV_X1    g026(.A(KEYINPUT25), .ZN(new_n164));
  NAND4_X1  g027(.A1(new_n155), .A2(new_n161), .A3(new_n164), .A4(new_n144), .ZN(new_n165));
  NAND3_X1  g028(.A1(new_n150), .A2(new_n163), .A3(new_n165), .ZN(new_n166));
  AND2_X1   g029(.A1(G226gat), .A2(G233gat), .ZN(new_n167));
  OR2_X1    g030(.A1(new_n167), .A2(KEYINPUT29), .ZN(new_n168));
  NAND2_X1  g031(.A1(new_n166), .A2(new_n168), .ZN(new_n169));
  XNOR2_X1  g032(.A(G197gat), .B(G204gat), .ZN(new_n170));
  INV_X1    g033(.A(KEYINPUT22), .ZN(new_n171));
  INV_X1    g034(.A(G211gat), .ZN(new_n172));
  INV_X1    g035(.A(G218gat), .ZN(new_n173));
  OAI21_X1  g036(.A(new_n171), .B1(new_n172), .B2(new_n173), .ZN(new_n174));
  NAND2_X1  g037(.A1(new_n170), .A2(new_n174), .ZN(new_n175));
  XNOR2_X1  g038(.A(G211gat), .B(G218gat), .ZN(new_n176));
  XNOR2_X1  g039(.A(new_n175), .B(new_n176), .ZN(new_n177));
  INV_X1    g040(.A(new_n167), .ZN(new_n178));
  NAND4_X1  g041(.A1(new_n150), .A2(new_n163), .A3(new_n178), .A4(new_n165), .ZN(new_n179));
  AND3_X1   g042(.A1(new_n169), .A2(new_n177), .A3(new_n179), .ZN(new_n180));
  AOI21_X1  g043(.A(new_n177), .B1(new_n169), .B2(new_n179), .ZN(new_n181));
  OAI21_X1  g044(.A(KEYINPUT37), .B1(new_n180), .B2(new_n181), .ZN(new_n182));
  NAND2_X1  g045(.A1(new_n169), .A2(new_n179), .ZN(new_n183));
  INV_X1    g046(.A(new_n177), .ZN(new_n184));
  NAND2_X1  g047(.A1(new_n183), .A2(new_n184), .ZN(new_n185));
  INV_X1    g048(.A(KEYINPUT37), .ZN(new_n186));
  NAND3_X1  g049(.A1(new_n169), .A2(new_n177), .A3(new_n179), .ZN(new_n187));
  NAND3_X1  g050(.A1(new_n185), .A2(new_n186), .A3(new_n187), .ZN(new_n188));
  AND2_X1   g051(.A1(new_n182), .A2(new_n188), .ZN(new_n189));
  XOR2_X1   g052(.A(G8gat), .B(G36gat), .Z(new_n190));
  XNOR2_X1  g053(.A(new_n190), .B(G64gat), .ZN(new_n191));
  XOR2_X1   g054(.A(new_n191), .B(G92gat), .Z(new_n192));
  INV_X1    g055(.A(new_n192), .ZN(new_n193));
  OAI21_X1  g056(.A(KEYINPUT38), .B1(new_n189), .B2(new_n193), .ZN(new_n194));
  NAND2_X1  g057(.A1(G225gat), .A2(G233gat), .ZN(new_n195));
  INV_X1    g058(.A(G120gat), .ZN(new_n196));
  NAND2_X1  g059(.A1(new_n196), .A2(G113gat), .ZN(new_n197));
  INV_X1    g060(.A(G113gat), .ZN(new_n198));
  NAND2_X1  g061(.A1(new_n198), .A2(G120gat), .ZN(new_n199));
  NAND2_X1  g062(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g063(.A(KEYINPUT1), .ZN(new_n201));
  INV_X1    g064(.A(G134gat), .ZN(new_n202));
  NAND2_X1  g065(.A1(new_n202), .A2(G127gat), .ZN(new_n203));
  INV_X1    g066(.A(G127gat), .ZN(new_n204));
  NAND2_X1  g067(.A1(new_n204), .A2(G134gat), .ZN(new_n205));
  NAND4_X1  g068(.A1(new_n200), .A2(new_n201), .A3(new_n203), .A4(new_n205), .ZN(new_n206));
  NAND2_X1  g069(.A1(new_n203), .A2(new_n205), .ZN(new_n207));
  XNOR2_X1  g070(.A(G113gat), .B(G120gat), .ZN(new_n208));
  OAI21_X1  g071(.A(new_n207), .B1(new_n208), .B2(KEYINPUT1), .ZN(new_n209));
  NAND2_X1  g072(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  AND2_X1   g073(.A1(G155gat), .A2(G162gat), .ZN(new_n211));
  NOR2_X1   g074(.A1(G155gat), .A2(G162gat), .ZN(new_n212));
  NOR2_X1   g075(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OR2_X1    g076(.A1(G141gat), .A2(G148gat), .ZN(new_n214));
  NAND2_X1  g077(.A1(G141gat), .A2(G148gat), .ZN(new_n215));
  NAND2_X1  g078(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g079(.A(KEYINPUT2), .ZN(new_n217));
  AOI21_X1  g080(.A(new_n217), .B1(G155gat), .B2(G162gat), .ZN(new_n218));
  OAI21_X1  g081(.A(new_n213), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g082(.A(G155gat), .B(G162gat), .ZN(new_n220));
  INV_X1    g083(.A(G155gat), .ZN(new_n221));
  INV_X1    g084(.A(G162gat), .ZN(new_n222));
  OAI21_X1  g085(.A(KEYINPUT2), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND4_X1  g086(.A1(new_n220), .A2(new_n223), .A3(new_n214), .A4(new_n215), .ZN(new_n224));
  NAND2_X1  g087(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g088(.A1(new_n210), .A2(new_n225), .ZN(new_n226));
  NAND4_X1  g089(.A1(new_n219), .A2(new_n206), .A3(new_n209), .A4(new_n224), .ZN(new_n227));
  AOI21_X1  g090(.A(new_n195), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g091(.A1(new_n225), .A2(KEYINPUT3), .ZN(new_n229));
  INV_X1    g092(.A(KEYINPUT3), .ZN(new_n230));
  NAND3_X1  g093(.A1(new_n219), .A2(new_n224), .A3(new_n230), .ZN(new_n231));
  NAND3_X1  g094(.A1(new_n229), .A2(new_n210), .A3(new_n231), .ZN(new_n232));
  AND2_X1   g095(.A1(new_n206), .A2(new_n209), .ZN(new_n233));
  NAND4_X1  g096(.A1(new_n233), .A2(KEYINPUT4), .A3(new_n219), .A4(new_n224), .ZN(new_n234));
  INV_X1    g097(.A(KEYINPUT4), .ZN(new_n235));
  NAND2_X1  g098(.A1(new_n227), .A2(new_n235), .ZN(new_n236));
  NAND4_X1  g099(.A1(new_n232), .A2(new_n234), .A3(new_n195), .A4(new_n236), .ZN(new_n237));
  INV_X1    g100(.A(KEYINPUT5), .ZN(new_n238));
  AOI21_X1  g101(.A(new_n228), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  AND3_X1   g102(.A1(new_n219), .A2(new_n224), .A3(new_n230), .ZN(new_n240));
  AOI21_X1  g103(.A(new_n230), .B1(new_n219), .B2(new_n224), .ZN(new_n241));
  NOR2_X1   g104(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI22_X1  g105(.A1(new_n242), .A2(new_n210), .B1(new_n235), .B2(new_n227), .ZN(new_n243));
  NAND4_X1  g106(.A1(new_n243), .A2(KEYINPUT5), .A3(new_n195), .A4(new_n234), .ZN(new_n244));
  XNOR2_X1  g107(.A(G1gat), .B(G29gat), .ZN(new_n245));
  XNOR2_X1  g108(.A(new_n245), .B(KEYINPUT0), .ZN(new_n246));
  XNOR2_X1  g109(.A(new_n246), .B(G57gat), .ZN(new_n247));
  XNOR2_X1  g110(.A(new_n247), .B(G85gat), .ZN(new_n248));
  NAND3_X1  g111(.A1(new_n239), .A2(new_n244), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g112(.A1(new_n249), .A2(KEYINPUT6), .ZN(new_n250));
  NAND2_X1  g113(.A1(new_n239), .A2(new_n244), .ZN(new_n251));
  INV_X1    g114(.A(new_n248), .ZN(new_n252));
  NAND2_X1  g115(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g116(.A(KEYINPUT6), .ZN(new_n254));
  NAND4_X1  g117(.A1(new_n239), .A2(new_n244), .A3(new_n248), .A4(new_n254), .ZN(new_n255));
  NAND3_X1  g118(.A1(new_n250), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  OAI21_X1  g119(.A(new_n193), .B1(new_n180), .B2(new_n181), .ZN(new_n257));
  AOI21_X1  g120(.A(new_n193), .B1(new_n182), .B2(new_n188), .ZN(new_n258));
  INV_X1    g121(.A(KEYINPUT38), .ZN(new_n259));
  NAND2_X1  g122(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g123(.A1(new_n194), .A2(new_n256), .A3(new_n257), .A4(new_n260), .ZN(new_n261));
  NAND3_X1  g124(.A1(new_n232), .A2(new_n234), .A3(new_n236), .ZN(new_n262));
  INV_X1    g125(.A(new_n195), .ZN(new_n263));
  NAND2_X1  g126(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g127(.A(KEYINPUT39), .ZN(new_n265));
  NAND2_X1  g128(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g129(.A1(new_n226), .A2(new_n195), .A3(new_n227), .ZN(new_n267));
  NAND3_X1  g130(.A1(new_n262), .A2(KEYINPUT39), .A3(new_n263), .ZN(new_n268));
  NAND3_X1  g131(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g132(.A1(new_n269), .A2(new_n252), .ZN(new_n270));
  INV_X1    g133(.A(KEYINPUT40), .ZN(new_n271));
  NAND2_X1  g134(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g135(.A1(new_n269), .A2(KEYINPUT40), .A3(new_n252), .ZN(new_n273));
  INV_X1    g136(.A(KEYINPUT30), .ZN(new_n274));
  NAND2_X1  g137(.A1(new_n257), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g138(.A1(new_n185), .A2(new_n187), .A3(new_n192), .ZN(new_n276));
  OAI211_X1 g139(.A(KEYINPUT30), .B(new_n193), .C1(new_n180), .C2(new_n181), .ZN(new_n277));
  NAND3_X1  g140(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND4_X1  g141(.A1(new_n272), .A2(new_n249), .A3(new_n273), .A4(new_n278), .ZN(new_n279));
  XNOR2_X1  g142(.A(G22gat), .B(G50gat), .ZN(new_n280));
  NAND2_X1  g143(.A1(G228gat), .A2(G233gat), .ZN(new_n281));
  XNOR2_X1  g144(.A(new_n280), .B(new_n281), .ZN(new_n282));
  INV_X1    g145(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g146(.A(new_n230), .B1(new_n177), .B2(KEYINPUT29), .ZN(new_n284));
  NAND2_X1  g147(.A1(new_n284), .A2(new_n225), .ZN(new_n285));
  XNOR2_X1  g148(.A(G78gat), .B(G106gat), .ZN(new_n286));
  XNOR2_X1  g149(.A(new_n286), .B(KEYINPUT31), .ZN(new_n287));
  OAI21_X1  g150(.A(new_n177), .B1(new_n240), .B2(KEYINPUT29), .ZN(new_n288));
  NAND3_X1  g151(.A1(new_n285), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  INV_X1    g152(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g153(.A(new_n287), .B1(new_n285), .B2(new_n288), .ZN(new_n291));
  OAI21_X1  g154(.A(new_n283), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g155(.A(new_n291), .ZN(new_n293));
  NAND3_X1  g156(.A1(new_n293), .A2(new_n282), .A3(new_n289), .ZN(new_n294));
  NAND2_X1  g157(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g158(.A(new_n295), .ZN(new_n296));
  NAND3_X1  g159(.A1(new_n261), .A2(new_n279), .A3(new_n296), .ZN(new_n297));
  OAI21_X1  g160(.A(new_n295), .B1(new_n256), .B2(new_n278), .ZN(new_n298));
  INV_X1    g161(.A(KEYINPUT36), .ZN(new_n299));
  NAND2_X1  g162(.A1(new_n166), .A2(new_n210), .ZN(new_n300));
  NAND2_X1  g163(.A1(G227gat), .A2(G233gat), .ZN(new_n301));
  NAND4_X1  g164(.A1(new_n233), .A2(new_n150), .A3(new_n163), .A4(new_n165), .ZN(new_n302));
  NAND3_X1  g165(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g166(.A(KEYINPUT32), .ZN(new_n304));
  NAND2_X1  g167(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g168(.A1(new_n300), .A2(new_n302), .ZN(new_n306));
  INV_X1    g169(.A(new_n301), .ZN(new_n307));
  NAND2_X1  g170(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g171(.A1(new_n300), .A2(KEYINPUT32), .A3(new_n301), .A4(new_n302), .ZN(new_n309));
  AND3_X1   g172(.A1(new_n305), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  XNOR2_X1  g173(.A(G15gat), .B(G43gat), .ZN(new_n311));
  XNOR2_X1  g174(.A(new_n311), .B(G71gat), .ZN(new_n312));
  INV_X1    g175(.A(G99gat), .ZN(new_n313));
  XNOR2_X1  g176(.A(new_n312), .B(new_n313), .ZN(new_n314));
  AOI21_X1  g177(.A(new_n301), .B1(new_n300), .B2(new_n302), .ZN(new_n315));
  OAI21_X1  g178(.A(new_n314), .B1(new_n315), .B2(KEYINPUT33), .ZN(new_n316));
  NAND2_X1  g179(.A1(new_n316), .A2(KEYINPUT34), .ZN(new_n317));
  INV_X1    g180(.A(KEYINPUT34), .ZN(new_n318));
  OAI211_X1 g181(.A(new_n318), .B(new_n314), .C1(new_n315), .C2(KEYINPUT33), .ZN(new_n319));
  AND3_X1   g182(.A1(new_n310), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g183(.A(new_n310), .B1(new_n317), .B2(new_n319), .ZN(new_n321));
  OAI21_X1  g184(.A(new_n299), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g185(.A1(new_n317), .A2(new_n319), .ZN(new_n323));
  INV_X1    g186(.A(new_n310), .ZN(new_n324));
  NAND2_X1  g187(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g188(.A1(new_n310), .A2(new_n317), .A3(new_n319), .ZN(new_n326));
  NAND3_X1  g189(.A1(new_n325), .A2(KEYINPUT36), .A3(new_n326), .ZN(new_n327));
  AND3_X1   g190(.A1(new_n298), .A2(new_n322), .A3(new_n327), .ZN(new_n328));
  AND3_X1   g191(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n329));
  NAND4_X1  g192(.A1(new_n329), .A2(new_n253), .A3(new_n250), .A4(new_n255), .ZN(new_n330));
  OAI21_X1  g193(.A(new_n296), .B1(new_n320), .B2(new_n321), .ZN(new_n331));
  OAI21_X1  g194(.A(KEYINPUT35), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g195(.A(new_n295), .B1(new_n325), .B2(new_n326), .ZN(new_n333));
  NOR2_X1   g196(.A1(new_n256), .A2(new_n278), .ZN(new_n334));
  INV_X1    g197(.A(KEYINPUT35), .ZN(new_n335));
  NAND3_X1  g198(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  AOI22_X1  g199(.A1(new_n297), .A2(new_n328), .B1(new_n332), .B2(new_n336), .ZN(new_n337));
  INV_X1    g200(.A(KEYINPUT17), .ZN(new_n338));
  INV_X1    g201(.A(KEYINPUT14), .ZN(new_n339));
  INV_X1    g202(.A(G29gat), .ZN(new_n340));
  INV_X1    g203(.A(G36gat), .ZN(new_n341));
  NAND3_X1  g204(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  OAI21_X1  g205(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n343));
  AOI22_X1  g206(.A1(new_n342), .A2(new_n343), .B1(G29gat), .B2(G36gat), .ZN(new_n344));
  XNOR2_X1  g207(.A(G43gat), .B(G50gat), .ZN(new_n345));
  NAND2_X1  g208(.A1(new_n345), .A2(KEYINPUT15), .ZN(new_n346));
  INV_X1    g209(.A(G43gat), .ZN(new_n347));
  INV_X1    g210(.A(G50gat), .ZN(new_n348));
  NAND2_X1  g211(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g212(.A(KEYINPUT15), .ZN(new_n350));
  NAND2_X1  g213(.A1(G43gat), .A2(G50gat), .ZN(new_n351));
  NAND3_X1  g214(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  AND3_X1   g215(.A1(new_n344), .A2(new_n346), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g216(.A(new_n346), .B1(new_n352), .B2(new_n344), .ZN(new_n354));
  OAI21_X1  g217(.A(new_n338), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g218(.A1(new_n344), .A2(new_n352), .ZN(new_n356));
  INV_X1    g219(.A(new_n346), .ZN(new_n357));
  NAND2_X1  g220(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g221(.A1(new_n344), .A2(new_n346), .A3(new_n352), .ZN(new_n359));
  NAND3_X1  g222(.A1(new_n358), .A2(KEYINPUT17), .A3(new_n359), .ZN(new_n360));
  XNOR2_X1  g223(.A(G99gat), .B(G106gat), .ZN(new_n361));
  NAND2_X1  g224(.A1(G85gat), .A2(G92gat), .ZN(new_n362));
  NAND2_X1  g225(.A1(new_n362), .A2(KEYINPUT7), .ZN(new_n363));
  INV_X1    g226(.A(KEYINPUT7), .ZN(new_n364));
  NAND3_X1  g227(.A1(new_n364), .A2(G85gat), .A3(G92gat), .ZN(new_n365));
  NAND2_X1  g228(.A1(G99gat), .A2(G106gat), .ZN(new_n366));
  AOI22_X1  g229(.A1(new_n363), .A2(new_n365), .B1(KEYINPUT8), .B2(new_n366), .ZN(new_n367));
  OR2_X1    g230(.A1(G85gat), .A2(G92gat), .ZN(new_n368));
  AOI21_X1  g231(.A(new_n361), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g232(.A1(new_n363), .A2(new_n365), .ZN(new_n370));
  NAND2_X1  g233(.A1(new_n366), .A2(KEYINPUT8), .ZN(new_n371));
  NAND3_X1  g234(.A1(new_n370), .A2(new_n368), .A3(new_n371), .ZN(new_n372));
  INV_X1    g235(.A(new_n361), .ZN(new_n373));
  NOR2_X1   g236(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI211_X1 g237(.A(new_n355), .B(new_n360), .C1(new_n369), .C2(new_n374), .ZN(new_n375));
  NOR2_X1   g238(.A1(new_n374), .A2(new_n369), .ZN(new_n376));
  NAND2_X1  g239(.A1(new_n358), .A2(new_n359), .ZN(new_n377));
  AND2_X1   g240(.A1(G232gat), .A2(G233gat), .ZN(new_n378));
  AOI22_X1  g241(.A1(new_n376), .A2(new_n377), .B1(KEYINPUT41), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g242(.A(G134gat), .B(G162gat), .ZN(new_n380));
  XNOR2_X1  g243(.A(new_n380), .B(G190gat), .ZN(new_n381));
  AND3_X1   g244(.A1(new_n375), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g245(.A(new_n381), .B1(new_n375), .B2(new_n379), .ZN(new_n383));
  NOR2_X1   g246(.A1(new_n378), .A2(KEYINPUT41), .ZN(new_n384));
  XNOR2_X1  g247(.A(new_n384), .B(new_n173), .ZN(new_n385));
  OR3_X1    g248(.A1(new_n382), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  OAI21_X1  g249(.A(new_n385), .B1(new_n382), .B2(new_n383), .ZN(new_n387));
  NAND2_X1  g250(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g251(.A(new_n388), .ZN(new_n389));
  INV_X1    g252(.A(KEYINPUT12), .ZN(new_n390));
  XNOR2_X1  g253(.A(G113gat), .B(G141gat), .ZN(new_n391));
  INV_X1    g254(.A(KEYINPUT11), .ZN(new_n392));
  OR2_X1    g255(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g256(.A1(new_n391), .A2(new_n392), .ZN(new_n394));
  AOI21_X1  g257(.A(new_n157), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g258(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g259(.A1(new_n393), .A2(new_n157), .A3(new_n394), .ZN(new_n397));
  AOI21_X1  g260(.A(G197gat), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g261(.A(new_n397), .ZN(new_n399));
  INV_X1    g262(.A(G197gat), .ZN(new_n400));
  NOR3_X1   g263(.A1(new_n399), .A2(new_n400), .A3(new_n395), .ZN(new_n401));
  OAI21_X1  g264(.A(new_n390), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g265(.A(new_n400), .B1(new_n399), .B2(new_n395), .ZN(new_n403));
  NAND3_X1  g266(.A1(new_n396), .A2(G197gat), .A3(new_n397), .ZN(new_n404));
  NAND3_X1  g267(.A1(new_n403), .A2(new_n404), .A3(KEYINPUT12), .ZN(new_n405));
  NAND2_X1  g268(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g269(.A1(G229gat), .A2(G233gat), .ZN(new_n407));
  XNOR2_X1  g270(.A(new_n407), .B(KEYINPUT13), .ZN(new_n408));
  XNOR2_X1  g271(.A(G15gat), .B(G22gat), .ZN(new_n409));
  INV_X1    g272(.A(G1gat), .ZN(new_n410));
  NAND2_X1  g273(.A1(new_n410), .A2(KEYINPUT16), .ZN(new_n411));
  NAND2_X1  g274(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  INV_X1    g275(.A(G8gat), .ZN(new_n413));
  OAI211_X1 g276(.A(new_n412), .B(new_n413), .C1(G1gat), .C2(new_n409), .ZN(new_n414));
  INV_X1    g277(.A(G22gat), .ZN(new_n415));
  NAND2_X1  g278(.A1(new_n415), .A2(G15gat), .ZN(new_n416));
  INV_X1    g279(.A(G15gat), .ZN(new_n417));
  NAND2_X1  g280(.A1(new_n417), .A2(G22gat), .ZN(new_n418));
  AND3_X1   g281(.A1(new_n411), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g282(.A(G1gat), .B1(new_n416), .B2(new_n418), .ZN(new_n420));
  OAI21_X1  g283(.A(G8gat), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g284(.A1(new_n414), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g285(.A1(new_n377), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g286(.A1(new_n358), .A2(new_n359), .A3(new_n421), .A4(new_n414), .ZN(new_n424));
  AOI21_X1  g287(.A(new_n408), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AND2_X1   g288(.A1(new_n414), .A2(new_n421), .ZN(new_n426));
  NAND3_X1  g289(.A1(new_n355), .A2(new_n360), .A3(new_n426), .ZN(new_n427));
  NAND3_X1  g290(.A1(new_n427), .A2(new_n407), .A3(new_n423), .ZN(new_n428));
  INV_X1    g291(.A(KEYINPUT18), .ZN(new_n429));
  AOI21_X1  g292(.A(new_n425), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND4_X1  g293(.A1(new_n427), .A2(KEYINPUT18), .A3(new_n407), .A4(new_n423), .ZN(new_n431));
  AOI21_X1  g294(.A(new_n406), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g295(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g296(.A1(new_n430), .A2(new_n431), .A3(new_n406), .ZN(new_n434));
  NAND2_X1  g297(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g298(.A(new_n435), .ZN(new_n436));
  XOR2_X1   g299(.A(G57gat), .B(G64gat), .Z(new_n437));
  INV_X1    g300(.A(G71gat), .ZN(new_n438));
  INV_X1    g301(.A(G78gat), .ZN(new_n439));
  NAND2_X1  g302(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g303(.A1(G71gat), .A2(G78gat), .ZN(new_n441));
  NAND2_X1  g304(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g305(.A(KEYINPUT9), .ZN(new_n443));
  NAND2_X1  g306(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g307(.A1(new_n437), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  XNOR2_X1  g308(.A(G57gat), .B(G64gat), .ZN(new_n446));
  OAI211_X1 g309(.A(new_n441), .B(new_n440), .C1(new_n446), .C2(new_n443), .ZN(new_n447));
  NAND2_X1  g310(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  INV_X1    g311(.A(KEYINPUT21), .ZN(new_n449));
  NAND2_X1  g312(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g313(.A1(G231gat), .A2(G233gat), .ZN(new_n451));
  XOR2_X1   g314(.A(new_n450), .B(new_n451), .Z(new_n452));
  XNOR2_X1  g315(.A(G127gat), .B(G155gat), .ZN(new_n453));
  XNOR2_X1  g316(.A(new_n453), .B(KEYINPUT19), .ZN(new_n454));
  XNOR2_X1  g317(.A(new_n454), .B(KEYINPUT20), .ZN(new_n455));
  XNOR2_X1  g318(.A(new_n452), .B(new_n455), .ZN(new_n456));
  INV_X1    g319(.A(new_n448), .ZN(new_n457));
  AOI21_X1  g320(.A(new_n422), .B1(KEYINPUT21), .B2(new_n457), .ZN(new_n458));
  XOR2_X1   g321(.A(G183gat), .B(G211gat), .Z(new_n459));
  XNOR2_X1  g322(.A(new_n458), .B(new_n459), .ZN(new_n460));
  XNOR2_X1  g323(.A(new_n456), .B(new_n460), .ZN(new_n461));
  OAI21_X1  g324(.A(new_n448), .B1(new_n374), .B2(new_n369), .ZN(new_n462));
  INV_X1    g325(.A(KEYINPUT10), .ZN(new_n463));
  NAND2_X1  g326(.A1(new_n372), .A2(new_n373), .ZN(new_n464));
  NAND3_X1  g327(.A1(new_n367), .A2(new_n361), .A3(new_n368), .ZN(new_n465));
  NAND4_X1  g328(.A1(new_n464), .A2(new_n465), .A3(new_n447), .A4(new_n445), .ZN(new_n466));
  NAND3_X1  g329(.A1(new_n462), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g330(.A1(new_n376), .A2(KEYINPUT10), .A3(new_n457), .ZN(new_n468));
  NAND2_X1  g331(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g332(.A1(G230gat), .A2(G233gat), .ZN(new_n470));
  NAND2_X1  g333(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g334(.A1(new_n462), .A2(new_n466), .ZN(new_n472));
  INV_X1    g335(.A(new_n470), .ZN(new_n473));
  NAND2_X1  g336(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g337(.A(G120gat), .B(G148gat), .ZN(new_n475));
  XNOR2_X1  g338(.A(new_n475), .B(new_n158), .ZN(new_n476));
  INV_X1    g339(.A(G204gat), .ZN(new_n477));
  XNOR2_X1  g340(.A(new_n476), .B(new_n477), .ZN(new_n478));
  INV_X1    g341(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g342(.A1(new_n471), .A2(new_n474), .A3(new_n479), .ZN(new_n480));
  INV_X1    g343(.A(new_n474), .ZN(new_n481));
  AOI21_X1  g344(.A(new_n473), .B1(new_n467), .B2(new_n468), .ZN(new_n482));
  OAI21_X1  g345(.A(new_n478), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g346(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  INV_X1    g347(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g348(.A1(new_n461), .A2(new_n485), .ZN(new_n486));
  NOR4_X1   g349(.A1(new_n337), .A2(new_n389), .A3(new_n436), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g350(.A1(new_n487), .A2(new_n256), .ZN(new_n488));
  XNOR2_X1  g351(.A(new_n488), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g352(.A1(new_n487), .A2(new_n278), .ZN(new_n490));
  INV_X1    g353(.A(KEYINPUT42), .ZN(new_n491));
  XNOR2_X1  g354(.A(KEYINPUT16), .B(G8gat), .ZN(new_n492));
  OR3_X1    g355(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g356(.A1(new_n490), .A2(G8gat), .ZN(new_n494));
  OAI21_X1  g357(.A(new_n491), .B1(new_n490), .B2(new_n492), .ZN(new_n495));
  NAND3_X1  g358(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(G1325gat));
  NOR2_X1   g359(.A1(new_n320), .A2(new_n321), .ZN(new_n497));
  INV_X1    g360(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g361(.A1(new_n487), .A2(new_n417), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g362(.A1(new_n322), .A2(new_n327), .ZN(new_n500));
  AND2_X1   g363(.A1(new_n487), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g364(.A(new_n499), .B1(new_n501), .B2(new_n417), .ZN(G1326gat));
  NAND2_X1  g365(.A1(new_n487), .A2(new_n295), .ZN(new_n503));
  XNOR2_X1  g366(.A(KEYINPUT43), .B(G22gat), .ZN(new_n504));
  XNOR2_X1  g367(.A(new_n503), .B(new_n504), .ZN(G1327gat));
  OAI21_X1  g368(.A(KEYINPUT44), .B1(new_n337), .B2(new_n388), .ZN(new_n506));
  AND3_X1   g369(.A1(new_n261), .A2(new_n279), .A3(new_n296), .ZN(new_n507));
  NAND3_X1  g370(.A1(new_n298), .A2(new_n322), .A3(new_n327), .ZN(new_n508));
  AND3_X1   g371(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n509));
  AOI21_X1  g372(.A(new_n335), .B1(new_n333), .B2(new_n334), .ZN(new_n510));
  OAI22_X1  g373(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g374(.A(KEYINPUT44), .ZN(new_n512));
  NAND3_X1  g375(.A1(new_n511), .A2(new_n512), .A3(new_n389), .ZN(new_n513));
  NAND2_X1  g376(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g377(.A1(new_n436), .A2(new_n461), .ZN(new_n515));
  NAND3_X1  g378(.A1(new_n514), .A2(new_n485), .A3(new_n515), .ZN(new_n516));
  INV_X1    g379(.A(new_n256), .ZN(new_n517));
  OAI21_X1  g380(.A(G29gat), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g381(.A(new_n515), .ZN(new_n519));
  NOR3_X1   g382(.A1(new_n337), .A2(new_n388), .A3(new_n519), .ZN(new_n520));
  NAND4_X1  g383(.A1(new_n520), .A2(new_n340), .A3(new_n256), .A4(new_n485), .ZN(new_n521));
  INV_X1    g384(.A(KEYINPUT45), .ZN(new_n522));
  NAND2_X1  g385(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OR2_X1    g386(.A1(new_n521), .A2(new_n522), .ZN(new_n524));
  NAND3_X1  g387(.A1(new_n518), .A2(new_n523), .A3(new_n524), .ZN(G1328gat));
  OAI21_X1  g388(.A(G36gat), .B1(new_n516), .B2(new_n329), .ZN(new_n526));
  NAND4_X1  g389(.A1(new_n520), .A2(new_n341), .A3(new_n278), .A4(new_n485), .ZN(new_n527));
  NAND2_X1  g390(.A1(new_n527), .A2(KEYINPUT46), .ZN(new_n528));
  OR2_X1    g391(.A1(new_n527), .A2(KEYINPUT46), .ZN(new_n529));
  NAND3_X1  g392(.A1(new_n526), .A2(new_n528), .A3(new_n529), .ZN(G1329gat));
  INV_X1    g393(.A(KEYINPUT47), .ZN(new_n531));
  AOI211_X1 g394(.A(new_n484), .B(new_n519), .C1(new_n506), .C2(new_n513), .ZN(new_n532));
  AOI21_X1  g395(.A(new_n347), .B1(new_n532), .B2(new_n500), .ZN(new_n533));
  NOR2_X1   g396(.A1(new_n484), .A2(G43gat), .ZN(new_n534));
  NAND3_X1  g397(.A1(new_n520), .A2(new_n498), .A3(new_n534), .ZN(new_n535));
  INV_X1    g398(.A(new_n535), .ZN(new_n536));
  OAI21_X1  g399(.A(new_n531), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  INV_X1    g400(.A(new_n500), .ZN(new_n538));
  OAI21_X1  g401(.A(G43gat), .B1(new_n516), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g402(.A1(new_n539), .A2(KEYINPUT47), .A3(new_n535), .ZN(new_n540));
  NAND2_X1  g403(.A1(new_n537), .A2(new_n540), .ZN(G1330gat));
  INV_X1    g404(.A(KEYINPUT48), .ZN(new_n542));
  AOI21_X1  g405(.A(new_n348), .B1(new_n532), .B2(new_n295), .ZN(new_n543));
  NAND4_X1  g406(.A1(new_n520), .A2(new_n348), .A3(new_n295), .A4(new_n485), .ZN(new_n544));
  INV_X1    g407(.A(new_n544), .ZN(new_n545));
  OAI21_X1  g408(.A(new_n542), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g409(.A(G50gat), .B1(new_n516), .B2(new_n296), .ZN(new_n547));
  NAND3_X1  g410(.A1(new_n547), .A2(KEYINPUT48), .A3(new_n544), .ZN(new_n548));
  NAND2_X1  g411(.A1(new_n546), .A2(new_n548), .ZN(G1331gat));
  NOR2_X1   g412(.A1(new_n337), .A2(new_n435), .ZN(new_n550));
  INV_X1    g413(.A(new_n461), .ZN(new_n551));
  NOR3_X1   g414(.A1(new_n551), .A2(new_n389), .A3(new_n485), .ZN(new_n552));
  NAND2_X1  g415(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  INV_X1    g416(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g417(.A1(new_n554), .A2(new_n256), .ZN(new_n555));
  XNOR2_X1  g418(.A(new_n555), .B(G57gat), .ZN(G1332gat));
  AOI211_X1 g419(.A(new_n329), .B(new_n553), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n557));
  NOR2_X1   g420(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n558));
  XNOR2_X1  g421(.A(new_n557), .B(new_n558), .ZN(G1333gat));
  NAND3_X1  g422(.A1(new_n554), .A2(new_n438), .A3(new_n498), .ZN(new_n560));
  OAI21_X1  g423(.A(G71gat), .B1(new_n553), .B2(new_n538), .ZN(new_n561));
  NAND2_X1  g424(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g425(.A(KEYINPUT50), .ZN(new_n563));
  XNOR2_X1  g426(.A(new_n562), .B(new_n563), .ZN(G1334gat));
  NOR2_X1   g427(.A1(new_n553), .A2(new_n296), .ZN(new_n565));
  XNOR2_X1  g428(.A(new_n565), .B(new_n439), .ZN(G1335gat));
  NOR2_X1   g429(.A1(new_n461), .A2(new_n435), .ZN(new_n567));
  NAND3_X1  g430(.A1(new_n511), .A2(new_n389), .A3(new_n567), .ZN(new_n568));
  INV_X1    g431(.A(KEYINPUT51), .ZN(new_n569));
  NAND2_X1  g432(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g433(.A1(new_n511), .A2(KEYINPUT51), .A3(new_n389), .A4(new_n567), .ZN(new_n571));
  AOI21_X1  g434(.A(new_n485), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g435(.A(G85gat), .B1(new_n572), .B2(new_n256), .ZN(new_n573));
  NAND2_X1  g436(.A1(new_n567), .A2(new_n484), .ZN(new_n574));
  AOI21_X1  g437(.A(new_n574), .B1(new_n506), .B2(new_n513), .ZN(new_n575));
  AND2_X1   g438(.A1(new_n575), .A2(new_n256), .ZN(new_n576));
  AOI21_X1  g439(.A(new_n573), .B1(G85gat), .B2(new_n576), .ZN(G1336gat));
  INV_X1    g440(.A(KEYINPUT52), .ZN(new_n578));
  AOI21_X1  g441(.A(G92gat), .B1(new_n572), .B2(new_n278), .ZN(new_n579));
  NAND3_X1  g442(.A1(new_n575), .A2(G92gat), .A3(new_n278), .ZN(new_n580));
  INV_X1    g443(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g444(.A(new_n578), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  AOI211_X1 g445(.A(new_n329), .B(new_n485), .C1(new_n570), .C2(new_n571), .ZN(new_n583));
  OAI211_X1 g446(.A(KEYINPUT52), .B(new_n580), .C1(new_n583), .C2(G92gat), .ZN(new_n584));
  NAND2_X1  g447(.A1(new_n582), .A2(new_n584), .ZN(G1337gat));
  NAND3_X1  g448(.A1(new_n572), .A2(new_n313), .A3(new_n498), .ZN(new_n586));
  AND2_X1   g449(.A1(new_n575), .A2(new_n500), .ZN(new_n587));
  OAI21_X1  g450(.A(new_n586), .B1(new_n313), .B2(new_n587), .ZN(G1338gat));
  NAND2_X1  g451(.A1(new_n570), .A2(new_n571), .ZN(new_n589));
  NOR3_X1   g452(.A1(new_n296), .A2(G106gat), .A3(new_n485), .ZN(new_n590));
  NAND2_X1  g453(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g454(.A(new_n591), .ZN(new_n592));
  INV_X1    g455(.A(G106gat), .ZN(new_n593));
  AOI21_X1  g456(.A(new_n593), .B1(new_n575), .B2(new_n295), .ZN(new_n594));
  OAI21_X1  g457(.A(KEYINPUT53), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  INV_X1    g458(.A(KEYINPUT53), .ZN(new_n596));
  AND2_X1   g459(.A1(new_n575), .A2(new_n295), .ZN(new_n597));
  OAI211_X1 g460(.A(new_n591), .B(new_n596), .C1(new_n597), .C2(new_n593), .ZN(new_n598));
  NAND2_X1  g461(.A1(new_n595), .A2(new_n598), .ZN(G1339gat));
  NOR3_X1   g462(.A1(new_n486), .A2(new_n389), .A3(new_n435), .ZN(new_n600));
  AOI21_X1  g463(.A(KEYINPUT54), .B1(new_n469), .B2(new_n470), .ZN(new_n601));
  INV_X1    g464(.A(KEYINPUT54), .ZN(new_n602));
  AOI211_X1 g465(.A(new_n602), .B(new_n473), .C1(new_n467), .C2(new_n468), .ZN(new_n603));
  AND3_X1   g466(.A1(new_n467), .A2(new_n473), .A3(new_n468), .ZN(new_n604));
  NOR3_X1   g467(.A1(new_n601), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  OAI21_X1  g468(.A(KEYINPUT55), .B1(new_n605), .B2(new_n479), .ZN(new_n606));
  INV_X1    g469(.A(KEYINPUT55), .ZN(new_n607));
  NAND2_X1  g470(.A1(new_n471), .A2(new_n602), .ZN(new_n608));
  NAND2_X1  g471(.A1(new_n482), .A2(KEYINPUT54), .ZN(new_n609));
  NAND2_X1  g472(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI211_X1 g473(.A(new_n607), .B(new_n478), .C1(new_n610), .C2(new_n604), .ZN(new_n611));
  NAND2_X1  g474(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g475(.A(new_n407), .B1(new_n427), .B2(new_n423), .ZN(new_n613));
  AND3_X1   g476(.A1(new_n423), .A2(new_n424), .A3(new_n408), .ZN(new_n614));
  OAI211_X1 g477(.A(new_n404), .B(new_n403), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  AND3_X1   g478(.A1(new_n386), .A2(new_n387), .A3(new_n615), .ZN(new_n616));
  NAND4_X1  g479(.A1(new_n612), .A2(new_n434), .A3(new_n480), .A4(new_n616), .ZN(new_n617));
  AND3_X1   g480(.A1(new_n484), .A2(new_n434), .A3(new_n615), .ZN(new_n618));
  INV_X1    g481(.A(new_n480), .ZN(new_n619));
  AOI21_X1  g482(.A(new_n619), .B1(new_n433), .B2(new_n434), .ZN(new_n620));
  AOI21_X1  g483(.A(new_n618), .B1(new_n612), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g484(.A(new_n617), .B1(new_n621), .B2(new_n389), .ZN(new_n622));
  AOI21_X1  g485(.A(new_n600), .B1(new_n622), .B2(new_n551), .ZN(new_n623));
  NOR2_X1   g486(.A1(new_n623), .A2(new_n331), .ZN(new_n624));
  NOR2_X1   g487(.A1(new_n517), .A2(new_n278), .ZN(new_n625));
  NAND2_X1  g488(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g489(.A1(new_n626), .A2(new_n436), .ZN(new_n627));
  XNOR2_X1  g490(.A(new_n627), .B(new_n198), .ZN(G1340gat));
  NOR2_X1   g491(.A1(new_n626), .A2(new_n485), .ZN(new_n629));
  XNOR2_X1  g492(.A(new_n629), .B(new_n196), .ZN(G1341gat));
  NOR2_X1   g493(.A1(new_n626), .A2(new_n551), .ZN(new_n631));
  XNOR2_X1  g494(.A(new_n631), .B(new_n204), .ZN(G1342gat));
  AND2_X1   g495(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n633));
  NOR3_X1   g496(.A1(new_n626), .A2(new_n388), .A3(new_n633), .ZN(new_n634));
  NOR2_X1   g497(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n635));
  XNOR2_X1  g498(.A(new_n634), .B(new_n635), .ZN(G1343gat));
  NOR3_X1   g499(.A1(new_n623), .A2(new_n296), .A3(new_n500), .ZN(new_n637));
  NAND3_X1  g500(.A1(new_n637), .A2(new_n435), .A3(new_n625), .ZN(new_n638));
  INV_X1    g501(.A(G141gat), .ZN(new_n639));
  NAND2_X1  g502(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g503(.A(KEYINPUT57), .ZN(new_n641));
  OAI21_X1  g504(.A(new_n641), .B1(new_n623), .B2(new_n296), .ZN(new_n642));
  AND3_X1   g505(.A1(new_n430), .A2(new_n431), .A3(new_n406), .ZN(new_n643));
  OAI21_X1  g506(.A(new_n480), .B1(new_n643), .B2(new_n432), .ZN(new_n644));
  AOI21_X1  g507(.A(new_n644), .B1(new_n606), .B2(new_n611), .ZN(new_n645));
  OAI21_X1  g508(.A(new_n388), .B1(new_n645), .B2(new_n618), .ZN(new_n646));
  AOI21_X1  g509(.A(new_n461), .B1(new_n646), .B2(new_n617), .ZN(new_n647));
  OAI211_X1 g510(.A(KEYINPUT57), .B(new_n295), .C1(new_n647), .C2(new_n600), .ZN(new_n648));
  NAND2_X1  g511(.A1(new_n642), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g512(.A1(new_n649), .A2(new_n538), .A3(new_n435), .A4(new_n625), .ZN(new_n650));
  OAI21_X1  g513(.A(new_n640), .B1(new_n650), .B2(new_n639), .ZN(new_n651));
  INV_X1    g514(.A(KEYINPUT58), .ZN(new_n652));
  NAND2_X1  g515(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  OAI211_X1 g516(.A(KEYINPUT58), .B(new_n640), .C1(new_n650), .C2(new_n639), .ZN(new_n654));
  NAND2_X1  g517(.A1(new_n653), .A2(new_n654), .ZN(G1344gat));
  NOR2_X1   g518(.A1(new_n278), .A2(G148gat), .ZN(new_n656));
  NAND4_X1  g519(.A1(new_n637), .A2(new_n256), .A3(new_n484), .A4(new_n656), .ZN(new_n657));
  NAND4_X1  g520(.A1(new_n649), .A2(new_n538), .A3(new_n484), .A4(new_n625), .ZN(new_n658));
  INV_X1    g521(.A(KEYINPUT59), .ZN(new_n659));
  AND3_X1   g522(.A1(new_n658), .A2(new_n659), .A3(G148gat), .ZN(new_n660));
  AOI21_X1  g523(.A(new_n659), .B1(new_n658), .B2(G148gat), .ZN(new_n661));
  OAI21_X1  g524(.A(new_n657), .B1(new_n660), .B2(new_n661), .ZN(G1345gat));
  AND2_X1   g525(.A1(new_n637), .A2(new_n625), .ZN(new_n663));
  AOI21_X1  g526(.A(G155gat), .B1(new_n663), .B2(new_n461), .ZN(new_n664));
  AOI21_X1  g527(.A(new_n500), .B1(new_n642), .B2(new_n648), .ZN(new_n665));
  AND3_X1   g528(.A1(new_n665), .A2(new_n461), .A3(new_n625), .ZN(new_n666));
  AOI21_X1  g529(.A(new_n664), .B1(G155gat), .B2(new_n666), .ZN(G1346gat));
  NAND3_X1  g530(.A1(new_n663), .A2(new_n222), .A3(new_n389), .ZN(new_n668));
  AND3_X1   g531(.A1(new_n665), .A2(new_n389), .A3(new_n625), .ZN(new_n669));
  OAI21_X1  g532(.A(new_n668), .B1(new_n669), .B2(new_n222), .ZN(G1347gat));
  NOR2_X1   g533(.A1(new_n256), .A2(new_n329), .ZN(new_n671));
  NAND2_X1  g534(.A1(new_n624), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g535(.A1(new_n672), .A2(new_n436), .ZN(new_n673));
  XNOR2_X1  g536(.A(new_n673), .B(new_n157), .ZN(G1348gat));
  NOR2_X1   g537(.A1(new_n672), .A2(new_n485), .ZN(new_n675));
  XNOR2_X1  g538(.A(new_n675), .B(new_n158), .ZN(G1349gat));
  NAND3_X1  g539(.A1(new_n624), .A2(new_n461), .A3(new_n671), .ZN(new_n677));
  NAND2_X1  g540(.A1(new_n677), .A2(G183gat), .ZN(new_n678));
  NOR2_X1   g541(.A1(new_n139), .A2(new_n140), .ZN(new_n679));
  OAI21_X1  g542(.A(new_n678), .B1(new_n679), .B2(new_n677), .ZN(new_n680));
  XNOR2_X1  g543(.A(new_n680), .B(KEYINPUT60), .ZN(G1350gat));
  NOR2_X1   g544(.A1(new_n672), .A2(new_n388), .ZN(new_n682));
  INV_X1    g545(.A(KEYINPUT61), .ZN(new_n683));
  OAI21_X1  g546(.A(new_n682), .B1(new_n683), .B2(new_n138), .ZN(new_n684));
  XOR2_X1   g547(.A(KEYINPUT61), .B(G190gat), .Z(new_n685));
  OAI21_X1  g548(.A(new_n684), .B1(new_n682), .B2(new_n685), .ZN(G1351gat));
  AND2_X1   g549(.A1(new_n637), .A2(new_n671), .ZN(new_n687));
  NAND3_X1  g550(.A1(new_n687), .A2(new_n400), .A3(new_n435), .ZN(new_n688));
  AND3_X1   g551(.A1(new_n665), .A2(new_n435), .A3(new_n671), .ZN(new_n689));
  OAI21_X1  g552(.A(new_n688), .B1(new_n689), .B2(new_n400), .ZN(G1352gat));
  NAND3_X1  g553(.A1(new_n687), .A2(new_n477), .A3(new_n484), .ZN(new_n691));
  NAND2_X1  g554(.A1(new_n691), .A2(KEYINPUT62), .ZN(new_n692));
  INV_X1    g555(.A(KEYINPUT62), .ZN(new_n693));
  NAND4_X1  g556(.A1(new_n687), .A2(new_n693), .A3(new_n477), .A4(new_n484), .ZN(new_n694));
  AND3_X1   g557(.A1(new_n665), .A2(new_n484), .A3(new_n671), .ZN(new_n695));
  OAI211_X1 g558(.A(new_n692), .B(new_n694), .C1(new_n477), .C2(new_n695), .ZN(G1353gat));
  NAND3_X1  g559(.A1(new_n687), .A2(new_n172), .A3(new_n461), .ZN(new_n697));
  NAND4_X1  g560(.A1(new_n649), .A2(new_n538), .A3(new_n461), .A4(new_n671), .ZN(new_n698));
  AND3_X1   g561(.A1(new_n698), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n699));
  AOI21_X1  g562(.A(KEYINPUT63), .B1(new_n698), .B2(G211gat), .ZN(new_n700));
  OAI21_X1  g563(.A(new_n697), .B1(new_n699), .B2(new_n700), .ZN(G1354gat));
  NAND3_X1  g564(.A1(new_n687), .A2(new_n173), .A3(new_n389), .ZN(new_n702));
  AND3_X1   g565(.A1(new_n665), .A2(new_n389), .A3(new_n671), .ZN(new_n703));
  OAI21_X1  g566(.A(new_n702), .B1(new_n703), .B2(new_n173), .ZN(G1355gat));
endmodule


