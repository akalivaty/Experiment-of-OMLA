//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n555, new_n557, new_n558, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n572, new_n573, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  NAND2_X1  g033(.A1(G113), .A2(G2104), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G125), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  OR2_X1    g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n469), .A2(G137), .B1(G101), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n466), .A2(new_n473), .ZN(G160));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  OAI21_X1  g050(.A(KEYINPUT66), .B1(new_n462), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n467), .A2(new_n468), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT66), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n477), .A2(new_n478), .A3(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n480), .A2(KEYINPUT67), .A3(G124), .ZN(new_n484));
  AOI22_X1  g059(.A1(new_n483), .A2(new_n484), .B1(G136), .B2(new_n469), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NAND2_X1  g064(.A1(G114), .A2(G2104), .ZN(new_n490));
  INV_X1    g065(.A(G126), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n462), .B2(new_n491), .ZN(new_n492));
  AOI22_X1  g067(.A1(new_n492), .A2(G2105), .B1(G102), .B2(new_n471), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n469), .A2(new_n494), .A3(G138), .ZN(new_n495));
  OAI211_X1 g070(.A(G138), .B(new_n475), .C1(new_n460), .C2(new_n461), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n501), .B1(new_n502), .B2(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(KEYINPUT70), .A3(G543), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n503), .A2(new_n505), .B1(KEYINPUT5), .B2(new_n502), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n510), .B1(new_n508), .B2(KEYINPUT68), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT68), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(KEYINPUT6), .A3(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n506), .A2(new_n514), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n514), .A2(G50), .A3(G543), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT69), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n517), .B(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n516), .A2(new_n519), .ZN(G166));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n514), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n503), .A2(new_n505), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n502), .A2(KEYINPUT5), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n514), .A2(KEYINPUT71), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT71), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n511), .A2(new_n528), .A3(new_n513), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n527), .A2(G543), .A3(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G51), .ZN(new_n531));
  OAI221_X1 g106(.A(new_n522), .B1(new_n523), .B2(new_n526), .C1(new_n530), .C2(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  AND3_X1   g108(.A1(new_n527), .A2(G543), .A3(new_n529), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n534), .A2(G52), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n536), .A2(new_n508), .B1(new_n537), .B2(new_n515), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n535), .A2(new_n538), .ZN(G301));
  INV_X1    g114(.A(G301), .ZN(G171));
  XOR2_X1   g115(.A(KEYINPUT72), .B(G43), .Z(new_n541));
  NAND4_X1  g116(.A1(new_n527), .A2(G543), .A3(new_n529), .A4(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n506), .A2(G81), .A3(new_n514), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  OAI211_X1 g119(.A(new_n542), .B(new_n543), .C1(new_n544), .C2(new_n508), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(KEYINPUT73), .ZN(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n526), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT73), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n550), .A2(new_n551), .A3(new_n543), .A4(new_n542), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n546), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  AND3_X1   g129(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G36), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n558), .ZN(G188));
  AOI22_X1  g134(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT74), .B1(new_n560), .B2(new_n508), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n524), .A2(G65), .A3(new_n525), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT74), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n564), .A2(new_n565), .A3(G651), .ZN(new_n566));
  INV_X1    g141(.A(new_n515), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n561), .A2(new_n566), .B1(G91), .B2(new_n567), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n527), .A2(G53), .A3(G543), .A4(new_n529), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT9), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(G299));
  INV_X1    g146(.A(new_n516), .ZN(new_n572));
  INV_X1    g147(.A(new_n519), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(G303));
  INV_X1    g149(.A(KEYINPUT75), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n534), .A2(new_n575), .A3(G49), .ZN(new_n576));
  INV_X1    g151(.A(G49), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT75), .B1(new_n530), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n576), .A2(new_n578), .B1(G87), .B2(new_n567), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(G288));
  NAND3_X1  g156(.A1(new_n506), .A2(G86), .A3(new_n514), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n514), .A2(G48), .A3(G543), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n506), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n584));
  OAI211_X1 g159(.A(new_n582), .B(new_n583), .C1(new_n584), .C2(new_n508), .ZN(G305));
  NAND4_X1  g160(.A1(new_n527), .A2(G47), .A3(G543), .A4(new_n529), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n506), .A2(G85), .A3(new_n514), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  OAI211_X1 g163(.A(new_n586), .B(new_n587), .C1(new_n588), .C2(new_n508), .ZN(new_n589));
  AND2_X1   g164(.A1(new_n589), .A2(KEYINPUT76), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n589), .A2(KEYINPUT76), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G290));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  INV_X1    g169(.A(G92), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n515), .B2(new_n595), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n506), .A2(KEYINPUT10), .A3(G92), .A4(new_n514), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n506), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n599), .A2(new_n508), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n534), .A2(G54), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n598), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(G171), .B2(new_n603), .ZN(G284));
  OAI21_X1  g180(.A(new_n604), .B1(G171), .B2(new_n603), .ZN(G321));
  NAND2_X1  g181(.A1(G286), .A2(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n567), .A2(G91), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n565), .B1(new_n564), .B2(G651), .ZN(new_n609));
  AOI211_X1 g184(.A(KEYINPUT74), .B(new_n508), .C1(new_n562), .C2(new_n563), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT9), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n569), .B(new_n612), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n607), .B1(new_n614), .B2(G868), .ZN(G297));
  XNOR2_X1  g190(.A(G297), .B(KEYINPUT77), .ZN(G280));
  INV_X1    g191(.A(new_n602), .ZN(new_n617));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G860), .ZN(G148));
  NOR2_X1   g194(.A1(new_n602), .A2(G559), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n553), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n477), .A2(new_n471), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT12), .Z(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT13), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2100), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n475), .A2(G111), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n470), .B1(new_n629), .B2(KEYINPUT78), .ZN(new_n630));
  OAI221_X1 g205(.A(new_n630), .B1(KEYINPUT78), .B2(new_n629), .C1(G99), .C2(G2105), .ZN(new_n631));
  INV_X1    g206(.A(G135), .ZN(new_n632));
  INV_X1    g207(.A(new_n469), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n634), .B1(G123), .B2(new_n480), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2096), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n628), .A2(new_n636), .ZN(G156));
  XOR2_X1   g212(.A(G1341), .B(G1348), .Z(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2451), .B(G2454), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT80), .Z(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2427), .B(G2430), .Z(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n645), .A2(KEYINPUT79), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(KEYINPUT79), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(G2438), .A3(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  AOI21_X1  g224(.A(G2438), .B1(new_n646), .B2(new_n647), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n644), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n652), .A2(new_n643), .A3(new_n648), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n651), .A2(new_n653), .A3(KEYINPUT14), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n654), .A2(G2443), .ZN(new_n655));
  INV_X1    g230(.A(G2443), .ZN(new_n656));
  NAND4_X1  g231(.A1(new_n651), .A2(new_n653), .A3(KEYINPUT14), .A4(new_n656), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n642), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT16), .B(G2446), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n655), .A2(new_n657), .A3(new_n642), .ZN(new_n661));
  AND3_X1   g236(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n660), .B1(new_n659), .B2(new_n661), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n639), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT81), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n662), .A2(new_n663), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(new_n638), .ZN(new_n668));
  OAI211_X1 g243(.A(KEYINPUT81), .B(new_n639), .C1(new_n662), .C2(new_n663), .ZN(new_n669));
  NAND4_X1  g244(.A1(new_n666), .A2(new_n668), .A3(G14), .A4(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G401));
  XNOR2_X1  g246(.A(G2084), .B(G2090), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2072), .B(G2078), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT82), .ZN(new_n676));
  INV_X1    g251(.A(new_n673), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n674), .B(KEYINPUT17), .Z(new_n678));
  OAI21_X1  g253(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n672), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n678), .A2(new_n677), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n680), .A2(new_n673), .A3(new_n674), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT18), .Z(new_n683));
  NAND3_X1  g258(.A1(new_n679), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT83), .ZN(new_n685));
  XNOR2_X1  g260(.A(G2096), .B(G2100), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G227));
  XOR2_X1   g262(.A(G1956), .B(G2474), .Z(new_n688));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1971), .B(G1976), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT19), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n688), .A2(new_n689), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n697));
  AOI21_X1  g272(.A(new_n694), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n691), .A2(new_n693), .A3(new_n695), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n698), .B(new_n699), .C1(new_n696), .C2(new_n697), .ZN(new_n700));
  XOR2_X1   g275(.A(G1991), .B(G1996), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(G1981), .B(G1986), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT85), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n704), .B(new_n706), .Z(G229));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G26), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n469), .A2(G140), .ZN(new_n710));
  NOR2_X1   g285(.A1(G104), .A2(G2105), .ZN(new_n711));
  OAI21_X1  g286(.A(G2104), .B1(new_n475), .B2(G116), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(G128), .B2(new_n480), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n714), .A2(new_n708), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(new_n709), .ZN(new_n716));
  MUX2_X1   g291(.A(new_n709), .B(new_n716), .S(KEYINPUT28), .Z(new_n717));
  NOR2_X1   g292(.A1(new_n717), .A2(G2067), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n708), .A2(G35), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G162), .B2(new_n708), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT29), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G2090), .ZN(new_n722));
  INV_X1    g297(.A(G1961), .ZN(new_n723));
  NAND2_X1  g298(.A1(G171), .A2(G16), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G5), .B2(G16), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n722), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G16), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G21), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G168), .B2(new_n727), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT92), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G1966), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT93), .Z(new_n733));
  NAND2_X1  g308(.A1(new_n708), .A2(G32), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n480), .A2(G129), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n469), .A2(G141), .B1(G105), .B2(new_n471), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT26), .Z(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n734), .B1(new_n741), .B2(new_n708), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT91), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT27), .B(G1996), .Z(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NOR3_X1   g320(.A1(new_n726), .A2(new_n733), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n727), .A2(G20), .ZN(new_n747));
  OAI211_X1 g322(.A(KEYINPUT23), .B(new_n747), .C1(new_n614), .C2(new_n727), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(KEYINPUT23), .B2(new_n747), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT95), .B(G1956), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n721), .A2(G2090), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n727), .A2(KEYINPUT88), .A3(G19), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n553), .B2(new_n727), .ZN(new_n754));
  AOI21_X1  g329(.A(KEYINPUT88), .B1(new_n727), .B2(G19), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT89), .B(G1341), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n752), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n731), .A2(G1966), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT94), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n469), .A2(G139), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT90), .Z(new_n763));
  NAND2_X1  g338(.A1(new_n471), .A2(G103), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT25), .Z(new_n765));
  AOI22_X1  g340(.A1(new_n477), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n763), .B(new_n765), .C1(new_n475), .C2(new_n766), .ZN(new_n767));
  MUX2_X1   g342(.A(G33), .B(new_n767), .S(G29), .Z(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(G2072), .Z(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT31), .B(G11), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n708), .A2(G27), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G164), .B2(new_n708), .ZN(new_n772));
  INV_X1    g347(.A(G2078), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  OR2_X1    g349(.A1(KEYINPUT30), .A2(G28), .ZN(new_n775));
  NAND2_X1  g350(.A1(KEYINPUT30), .A2(G28), .ZN(new_n776));
  AOI21_X1  g351(.A(G29), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n635), .B2(G29), .ZN(new_n778));
  AND2_X1   g353(.A1(KEYINPUT24), .A2(G34), .ZN(new_n779));
  NOR2_X1   g354(.A1(KEYINPUT24), .A2(G34), .ZN(new_n780));
  NOR3_X1   g355(.A1(new_n779), .A2(new_n780), .A3(G29), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G160), .B2(new_n708), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n783), .A2(G2084), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(G2084), .ZN(new_n785));
  AND3_X1   g360(.A1(new_n778), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n769), .A2(new_n770), .A3(new_n774), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n717), .A2(G2067), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n727), .A2(G4), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n617), .B2(new_n727), .ZN(new_n790));
  INV_X1    g365(.A(G1348), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n725), .A2(new_n723), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n788), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NOR3_X1   g369(.A1(new_n761), .A2(new_n787), .A3(new_n794), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n746), .A2(new_n751), .A3(new_n759), .A4(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(G1976), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n727), .B1(new_n579), .B2(new_n580), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n727), .A2(G23), .ZN(new_n799));
  OAI21_X1  g374(.A(KEYINPUT33), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n798), .A2(KEYINPUT33), .A3(new_n799), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n797), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n727), .A2(G22), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G166), .B2(new_n727), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n805), .A2(G1971), .ZN(new_n806));
  OR3_X1    g381(.A1(new_n798), .A2(KEYINPUT33), .A3(new_n799), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n807), .A2(G1976), .A3(new_n800), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n805), .A2(G1971), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n803), .A2(new_n806), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  MUX2_X1   g385(.A(G6), .B(G305), .S(G16), .Z(new_n811));
  XOR2_X1   g386(.A(KEYINPUT86), .B(KEYINPUT32), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1981), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n811), .B(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(KEYINPUT34), .B1(new_n810), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(KEYINPUT87), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT87), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n817), .B(KEYINPUT34), .C1(new_n810), .C2(new_n814), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n592), .A2(new_n727), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(new_n727), .B2(G24), .ZN(new_n821));
  INV_X1    g396(.A(G1986), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n810), .A2(KEYINPUT34), .A3(new_n814), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n708), .A2(G25), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n480), .A2(G119), .ZN(new_n826));
  OR2_X1    g401(.A1(G95), .A2(G2105), .ZN(new_n827));
  INV_X1    g402(.A(G107), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n470), .B1(new_n828), .B2(G2105), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n469), .A2(G131), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n825), .B1(new_n831), .B2(new_n708), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT35), .B(G1991), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n832), .B(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n821), .B2(new_n822), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n824), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n819), .A2(new_n823), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT36), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT36), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n819), .A2(new_n840), .A3(new_n823), .A4(new_n837), .ZN(new_n841));
  AOI211_X1 g416(.A(new_n718), .B(new_n796), .C1(new_n839), .C2(new_n841), .ZN(G311));
  NAND2_X1  g417(.A1(new_n839), .A2(new_n841), .ZN(new_n843));
  INV_X1    g418(.A(new_n718), .ZN(new_n844));
  INV_X1    g419(.A(new_n796), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(G150));
  AND3_X1   g421(.A1(new_n504), .A2(KEYINPUT70), .A3(G543), .ZN(new_n847));
  AOI21_X1  g422(.A(KEYINPUT70), .B1(new_n504), .B2(G543), .ZN(new_n848));
  OAI211_X1 g423(.A(G67), .B(new_n525), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(G80), .A2(G543), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT96), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n849), .A2(KEYINPUT96), .A3(new_n850), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n853), .A2(G651), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(KEYINPUT97), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n534), .A2(G55), .B1(new_n567), .B2(G93), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT97), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n853), .A2(new_n858), .A3(new_n854), .A4(G651), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n856), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(G860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT37), .Z(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n553), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT98), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n856), .A2(new_n545), .A3(new_n857), .A4(new_n859), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n864), .B1(new_n863), .B2(new_n865), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n617), .A2(G559), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(KEYINPUT39), .Z(new_n871));
  OR2_X1    g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n869), .A2(new_n871), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n874), .B(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n878));
  INV_X1    g453(.A(G860), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n878), .B1(new_n877), .B2(new_n879), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n862), .B1(new_n880), .B2(new_n881), .ZN(G145));
  INV_X1    g457(.A(G37), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n480), .A2(G130), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT102), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n469), .A2(G142), .ZN(new_n886));
  NOR2_X1   g461(.A1(G106), .A2(G2105), .ZN(new_n887));
  OAI21_X1  g462(.A(G2104), .B1(new_n475), .B2(G118), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n885), .B(new_n886), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n889), .A2(new_n626), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(new_n626), .ZN(new_n891));
  INV_X1    g466(.A(new_n831), .ZN(new_n892));
  OR3_X1    g467(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n892), .B1(new_n890), .B2(new_n891), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n893), .A2(KEYINPUT103), .A3(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n714), .B(new_n499), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(new_n740), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT101), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(new_n898), .A3(new_n767), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n896), .B(new_n741), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n767), .B(KEYINPUT101), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n895), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(G160), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n488), .B(new_n905), .ZN(new_n906));
  XOR2_X1   g481(.A(new_n906), .B(new_n635), .Z(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n893), .A2(new_n894), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT103), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n910), .A2(new_n903), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n883), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n910), .A2(new_n903), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n910), .A2(new_n903), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n908), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT104), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n914), .A2(KEYINPUT103), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n907), .B1(new_n903), .B2(new_n895), .ZN(new_n920));
  AOI21_X1  g495(.A(G37), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n922));
  INV_X1    g497(.A(new_n916), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n907), .B1(new_n923), .B2(new_n914), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n921), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n918), .A2(new_n925), .A3(KEYINPUT40), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT40), .B1(new_n918), .B2(new_n925), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(G395));
  NAND2_X1  g503(.A1(new_n860), .A2(new_n603), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n869), .A2(new_n620), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n863), .A2(new_n865), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(KEYINPUT98), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n866), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n621), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n602), .A2(new_n568), .A3(new_n570), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n602), .B1(new_n568), .B2(new_n570), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT41), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n940), .B1(new_n936), .B2(new_n937), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT105), .ZN(new_n942));
  XOR2_X1   g517(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n943));
  NAND2_X1  g518(.A1(new_n938), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT105), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n945), .B(new_n940), .C1(new_n936), .C2(new_n937), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n942), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n939), .B1(new_n935), .B2(new_n947), .ZN(new_n948));
  XOR2_X1   g523(.A(G305), .B(KEYINPUT107), .Z(new_n949));
  NAND2_X1  g524(.A1(new_n589), .A2(KEYINPUT76), .ZN(new_n950));
  NAND2_X1  g525(.A1(G72), .A2(G543), .ZN(new_n951));
  INV_X1    g526(.A(G60), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n951), .B1(new_n526), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(G651), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT76), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n954), .A2(new_n955), .A3(new_n586), .A4(new_n587), .ZN(new_n956));
  AND3_X1   g531(.A1(G166), .A2(new_n950), .A3(new_n956), .ZN(new_n957));
  AOI22_X1  g532(.A1(new_n950), .A2(new_n956), .B1(new_n572), .B2(new_n573), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n949), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(G303), .B1(new_n590), .B2(new_n591), .ZN(new_n960));
  XNOR2_X1  g535(.A(G305), .B(KEYINPUT107), .ZN(new_n961));
  NAND3_X1  g536(.A1(G166), .A2(new_n950), .A3(new_n956), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n959), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(G288), .ZN(new_n965));
  INV_X1    g540(.A(G288), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n959), .A2(new_n963), .A3(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n965), .A2(KEYINPUT108), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT108), .B1(new_n965), .B2(new_n967), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT42), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n970), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT42), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(new_n973), .A3(new_n968), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  XOR2_X1   g550(.A(new_n948), .B(new_n975), .Z(new_n976));
  OAI21_X1  g551(.A(new_n929), .B1(new_n976), .B2(new_n603), .ZN(G295));
  OAI21_X1  g552(.A(new_n929), .B1(new_n976), .B2(new_n603), .ZN(G331));
  INV_X1    g553(.A(KEYINPUT43), .ZN(new_n979));
  INV_X1    g554(.A(new_n938), .ZN(new_n980));
  XNOR2_X1  g555(.A(G301), .B(G286), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n867), .A2(new_n868), .A3(new_n981), .ZN(new_n982));
  XNOR2_X1  g557(.A(G301), .B(G168), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n983), .B1(new_n932), .B2(new_n866), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n980), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n965), .A2(new_n967), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n981), .B1(new_n867), .B2(new_n868), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n932), .A2(new_n866), .A3(new_n983), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n947), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n985), .A2(new_n986), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n883), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT109), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n959), .A2(new_n963), .A3(new_n966), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n966), .B1(new_n959), .B2(new_n963), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n965), .A2(KEYINPUT109), .A3(new_n967), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n943), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n614), .A2(new_n602), .ZN(new_n999));
  NAND2_X1  g574(.A1(G299), .A2(new_n617), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1001), .B1(new_n940), .B2(new_n938), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n987), .A2(new_n988), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n997), .B1(new_n985), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT110), .B1(new_n991), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n985), .A2(new_n1003), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n995), .A2(new_n996), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT110), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1008), .A2(new_n1009), .A3(new_n883), .A4(new_n990), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n979), .B1(new_n1005), .B2(new_n1010), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n990), .A2(new_n883), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n985), .A2(new_n989), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n1007), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT43), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT44), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT44), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n979), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n991), .A2(new_n1004), .A3(KEYINPUT43), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1016), .A2(new_n1020), .ZN(G397));
  NAND3_X1  g596(.A1(new_n465), .A2(G40), .A3(new_n472), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT111), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT111), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n465), .A2(new_n1024), .A3(new_n472), .A4(G40), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT45), .ZN(new_n1027));
  INV_X1    g602(.A(G1384), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n499), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1026), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G1996), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n741), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G2067), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n714), .B(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n740), .A2(G1996), .ZN(new_n1036));
  OR3_X1    g611(.A1(new_n1033), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1037), .B1(new_n833), .B2(new_n892), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n831), .A2(new_n834), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n592), .A2(new_n822), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n592), .A2(new_n822), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1031), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n1045));
  OR3_X1    g620(.A1(G305), .A2(new_n1045), .A3(G1981), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1045), .B1(G305), .B2(G1981), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g623(.A(KEYINPUT117), .B(G86), .ZN(new_n1049));
  OAI221_X1 g624(.A(new_n583), .B1(new_n515), .B2(new_n1049), .C1(new_n584), .C2(new_n508), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(G1981), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT49), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1029), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1055));
  INV_X1    g630(.A(G8), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1048), .A2(KEYINPUT49), .A3(new_n1051), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1054), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(KEYINPUT113), .B1(G288), .B2(new_n797), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT113), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n579), .A2(new_n1062), .A3(G1976), .A4(new_n580), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1061), .A2(new_n1057), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT52), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT114), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT114), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1064), .A2(new_n1067), .A3(KEYINPUT52), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1060), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT50), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1029), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(G1384), .B1(new_n493), .B2(new_n498), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT50), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n1071), .A2(new_n1073), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1074));
  XOR2_X1   g649(.A(KEYINPUT112), .B(G2090), .Z(new_n1075));
  NAND2_X1  g650(.A1(new_n1029), .A2(new_n1027), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1072), .A2(KEYINPUT45), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1076), .A2(new_n1026), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G1971), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1074), .A2(new_n1075), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  OR2_X1    g655(.A1(new_n1080), .A2(new_n1056), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT55), .ZN(new_n1083));
  NOR3_X1   g658(.A1(G166), .A2(new_n1083), .A3(new_n1056), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  OR2_X1    g660(.A1(new_n1056), .A2(KEYINPUT119), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1081), .A2(new_n1087), .ZN(new_n1088));
  OR3_X1    g663(.A1(new_n1087), .A2(new_n1080), .A3(new_n1056), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1061), .A2(new_n1057), .A3(new_n1063), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT115), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT52), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n966), .A2(G1976), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .A4(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1061), .A2(new_n1057), .A3(new_n1093), .A4(new_n1063), .ZN(new_n1097));
  OAI21_X1  g672(.A(KEYINPUT115), .B1(new_n1097), .B2(new_n1094), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1069), .A2(new_n1090), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT50), .B1(new_n499), .B2(new_n1028), .ZN(new_n1102));
  AOI211_X1 g677(.A(new_n1070), .B(G1384), .C1(new_n493), .C2(new_n498), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1026), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1101), .B1(new_n1104), .B2(G2084), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1106));
  INV_X1    g681(.A(G2084), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1106), .A2(KEYINPUT120), .A3(new_n1107), .A4(new_n1026), .ZN(new_n1108));
  INV_X1    g683(.A(G1966), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1078), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1105), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(G168), .A2(new_n1056), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT51), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1111), .A2(G8), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1112), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1114), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  AOI211_X1 g692(.A(KEYINPUT51), .B(new_n1112), .C1(new_n1111), .C2(G8), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1113), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  OR2_X1    g694(.A1(new_n1078), .A2(G2078), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT53), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1120), .A2(new_n1121), .B1(new_n723), .B2(new_n1104), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1022), .A2(new_n1121), .A3(G2078), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1076), .A2(new_n1077), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  XOR2_X1   g700(.A(G301), .B(KEYINPUT54), .Z(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1122), .B1(new_n1121), .B2(new_n1120), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1127), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1104), .A2(new_n791), .B1(new_n1055), .B2(new_n1034), .ZN(new_n1130));
  OR2_X1    g705(.A1(new_n1130), .A2(KEYINPUT60), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1104), .A2(new_n791), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1055), .A2(new_n1034), .ZN(new_n1133));
  AND4_X1   g708(.A1(KEYINPUT60), .A2(new_n1132), .A3(new_n602), .A4(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n602), .B1(new_n1130), .B2(KEYINPUT60), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1131), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g711(.A(KEYINPUT58), .B(G1341), .ZN(new_n1137));
  OAI22_X1  g712(.A1(new_n1078), .A2(G1996), .B1(new_n1055), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n553), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT59), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT59), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1138), .A2(new_n1141), .A3(new_n553), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(G1956), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1104), .A2(new_n1144), .ZN(new_n1145));
  XOR2_X1   g720(.A(KEYINPUT123), .B(G2072), .Z(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(KEYINPUT56), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1076), .A2(new_n1026), .A3(new_n1077), .A4(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(KEYINPUT122), .B1(new_n611), .B2(new_n613), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT122), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n568), .A2(new_n1151), .A3(new_n570), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1150), .A2(KEYINPUT57), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT57), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1149), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT57), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n611), .A2(new_n613), .A3(KEYINPUT122), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1151), .B1(new_n568), .B2(new_n570), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1156), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1150), .A2(new_n1152), .A3(KEYINPUT57), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1159), .A2(new_n1145), .A3(new_n1148), .A4(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1155), .A2(new_n1161), .A3(KEYINPUT61), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1136), .A2(new_n1143), .A3(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT61), .ZN(new_n1164));
  OR2_X1    g739(.A1(new_n1161), .A2(KEYINPUT124), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1161), .A2(KEYINPUT124), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1165), .A2(new_n1155), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1163), .B1(new_n1164), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1155), .B1(new_n602), .B2(new_n1130), .ZN(new_n1169));
  AND3_X1   g744(.A1(new_n1165), .A2(new_n1169), .A3(new_n1166), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1119), .B(new_n1129), .C1(new_n1168), .C2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1119), .A2(KEYINPUT62), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n1173));
  OAI211_X1 g748(.A(new_n1173), .B(new_n1113), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1172), .A2(G171), .A3(new_n1128), .A4(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1100), .B1(new_n1171), .B2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1111), .A2(G8), .A3(G168), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1177), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1069), .A2(new_n1090), .A3(new_n1099), .A4(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT63), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1082), .A2(new_n1084), .A3(KEYINPUT121), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1081), .A2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1183), .A2(new_n1177), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1180), .B1(new_n1081), .B2(new_n1182), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1184), .A2(new_n1069), .A3(new_n1099), .A4(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1181), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT118), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1081), .A2(new_n1085), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1069), .A2(new_n1099), .A3(new_n1189), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1059), .A2(new_n797), .A3(new_n966), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1191), .A2(new_n1048), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1192), .A2(new_n1057), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1188), .B1(new_n1190), .B2(new_n1193), .ZN(new_n1194));
  AND3_X1   g769(.A1(new_n1190), .A2(new_n1188), .A3(new_n1193), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1187), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1044), .B1(new_n1176), .B2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1031), .B1(new_n740), .B2(new_n1035), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1031), .A2(KEYINPUT46), .A3(new_n1032), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT46), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1200), .B1(new_n1030), .B2(G1996), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1198), .A2(new_n1199), .A3(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1202), .B(KEYINPUT125), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1203), .B(KEYINPUT47), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n714), .A2(new_n1034), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1205), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1206), .A2(new_n1031), .ZN(new_n1207));
  NOR2_X1   g782(.A1(new_n1041), .A2(new_n1030), .ZN(new_n1208));
  XNOR2_X1  g783(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1209));
  XNOR2_X1  g784(.A(new_n1208), .B(new_n1209), .ZN(new_n1210));
  OAI21_X1  g785(.A(new_n1210), .B1(new_n1040), .B2(new_n1030), .ZN(new_n1211));
  AND3_X1   g786(.A1(new_n1204), .A2(new_n1207), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1197), .A2(new_n1212), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g788(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1215));
  NAND2_X1  g789(.A1(new_n1215), .A2(KEYINPUT43), .ZN(new_n1216));
  INV_X1    g790(.A(new_n1019), .ZN(new_n1217));
  NAND2_X1  g791(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g792(.A(G227), .ZN(new_n1219));
  NAND3_X1  g793(.A1(new_n670), .A2(G319), .A3(new_n1219), .ZN(new_n1220));
  INV_X1    g794(.A(KEYINPUT127), .ZN(new_n1221));
  NAND2_X1  g795(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NAND4_X1  g796(.A1(new_n670), .A2(KEYINPUT127), .A3(G319), .A4(new_n1219), .ZN(new_n1223));
  NAND2_X1  g797(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g798(.A(G229), .B1(new_n921), .B2(new_n924), .ZN(new_n1225));
  AND3_X1   g799(.A1(new_n1218), .A2(new_n1224), .A3(new_n1225), .ZN(G308));
  NAND3_X1  g800(.A1(new_n1218), .A2(new_n1224), .A3(new_n1225), .ZN(G225));
endmodule


