

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X4 U547 ( .A1(n518), .A2(n519), .ZN(n884) );
  NOR2_X1 U548 ( .A1(n627), .A2(n934), .ZN(n620) );
  BUF_X2 U549 ( .A(n608), .Z(n648) );
  NOR2_X2 U550 ( .A1(G2104), .A2(G2105), .ZN(n515) );
  BUF_X1 U551 ( .A(n518), .Z(n520) );
  NAND2_X1 U552 ( .A1(n596), .A2(n595), .ZN(n939) );
  NOR2_X1 U553 ( .A1(G651), .A2(n563), .ZN(n794) );
  NAND2_X1 U554 ( .A1(n757), .A2(n756), .ZN(n759) );
  AND2_X1 U555 ( .A1(n927), .A2(n681), .ZN(n513) );
  XNOR2_X1 U556 ( .A(KEYINPUT65), .B(KEYINPUT26), .ZN(n514) );
  XNOR2_X1 U557 ( .A(n606), .B(n514), .ZN(n607) );
  INV_X1 U558 ( .A(KEYINPUT100), .ZN(n619) );
  INV_X1 U559 ( .A(KEYINPUT103), .ZN(n630) );
  XNOR2_X1 U560 ( .A(n651), .B(KEYINPUT30), .ZN(n652) );
  INV_X1 U561 ( .A(KEYINPUT29), .ZN(n641) );
  XNOR2_X1 U562 ( .A(n604), .B(KEYINPUT64), .ZN(n608) );
  INV_X1 U563 ( .A(KEYINPUT107), .ZN(n679) );
  INV_X1 U564 ( .A(KEYINPUT75), .ZN(n588) );
  INV_X1 U565 ( .A(n919), .ZN(n686) );
  XNOR2_X1 U566 ( .A(n589), .B(n588), .ZN(n590) );
  INV_X1 U567 ( .A(G651), .ZN(n529) );
  NOR2_X1 U568 ( .A1(n594), .A2(n593), .ZN(n596) );
  NOR2_X1 U569 ( .A1(G651), .A2(G543), .ZN(n799) );
  XNOR2_X1 U570 ( .A(n602), .B(KEYINPUT68), .ZN(n761) );
  INV_X1 U571 ( .A(KEYINPUT40), .ZN(n758) );
  XNOR2_X1 U572 ( .A(n759), .B(n758), .ZN(G329) );
  XOR2_X2 U573 ( .A(KEYINPUT17), .B(n515), .Z(n883) );
  NAND2_X1 U574 ( .A1(G138), .A2(n883), .ZN(n517) );
  XNOR2_X2 U575 ( .A(G2104), .B(KEYINPUT66), .ZN(n518) );
  INV_X1 U576 ( .A(G2105), .ZN(n519) );
  NAND2_X1 U577 ( .A1(G102), .A2(n884), .ZN(n516) );
  NAND2_X1 U578 ( .A1(n517), .A2(n516), .ZN(n524) );
  AND2_X1 U579 ( .A1(G2104), .A2(G2105), .ZN(n887) );
  NAND2_X1 U580 ( .A1(G114), .A2(n887), .ZN(n522) );
  NOR2_X4 U581 ( .A1(n520), .A2(n519), .ZN(n888) );
  NAND2_X1 U582 ( .A1(G126), .A2(n888), .ZN(n521) );
  NAND2_X1 U583 ( .A1(n522), .A2(n521), .ZN(n523) );
  NOR2_X1 U584 ( .A1(n524), .A2(n523), .ZN(G164) );
  NAND2_X1 U585 ( .A1(n799), .A2(G91), .ZN(n528) );
  NOR2_X1 U586 ( .A1(G543), .A2(n529), .ZN(n525) );
  XOR2_X1 U587 ( .A(KEYINPUT70), .B(n525), .Z(n526) );
  XNOR2_X2 U588 ( .A(KEYINPUT1), .B(n526), .ZN(n795) );
  NAND2_X1 U589 ( .A1(G65), .A2(n795), .ZN(n527) );
  NAND2_X1 U590 ( .A1(n528), .A2(n527), .ZN(n532) );
  XOR2_X1 U591 ( .A(KEYINPUT0), .B(G543), .Z(n563) );
  NOR2_X2 U592 ( .A1(n563), .A2(n529), .ZN(n798) );
  NAND2_X1 U593 ( .A1(G78), .A2(n798), .ZN(n530) );
  XNOR2_X1 U594 ( .A(KEYINPUT73), .B(n530), .ZN(n531) );
  NOR2_X1 U595 ( .A1(n532), .A2(n531), .ZN(n534) );
  NAND2_X1 U596 ( .A1(n794), .A2(G53), .ZN(n533) );
  NAND2_X1 U597 ( .A1(n534), .A2(n533), .ZN(G299) );
  NAND2_X1 U598 ( .A1(n794), .A2(G52), .ZN(n536) );
  NAND2_X1 U599 ( .A1(G64), .A2(n795), .ZN(n535) );
  NAND2_X1 U600 ( .A1(n536), .A2(n535), .ZN(n542) );
  NAND2_X1 U601 ( .A1(n799), .A2(G90), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n537), .B(KEYINPUT72), .ZN(n539) );
  NAND2_X1 U603 ( .A1(G77), .A2(n798), .ZN(n538) );
  NAND2_X1 U604 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U605 ( .A(KEYINPUT9), .B(n540), .Z(n541) );
  NOR2_X1 U606 ( .A1(n542), .A2(n541), .ZN(G171) );
  NAND2_X1 U607 ( .A1(n799), .A2(G89), .ZN(n543) );
  XNOR2_X1 U608 ( .A(n543), .B(KEYINPUT4), .ZN(n545) );
  NAND2_X1 U609 ( .A1(G76), .A2(n798), .ZN(n544) );
  NAND2_X1 U610 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n546), .B(KEYINPUT5), .ZN(n551) );
  NAND2_X1 U612 ( .A1(n794), .A2(G51), .ZN(n548) );
  NAND2_X1 U613 ( .A1(G63), .A2(n795), .ZN(n547) );
  NAND2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U615 ( .A(KEYINPUT6), .B(n549), .Z(n550) );
  NAND2_X1 U616 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U617 ( .A(n552), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U618 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U619 ( .A1(G75), .A2(n798), .ZN(n554) );
  NAND2_X1 U620 ( .A1(G88), .A2(n799), .ZN(n553) );
  NAND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(KEYINPUT88), .B(n555), .ZN(n559) );
  NAND2_X1 U623 ( .A1(n794), .A2(G50), .ZN(n557) );
  NAND2_X1 U624 ( .A1(G62), .A2(n795), .ZN(n556) );
  NAND2_X1 U625 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U626 ( .A1(n559), .A2(n558), .ZN(G166) );
  XOR2_X1 U627 ( .A(KEYINPUT92), .B(G166), .Z(G303) );
  NAND2_X1 U628 ( .A1(G49), .A2(n794), .ZN(n561) );
  NAND2_X1 U629 ( .A1(G74), .A2(G651), .ZN(n560) );
  NAND2_X1 U630 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U631 ( .A1(n795), .A2(n562), .ZN(n566) );
  NAND2_X1 U632 ( .A1(G87), .A2(n563), .ZN(n564) );
  XOR2_X1 U633 ( .A(KEYINPUT85), .B(n564), .Z(n565) );
  NAND2_X1 U634 ( .A1(n566), .A2(n565), .ZN(G288) );
  NAND2_X1 U635 ( .A1(G61), .A2(n795), .ZN(n574) );
  XOR2_X1 U636 ( .A(KEYINPUT86), .B(KEYINPUT2), .Z(n568) );
  NAND2_X1 U637 ( .A1(G73), .A2(n798), .ZN(n567) );
  XNOR2_X1 U638 ( .A(n568), .B(n567), .ZN(n572) );
  NAND2_X1 U639 ( .A1(G86), .A2(n799), .ZN(n570) );
  NAND2_X1 U640 ( .A1(G48), .A2(n794), .ZN(n569) );
  NAND2_X1 U641 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U642 ( .A1(n572), .A2(n571), .ZN(n573) );
  NAND2_X1 U643 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U644 ( .A(KEYINPUT87), .B(n575), .Z(G305) );
  NAND2_X1 U645 ( .A1(G72), .A2(n798), .ZN(n576) );
  XNOR2_X1 U646 ( .A(n576), .B(KEYINPUT69), .ZN(n581) );
  NAND2_X1 U647 ( .A1(n794), .A2(G47), .ZN(n578) );
  NAND2_X1 U648 ( .A1(G60), .A2(n795), .ZN(n577) );
  NAND2_X1 U649 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U650 ( .A(KEYINPUT71), .B(n579), .Z(n580) );
  NOR2_X1 U651 ( .A1(n581), .A2(n580), .ZN(n583) );
  NAND2_X1 U652 ( .A1(n799), .A2(G85), .ZN(n582) );
  NAND2_X1 U653 ( .A1(n583), .A2(n582), .ZN(G290) );
  NAND2_X1 U654 ( .A1(n795), .A2(G56), .ZN(n584) );
  XOR2_X1 U655 ( .A(KEYINPUT14), .B(n584), .Z(n594) );
  NAND2_X1 U656 ( .A1(n798), .A2(G68), .ZN(n585) );
  XNOR2_X1 U657 ( .A(KEYINPUT77), .B(n585), .ZN(n591) );
  XOR2_X1 U658 ( .A(KEYINPUT12), .B(KEYINPUT76), .Z(n587) );
  NAND2_X1 U659 ( .A1(G81), .A2(n799), .ZN(n586) );
  XNOR2_X1 U660 ( .A(n587), .B(n586), .ZN(n589) );
  NOR2_X1 U661 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U662 ( .A(n592), .B(KEYINPUT13), .ZN(n593) );
  NAND2_X1 U663 ( .A1(n794), .A2(G43), .ZN(n595) );
  NAND2_X1 U664 ( .A1(G101), .A2(n884), .ZN(n597) );
  XNOR2_X1 U665 ( .A(n597), .B(KEYINPUT23), .ZN(n598) );
  XNOR2_X1 U666 ( .A(n598), .B(KEYINPUT67), .ZN(n760) );
  NAND2_X1 U667 ( .A1(G113), .A2(n887), .ZN(n600) );
  NAND2_X1 U668 ( .A1(G125), .A2(n888), .ZN(n599) );
  AND2_X1 U669 ( .A1(n600), .A2(n599), .ZN(n762) );
  AND2_X1 U670 ( .A1(G40), .A2(n762), .ZN(n601) );
  AND2_X1 U671 ( .A1(n760), .A2(n601), .ZN(n711) );
  NAND2_X1 U672 ( .A1(G137), .A2(n883), .ZN(n602) );
  AND2_X1 U673 ( .A1(n711), .A2(n761), .ZN(n603) );
  NOR2_X1 U674 ( .A1(G164), .A2(G1384), .ZN(n713) );
  NAND2_X1 U675 ( .A1(n603), .A2(n713), .ZN(n604) );
  INV_X1 U676 ( .A(n608), .ZN(n605) );
  NAND2_X1 U677 ( .A1(n605), .A2(G1996), .ZN(n606) );
  NOR2_X1 U678 ( .A1(n939), .A2(n607), .ZN(n610) );
  NAND2_X1 U679 ( .A1(n648), .A2(G1341), .ZN(n609) );
  NAND2_X1 U680 ( .A1(n610), .A2(n609), .ZN(n627) );
  NAND2_X1 U681 ( .A1(n794), .A2(G54), .ZN(n617) );
  NAND2_X1 U682 ( .A1(n799), .A2(G92), .ZN(n612) );
  NAND2_X1 U683 ( .A1(G66), .A2(n795), .ZN(n611) );
  NAND2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n615) );
  NAND2_X1 U685 ( .A1(n798), .A2(G79), .ZN(n613) );
  XOR2_X1 U686 ( .A(KEYINPUT78), .B(n613), .Z(n614) );
  NOR2_X1 U687 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U688 ( .A1(n617), .A2(n616), .ZN(n618) );
  XOR2_X1 U689 ( .A(KEYINPUT15), .B(n618), .Z(n934) );
  XNOR2_X1 U690 ( .A(n620), .B(n619), .ZN(n626) );
  NAND2_X1 U691 ( .A1(n648), .A2(G1348), .ZN(n621) );
  XOR2_X1 U692 ( .A(KEYINPUT101), .B(n621), .Z(n623) );
  INV_X1 U693 ( .A(n648), .ZN(n643) );
  NAND2_X1 U694 ( .A1(G2067), .A2(n643), .ZN(n622) );
  NAND2_X1 U695 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U696 ( .A(KEYINPUT102), .B(n624), .ZN(n625) );
  NAND2_X1 U697 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U698 ( .A1(n627), .A2(n934), .ZN(n628) );
  NAND2_X1 U699 ( .A1(n629), .A2(n628), .ZN(n631) );
  XNOR2_X1 U700 ( .A(n631), .B(n630), .ZN(n636) );
  NAND2_X1 U701 ( .A1(G2072), .A2(n643), .ZN(n632) );
  XNOR2_X1 U702 ( .A(n632), .B(KEYINPUT27), .ZN(n634) );
  INV_X1 U703 ( .A(G1956), .ZN(n923) );
  NOR2_X1 U704 ( .A1(n643), .A2(n923), .ZN(n633) );
  NOR2_X1 U705 ( .A1(n634), .A2(n633), .ZN(n637) );
  INV_X1 U706 ( .A(G299), .ZN(n924) );
  NAND2_X1 U707 ( .A1(n637), .A2(n924), .ZN(n635) );
  NAND2_X1 U708 ( .A1(n636), .A2(n635), .ZN(n640) );
  NOR2_X1 U709 ( .A1(n637), .A2(n924), .ZN(n638) );
  XOR2_X1 U710 ( .A(n638), .B(KEYINPUT28), .Z(n639) );
  NAND2_X1 U711 ( .A1(n640), .A2(n639), .ZN(n642) );
  XNOR2_X1 U712 ( .A(n642), .B(n641), .ZN(n647) );
  XNOR2_X1 U713 ( .A(KEYINPUT25), .B(G2078), .ZN(n981) );
  NAND2_X1 U714 ( .A1(n643), .A2(n981), .ZN(n645) );
  OR2_X1 U715 ( .A1(n643), .A2(G1961), .ZN(n644) );
  NAND2_X1 U716 ( .A1(n645), .A2(n644), .ZN(n653) );
  NAND2_X1 U717 ( .A1(n653), .A2(G171), .ZN(n646) );
  NAND2_X1 U718 ( .A1(n647), .A2(n646), .ZN(n658) );
  NAND2_X1 U719 ( .A1(n648), .A2(G8), .ZN(n649) );
  XNOR2_X2 U720 ( .A(n649), .B(KEYINPUT98), .ZN(n698) );
  NOR2_X1 U721 ( .A1(n698), .A2(G1966), .ZN(n670) );
  NOR2_X1 U722 ( .A1(n648), .A2(G2084), .ZN(n667) );
  NOR2_X1 U723 ( .A1(n670), .A2(n667), .ZN(n650) );
  NAND2_X1 U724 ( .A1(G8), .A2(n650), .ZN(n651) );
  NOR2_X1 U725 ( .A1(n652), .A2(G168), .ZN(n655) );
  NOR2_X1 U726 ( .A1(G171), .A2(n653), .ZN(n654) );
  NOR2_X1 U727 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U728 ( .A(KEYINPUT31), .B(n656), .Z(n657) );
  NAND2_X1 U729 ( .A1(n658), .A2(n657), .ZN(n668) );
  NAND2_X1 U730 ( .A1(n668), .A2(G286), .ZN(n659) );
  XNOR2_X1 U731 ( .A(n659), .B(KEYINPUT104), .ZN(n664) );
  NOR2_X1 U732 ( .A1(n698), .A2(G1971), .ZN(n661) );
  NOR2_X1 U733 ( .A1(n648), .A2(G2090), .ZN(n660) );
  NOR2_X1 U734 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U735 ( .A1(n662), .A2(G303), .ZN(n663) );
  NAND2_X1 U736 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U737 ( .A1(n665), .A2(G8), .ZN(n666) );
  XNOR2_X1 U738 ( .A(n666), .B(KEYINPUT32), .ZN(n674) );
  NAND2_X1 U739 ( .A1(G8), .A2(n667), .ZN(n672) );
  INV_X1 U740 ( .A(n668), .ZN(n669) );
  NOR2_X1 U741 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U742 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U743 ( .A1(n674), .A2(n673), .ZN(n694) );
  NOR2_X1 U744 ( .A1(G1976), .A2(G288), .ZN(n926) );
  NOR2_X1 U745 ( .A1(G303), .A2(G1971), .ZN(n675) );
  XOR2_X1 U746 ( .A(n675), .B(KEYINPUT105), .Z(n676) );
  NOR2_X1 U747 ( .A1(n926), .A2(n676), .ZN(n677) );
  XNOR2_X1 U748 ( .A(n677), .B(KEYINPUT106), .ZN(n678) );
  NAND2_X1 U749 ( .A1(n694), .A2(n678), .ZN(n680) );
  XNOR2_X1 U750 ( .A(n680), .B(n679), .ZN(n682) );
  NAND2_X1 U751 ( .A1(G1976), .A2(G288), .ZN(n927) );
  INV_X1 U752 ( .A(n698), .ZN(n681) );
  NAND2_X1 U753 ( .A1(n682), .A2(n513), .ZN(n684) );
  INV_X1 U754 ( .A(KEYINPUT33), .ZN(n683) );
  NAND2_X1 U755 ( .A1(n684), .A2(n683), .ZN(n689) );
  NAND2_X1 U756 ( .A1(n926), .A2(KEYINPUT33), .ZN(n685) );
  NOR2_X1 U757 ( .A1(n698), .A2(n685), .ZN(n687) );
  XOR2_X1 U758 ( .A(G1981), .B(G305), .Z(n919) );
  NOR2_X1 U759 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U760 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U761 ( .A(n690), .B(KEYINPUT108), .ZN(n747) );
  NOR2_X1 U762 ( .A1(G1981), .A2(G305), .ZN(n691) );
  XNOR2_X1 U763 ( .A(KEYINPUT24), .B(n691), .ZN(n692) );
  XNOR2_X1 U764 ( .A(KEYINPUT99), .B(n692), .ZN(n693) );
  OR2_X1 U765 ( .A1(n698), .A2(n693), .ZN(n745) );
  NOR2_X1 U766 ( .A1(G2090), .A2(G303), .ZN(n695) );
  NAND2_X1 U767 ( .A1(G8), .A2(n695), .ZN(n696) );
  NAND2_X1 U768 ( .A1(n694), .A2(n696), .ZN(n697) );
  NAND2_X1 U769 ( .A1(n698), .A2(n697), .ZN(n743) );
  XOR2_X1 U770 ( .A(G2067), .B(KEYINPUT37), .Z(n738) );
  NAND2_X1 U771 ( .A1(G140), .A2(n883), .ZN(n700) );
  NAND2_X1 U772 ( .A1(G104), .A2(n884), .ZN(n699) );
  NAND2_X1 U773 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U774 ( .A(KEYINPUT34), .B(n701), .ZN(n708) );
  XNOR2_X1 U775 ( .A(KEYINPUT35), .B(KEYINPUT94), .ZN(n706) );
  NAND2_X1 U776 ( .A1(n887), .A2(G116), .ZN(n704) );
  NAND2_X1 U777 ( .A1(n888), .A2(G128), .ZN(n702) );
  XOR2_X1 U778 ( .A(KEYINPUT93), .B(n702), .Z(n703) );
  NAND2_X1 U779 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U780 ( .A(n706), .B(n705), .Z(n707) );
  NOR2_X1 U781 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U782 ( .A(n709), .B(KEYINPUT36), .Z(n710) );
  XOR2_X1 U783 ( .A(KEYINPUT95), .B(n710), .Z(n894) );
  AND2_X1 U784 ( .A1(n738), .A2(n894), .ZN(n1016) );
  NAND2_X1 U785 ( .A1(n761), .A2(n711), .ZN(n712) );
  NOR2_X1 U786 ( .A1(n713), .A2(n712), .ZN(n750) );
  NAND2_X1 U787 ( .A1(n1016), .A2(n750), .ZN(n752) );
  INV_X1 U788 ( .A(n752), .ZN(n742) );
  INV_X1 U789 ( .A(G1996), .ZN(n729) );
  NAND2_X1 U790 ( .A1(G105), .A2(n884), .ZN(n714) );
  XNOR2_X1 U791 ( .A(n714), .B(KEYINPUT38), .ZN(n716) );
  NAND2_X1 U792 ( .A1(n883), .A2(G141), .ZN(n715) );
  NAND2_X1 U793 ( .A1(n716), .A2(n715), .ZN(n720) );
  NAND2_X1 U794 ( .A1(G117), .A2(n887), .ZN(n718) );
  NAND2_X1 U795 ( .A1(G129), .A2(n888), .ZN(n717) );
  NAND2_X1 U796 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U797 ( .A1(n720), .A2(n719), .ZN(n863) );
  AND2_X1 U798 ( .A1(n729), .A2(n863), .ZN(n995) );
  NAND2_X1 U799 ( .A1(G107), .A2(n887), .ZN(n721) );
  XNOR2_X1 U800 ( .A(n721), .B(KEYINPUT96), .ZN(n724) );
  NAND2_X1 U801 ( .A1(G131), .A2(n883), .ZN(n722) );
  XOR2_X1 U802 ( .A(KEYINPUT97), .B(n722), .Z(n723) );
  NAND2_X1 U803 ( .A1(n724), .A2(n723), .ZN(n728) );
  NAND2_X1 U804 ( .A1(G95), .A2(n884), .ZN(n726) );
  NAND2_X1 U805 ( .A1(G119), .A2(n888), .ZN(n725) );
  NAND2_X1 U806 ( .A1(n726), .A2(n725), .ZN(n727) );
  OR2_X1 U807 ( .A1(n728), .A2(n727), .ZN(n864) );
  AND2_X1 U808 ( .A1(n864), .A2(G1991), .ZN(n731) );
  NOR2_X1 U809 ( .A1(n729), .A2(n863), .ZN(n730) );
  NOR2_X1 U810 ( .A1(n731), .A2(n730), .ZN(n749) );
  INV_X1 U811 ( .A(n749), .ZN(n1005) );
  NOR2_X1 U812 ( .A1(G1986), .A2(G290), .ZN(n732) );
  NOR2_X1 U813 ( .A1(G1991), .A2(n864), .ZN(n1000) );
  NOR2_X1 U814 ( .A1(n732), .A2(n1000), .ZN(n733) );
  XOR2_X1 U815 ( .A(KEYINPUT109), .B(n733), .Z(n734) );
  NOR2_X1 U816 ( .A1(n1005), .A2(n734), .ZN(n735) );
  NOR2_X1 U817 ( .A1(n995), .A2(n735), .ZN(n736) );
  XNOR2_X1 U818 ( .A(KEYINPUT39), .B(n736), .ZN(n737) );
  NAND2_X1 U819 ( .A1(n737), .A2(n750), .ZN(n740) );
  NOR2_X1 U820 ( .A1(n738), .A2(n894), .ZN(n1012) );
  NAND2_X1 U821 ( .A1(n1012), .A2(n750), .ZN(n739) );
  AND2_X1 U822 ( .A1(n740), .A2(n739), .ZN(n741) );
  OR2_X1 U823 ( .A1(n742), .A2(n741), .ZN(n748) );
  AND2_X1 U824 ( .A1(n743), .A2(n748), .ZN(n744) );
  AND2_X1 U825 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U826 ( .A1(n747), .A2(n746), .ZN(n757) );
  INV_X1 U827 ( .A(n748), .ZN(n755) );
  XOR2_X1 U828 ( .A(G1986), .B(G290), .Z(n931) );
  NAND2_X1 U829 ( .A1(n931), .A2(n749), .ZN(n751) );
  NAND2_X1 U830 ( .A1(n751), .A2(n750), .ZN(n753) );
  AND2_X1 U831 ( .A1(n753), .A2(n752), .ZN(n754) );
  OR2_X1 U832 ( .A1(n755), .A2(n754), .ZN(n756) );
  AND2_X1 U833 ( .A1(n761), .A2(n760), .ZN(n763) );
  AND2_X1 U834 ( .A1(n763), .A2(n762), .ZN(G160) );
  AND2_X1 U835 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U836 ( .A(G132), .ZN(G219) );
  INV_X1 U837 ( .A(G57), .ZN(G237) );
  NAND2_X1 U838 ( .A1(G7), .A2(G661), .ZN(n764) );
  XNOR2_X1 U839 ( .A(n764), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U840 ( .A(G223), .ZN(n831) );
  NAND2_X1 U841 ( .A1(n831), .A2(G567), .ZN(n765) );
  XOR2_X1 U842 ( .A(KEYINPUT11), .B(n765), .Z(G234) );
  INV_X1 U843 ( .A(n939), .ZN(n766) );
  NAND2_X1 U844 ( .A1(n766), .A2(G860), .ZN(G153) );
  INV_X1 U845 ( .A(G171), .ZN(G301) );
  NAND2_X1 U846 ( .A1(G868), .A2(G301), .ZN(n768) );
  INV_X1 U847 ( .A(n934), .ZN(n792) );
  OR2_X1 U848 ( .A1(n792), .A2(G868), .ZN(n767) );
  NAND2_X1 U849 ( .A1(n768), .A2(n767), .ZN(G284) );
  XNOR2_X1 U850 ( .A(KEYINPUT79), .B(G868), .ZN(n769) );
  NOR2_X1 U851 ( .A1(G286), .A2(n769), .ZN(n771) );
  NOR2_X1 U852 ( .A1(G868), .A2(G299), .ZN(n770) );
  NOR2_X1 U853 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U854 ( .A(KEYINPUT80), .B(n772), .ZN(G297) );
  INV_X1 U855 ( .A(G559), .ZN(n773) );
  NOR2_X1 U856 ( .A1(G860), .A2(n773), .ZN(n774) );
  XNOR2_X1 U857 ( .A(KEYINPUT81), .B(n774), .ZN(n775) );
  NAND2_X1 U858 ( .A1(n775), .A2(n792), .ZN(n776) );
  XNOR2_X1 U859 ( .A(n776), .B(KEYINPUT83), .ZN(n778) );
  XOR2_X1 U860 ( .A(KEYINPUT16), .B(KEYINPUT82), .Z(n777) );
  XNOR2_X1 U861 ( .A(n778), .B(n777), .ZN(G148) );
  NOR2_X1 U862 ( .A1(G868), .A2(n939), .ZN(n779) );
  XNOR2_X1 U863 ( .A(KEYINPUT84), .B(n779), .ZN(n782) );
  NAND2_X1 U864 ( .A1(G868), .A2(n792), .ZN(n780) );
  NOR2_X1 U865 ( .A1(G559), .A2(n780), .ZN(n781) );
  NOR2_X1 U866 ( .A1(n782), .A2(n781), .ZN(G282) );
  NAND2_X1 U867 ( .A1(G135), .A2(n883), .ZN(n784) );
  NAND2_X1 U868 ( .A1(G111), .A2(n887), .ZN(n783) );
  NAND2_X1 U869 ( .A1(n784), .A2(n783), .ZN(n789) );
  NAND2_X1 U870 ( .A1(G123), .A2(n888), .ZN(n785) );
  XNOR2_X1 U871 ( .A(n785), .B(KEYINPUT18), .ZN(n787) );
  NAND2_X1 U872 ( .A1(n884), .A2(G99), .ZN(n786) );
  NAND2_X1 U873 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U874 ( .A1(n789), .A2(n788), .ZN(n999) );
  XNOR2_X1 U875 ( .A(n999), .B(G2096), .ZN(n791) );
  INV_X1 U876 ( .A(G2100), .ZN(n790) );
  NAND2_X1 U877 ( .A1(n791), .A2(n790), .ZN(G156) );
  NAND2_X1 U878 ( .A1(G559), .A2(n792), .ZN(n793) );
  XNOR2_X1 U879 ( .A(n939), .B(n793), .ZN(n812) );
  NOR2_X1 U880 ( .A1(n812), .A2(G860), .ZN(n804) );
  NAND2_X1 U881 ( .A1(n794), .A2(G55), .ZN(n797) );
  NAND2_X1 U882 ( .A1(G67), .A2(n795), .ZN(n796) );
  NAND2_X1 U883 ( .A1(n797), .A2(n796), .ZN(n803) );
  NAND2_X1 U884 ( .A1(G80), .A2(n798), .ZN(n801) );
  NAND2_X1 U885 ( .A1(G93), .A2(n799), .ZN(n800) );
  NAND2_X1 U886 ( .A1(n801), .A2(n800), .ZN(n802) );
  NOR2_X1 U887 ( .A1(n803), .A2(n802), .ZN(n808) );
  XNOR2_X1 U888 ( .A(n804), .B(n808), .ZN(G145) );
  NOR2_X1 U889 ( .A1(G868), .A2(n808), .ZN(n805) );
  XNOR2_X1 U890 ( .A(n805), .B(KEYINPUT89), .ZN(n815) );
  XOR2_X1 U891 ( .A(G166), .B(KEYINPUT19), .Z(n806) );
  XNOR2_X1 U892 ( .A(G288), .B(n806), .ZN(n807) );
  XNOR2_X1 U893 ( .A(n808), .B(n807), .ZN(n810) );
  XNOR2_X1 U894 ( .A(G305), .B(n924), .ZN(n809) );
  XNOR2_X1 U895 ( .A(n810), .B(n809), .ZN(n811) );
  XNOR2_X1 U896 ( .A(n811), .B(G290), .ZN(n898) );
  XOR2_X1 U897 ( .A(n898), .B(n812), .Z(n813) );
  NAND2_X1 U898 ( .A1(G868), .A2(n813), .ZN(n814) );
  NAND2_X1 U899 ( .A1(n815), .A2(n814), .ZN(G295) );
  NAND2_X1 U900 ( .A1(G2078), .A2(G2084), .ZN(n816) );
  XOR2_X1 U901 ( .A(KEYINPUT20), .B(n816), .Z(n817) );
  NAND2_X1 U902 ( .A1(G2090), .A2(n817), .ZN(n818) );
  XNOR2_X1 U903 ( .A(KEYINPUT21), .B(n818), .ZN(n819) );
  NAND2_X1 U904 ( .A1(n819), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U905 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U906 ( .A(KEYINPUT74), .B(G82), .Z(G220) );
  NAND2_X1 U907 ( .A1(G69), .A2(G120), .ZN(n820) );
  NOR2_X1 U908 ( .A1(G237), .A2(n820), .ZN(n821) );
  NAND2_X1 U909 ( .A1(G108), .A2(n821), .ZN(n836) );
  NAND2_X1 U910 ( .A1(G567), .A2(n836), .ZN(n822) );
  XNOR2_X1 U911 ( .A(KEYINPUT91), .B(n822), .ZN(n828) );
  NOR2_X1 U912 ( .A1(G220), .A2(G219), .ZN(n823) );
  XOR2_X1 U913 ( .A(KEYINPUT22), .B(n823), .Z(n824) );
  NOR2_X1 U914 ( .A1(G218), .A2(n824), .ZN(n825) );
  NAND2_X1 U915 ( .A1(G96), .A2(n825), .ZN(n835) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n835), .ZN(n826) );
  XOR2_X1 U917 ( .A(KEYINPUT90), .B(n826), .Z(n827) );
  NOR2_X1 U918 ( .A1(n828), .A2(n827), .ZN(G319) );
  INV_X1 U919 ( .A(G319), .ZN(n830) );
  NAND2_X1 U920 ( .A1(G483), .A2(G661), .ZN(n829) );
  NOR2_X1 U921 ( .A1(n830), .A2(n829), .ZN(n834) );
  NAND2_X1 U922 ( .A1(n834), .A2(G36), .ZN(G176) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n831), .ZN(G217) );
  AND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n832) );
  NAND2_X1 U925 ( .A1(G661), .A2(n832), .ZN(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n833) );
  NAND2_X1 U927 ( .A1(n834), .A2(n833), .ZN(G188) );
  INV_X1 U929 ( .A(G120), .ZN(G236) );
  INV_X1 U930 ( .A(G96), .ZN(G221) );
  INV_X1 U931 ( .A(G69), .ZN(G235) );
  NOR2_X1 U932 ( .A1(n836), .A2(n835), .ZN(G325) );
  INV_X1 U933 ( .A(G325), .ZN(G261) );
  XOR2_X1 U934 ( .A(KEYINPUT41), .B(G1991), .Z(n838) );
  XNOR2_X1 U935 ( .A(G1956), .B(G1996), .ZN(n837) );
  XNOR2_X1 U936 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U937 ( .A(n839), .B(KEYINPUT111), .Z(n841) );
  XNOR2_X1 U938 ( .A(G1981), .B(G1966), .ZN(n840) );
  XNOR2_X1 U939 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U940 ( .A(G1986), .B(G1976), .Z(n843) );
  XNOR2_X1 U941 ( .A(G1961), .B(G1971), .ZN(n842) );
  XNOR2_X1 U942 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U943 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U944 ( .A(KEYINPUT110), .B(G2474), .ZN(n846) );
  XNOR2_X1 U945 ( .A(n847), .B(n846), .ZN(G229) );
  XOR2_X1 U946 ( .A(G2678), .B(KEYINPUT42), .Z(n849) );
  XNOR2_X1 U947 ( .A(G2096), .B(G2100), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U949 ( .A(KEYINPUT43), .B(G2090), .Z(n851) );
  XNOR2_X1 U950 ( .A(G2072), .B(G2067), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U952 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U953 ( .A(G2078), .B(G2084), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(G227) );
  NAND2_X1 U955 ( .A1(G136), .A2(n883), .ZN(n857) );
  NAND2_X1 U956 ( .A1(G112), .A2(n887), .ZN(n856) );
  NAND2_X1 U957 ( .A1(n857), .A2(n856), .ZN(n862) );
  NAND2_X1 U958 ( .A1(G124), .A2(n888), .ZN(n858) );
  XNOR2_X1 U959 ( .A(n858), .B(KEYINPUT44), .ZN(n860) );
  NAND2_X1 U960 ( .A1(n884), .A2(G100), .ZN(n859) );
  NAND2_X1 U961 ( .A1(n860), .A2(n859), .ZN(n861) );
  NOR2_X1 U962 ( .A1(n862), .A2(n861), .ZN(G162) );
  XOR2_X1 U963 ( .A(G162), .B(n999), .Z(n866) );
  XOR2_X1 U964 ( .A(n864), .B(n863), .Z(n865) );
  XNOR2_X1 U965 ( .A(n866), .B(n865), .ZN(n870) );
  XOR2_X1 U966 ( .A(KEYINPUT46), .B(KEYINPUT113), .Z(n868) );
  XNOR2_X1 U967 ( .A(KEYINPUT114), .B(KEYINPUT48), .ZN(n867) );
  XNOR2_X1 U968 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U969 ( .A(n870), .B(n869), .Z(n872) );
  XNOR2_X1 U970 ( .A(G160), .B(G164), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(n882) );
  NAND2_X1 U972 ( .A1(G142), .A2(n883), .ZN(n874) );
  NAND2_X1 U973 ( .A1(G106), .A2(n884), .ZN(n873) );
  NAND2_X1 U974 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U975 ( .A(n875), .B(KEYINPUT45), .ZN(n877) );
  NAND2_X1 U976 ( .A1(G130), .A2(n888), .ZN(n876) );
  NAND2_X1 U977 ( .A1(n877), .A2(n876), .ZN(n880) );
  NAND2_X1 U978 ( .A1(n887), .A2(G118), .ZN(n878) );
  XOR2_X1 U979 ( .A(KEYINPUT112), .B(n878), .Z(n879) );
  NOR2_X1 U980 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U981 ( .A(n882), .B(n881), .Z(n896) );
  NAND2_X1 U982 ( .A1(G139), .A2(n883), .ZN(n886) );
  NAND2_X1 U983 ( .A1(G103), .A2(n884), .ZN(n885) );
  NAND2_X1 U984 ( .A1(n886), .A2(n885), .ZN(n893) );
  NAND2_X1 U985 ( .A1(G115), .A2(n887), .ZN(n890) );
  NAND2_X1 U986 ( .A1(G127), .A2(n888), .ZN(n889) );
  NAND2_X1 U987 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U988 ( .A(KEYINPUT47), .B(n891), .Z(n892) );
  NOR2_X1 U989 ( .A1(n893), .A2(n892), .ZN(n1006) );
  XNOR2_X1 U990 ( .A(n894), .B(n1006), .ZN(n895) );
  XNOR2_X1 U991 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U992 ( .A1(G37), .A2(n897), .ZN(G395) );
  XNOR2_X1 U993 ( .A(G171), .B(KEYINPUT115), .ZN(n901) );
  XNOR2_X1 U994 ( .A(n898), .B(n934), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n899), .B(n939), .ZN(n900) );
  XNOR2_X1 U996 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U997 ( .A(n902), .B(G286), .ZN(n903) );
  NOR2_X1 U998 ( .A1(G37), .A2(n903), .ZN(G397) );
  XOR2_X1 U999 ( .A(G2427), .B(G2430), .Z(n905) );
  XNOR2_X1 U1000 ( .A(G2438), .B(G2443), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n911) );
  XOR2_X1 U1002 ( .A(G2435), .B(G2454), .Z(n907) );
  XNOR2_X1 U1003 ( .A(G1341), .B(G1348), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n909) );
  XOR2_X1 U1005 ( .A(G2451), .B(G2446), .Z(n908) );
  XNOR2_X1 U1006 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1007 ( .A(n911), .B(n910), .Z(n912) );
  NAND2_X1 U1008 ( .A1(G14), .A2(n912), .ZN(n918) );
  NAND2_X1 U1009 ( .A1(G319), .A2(n918), .ZN(n915) );
  NOR2_X1 U1010 ( .A1(G229), .A2(G227), .ZN(n913) );
  XNOR2_X1 U1011 ( .A(KEYINPUT49), .B(n913), .ZN(n914) );
  NOR2_X1 U1012 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1014 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(G108), .ZN(G238) );
  INV_X1 U1017 ( .A(n918), .ZN(G401) );
  XNOR2_X1 U1018 ( .A(KEYINPUT56), .B(G16), .ZN(n946) );
  XNOR2_X1 U1019 ( .A(G1966), .B(G168), .ZN(n920) );
  NAND2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1021 ( .A(n921), .B(KEYINPUT57), .ZN(n922) );
  XNOR2_X1 U1022 ( .A(KEYINPUT122), .B(n922), .ZN(n944) );
  XNOR2_X1 U1023 ( .A(n924), .B(n923), .ZN(n925) );
  NOR2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n928) );
  NAND2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n930) );
  XNOR2_X1 U1026 ( .A(G1971), .B(G303), .ZN(n929) );
  NOR2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n932) );
  NAND2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1029 ( .A(n933), .B(KEYINPUT123), .ZN(n938) );
  XNOR2_X1 U1030 ( .A(G301), .B(G1961), .ZN(n936) );
  XNOR2_X1 U1031 ( .A(n934), .B(G1348), .ZN(n935) );
  NOR2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n942) );
  XNOR2_X1 U1034 ( .A(G1341), .B(n939), .ZN(n940) );
  XNOR2_X1 U1035 ( .A(KEYINPUT124), .B(n940), .ZN(n941) );
  NOR2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1037 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1038 ( .A1(n946), .A2(n945), .ZN(n1026) );
  XNOR2_X1 U1039 ( .A(G1348), .B(KEYINPUT59), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(n947), .B(G4), .ZN(n951) );
  XNOR2_X1 U1041 ( .A(G1981), .B(G6), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(G1341), .B(G19), .ZN(n948) );
  NOR2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1044 ( .A1(n951), .A2(n950), .ZN(n954) );
  XOR2_X1 U1045 ( .A(KEYINPUT127), .B(G1956), .Z(n952) );
  XNOR2_X1 U1046 ( .A(G20), .B(n952), .ZN(n953) );
  NOR2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1048 ( .A(KEYINPUT60), .B(n955), .ZN(n965) );
  XNOR2_X1 U1049 ( .A(G1961), .B(KEYINPUT126), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(n956), .B(G5), .ZN(n963) );
  XNOR2_X1 U1051 ( .A(G1971), .B(G22), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(G23), .B(G1976), .ZN(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n960) );
  XOR2_X1 U1054 ( .A(G1986), .B(G24), .Z(n959) );
  NAND2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1056 ( .A(KEYINPUT58), .B(n961), .ZN(n962) );
  NOR2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n967) );
  XNOR2_X1 U1059 ( .A(G21), .B(G1966), .ZN(n966) );
  NOR2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(n968), .B(KEYINPUT61), .ZN(n970) );
  XNOR2_X1 U1062 ( .A(G16), .B(KEYINPUT125), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1064 ( .A1(G11), .A2(n971), .ZN(n1024) );
  XNOR2_X1 U1065 ( .A(G2090), .B(G35), .ZN(n987) );
  XNOR2_X1 U1066 ( .A(KEYINPUT119), .B(G2067), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(n972), .B(G26), .ZN(n980) );
  XNOR2_X1 U1068 ( .A(G2072), .B(G33), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(G1996), .B(G32), .ZN(n973) );
  NOR2_X1 U1070 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1071 ( .A1(G28), .A2(n975), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(G25), .B(G1991), .ZN(n976) );
  XNOR2_X1 U1073 ( .A(KEYINPUT118), .B(n976), .ZN(n977) );
  NOR2_X1 U1074 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n984) );
  XOR2_X1 U1076 ( .A(G27), .B(n981), .Z(n982) );
  XNOR2_X1 U1077 ( .A(KEYINPUT120), .B(n982), .ZN(n983) );
  NOR2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1079 ( .A(KEYINPUT53), .B(n985), .ZN(n986) );
  NOR2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n990) );
  XOR2_X1 U1081 ( .A(G2084), .B(G34), .Z(n988) );
  XNOR2_X1 U1082 ( .A(KEYINPUT54), .B(n988), .ZN(n989) );
  NAND2_X1 U1083 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1084 ( .A(KEYINPUT55), .B(n991), .ZN(n992) );
  NOR2_X1 U1085 ( .A1(G29), .A2(n992), .ZN(n993) );
  XNOR2_X1 U1086 ( .A(n993), .B(KEYINPUT121), .ZN(n1022) );
  XOR2_X1 U1087 ( .A(G160), .B(G2084), .Z(n998) );
  XOR2_X1 U1088 ( .A(G2090), .B(G162), .Z(n994) );
  NOR2_X1 U1089 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1090 ( .A(KEYINPUT51), .B(n996), .ZN(n997) );
  NOR2_X1 U1091 ( .A1(n998), .A2(n997), .ZN(n1003) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1093 ( .A(n1001), .B(KEYINPUT116), .ZN(n1002) );
  NAND2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1014) );
  XNOR2_X1 U1096 ( .A(G2072), .B(n1006), .ZN(n1009) );
  XOR2_X1 U1097 ( .A(G164), .B(G2078), .Z(n1007) );
  XNOR2_X1 U1098 ( .A(KEYINPUT117), .B(n1007), .ZN(n1008) );
  NAND2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(n1010), .B(KEYINPUT50), .ZN(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1104 ( .A(n1017), .B(KEYINPUT52), .ZN(n1019) );
  INV_X1 U1105 ( .A(KEYINPUT55), .ZN(n1018) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1107 ( .A1(G29), .A2(n1020), .ZN(n1021) );
  NAND2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1111 ( .A(KEYINPUT62), .B(n1027), .Z(G311) );
  INV_X1 U1112 ( .A(G311), .ZN(G150) );
endmodule

