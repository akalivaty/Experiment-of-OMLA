//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 0 0 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n548, new_n549, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n573,
    new_n574, new_n575, new_n576, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT65), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT68), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n463), .B1(new_n464), .B2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(KEYINPUT69), .A3(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n464), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G137), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(new_n468), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n478), .A2(G101), .A3(G2104), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n471), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  AND2_X1   g056(.A1(new_n470), .A2(G136), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G112), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n465), .A2(new_n467), .A3(G2105), .A4(new_n468), .ZN(new_n486));
  OR2_X1    g061(.A1(new_n486), .A2(KEYINPUT70), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(KEYINPUT70), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI211_X1 g064(.A(new_n482), .B(new_n485), .C1(new_n489), .C2(G124), .ZN(G162));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n465), .A2(new_n467), .A3(new_n492), .A4(new_n468), .ZN(new_n493));
  AND2_X1   g068(.A1(new_n473), .A2(new_n468), .ZN(new_n494));
  NOR3_X1   g069(.A1(new_n491), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n493), .A2(KEYINPUT4), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G126), .ZN(new_n497));
  OR2_X1    g072(.A1(KEYINPUT71), .A2(G114), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT71), .A2(G114), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n478), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n501));
  OAI22_X1  g076(.A1(new_n486), .A2(new_n497), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n496), .A2(new_n502), .ZN(G164));
  XNOR2_X1  g078(.A(KEYINPUT5), .B(G543), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n508), .A2(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  OAI21_X1  g088(.A(G543), .B1(new_n510), .B2(new_n511), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n507), .A2(new_n516), .ZN(G166));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT7), .ZN(new_n519));
  INV_X1    g094(.A(G51), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n519), .B1(new_n520), .B2(new_n514), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n509), .A2(new_n508), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT6), .B(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G89), .ZN(new_n524));
  NAND2_X1  g099(.A1(G63), .A2(G651), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n522), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n521), .A2(new_n526), .ZN(G168));
  AOI22_X1  g102(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(new_n506), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n504), .A2(new_n523), .A3(G90), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n523), .A2(G52), .A3(G543), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT72), .ZN(new_n532));
  AND3_X1   g107(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n532), .B1(new_n530), .B2(new_n531), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n529), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(G171));
  NAND3_X1  g111(.A1(new_n504), .A2(new_n523), .A3(G81), .ZN(new_n537));
  OR2_X1    g112(.A1(KEYINPUT73), .A2(G43), .ZN(new_n538));
  NAND2_X1  g113(.A1(KEYINPUT73), .A2(G43), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n523), .A2(G543), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(G68), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n542), .B1(new_n504), .B2(G56), .ZN(new_n543));
  OAI211_X1 g118(.A(new_n537), .B(new_n540), .C1(new_n543), .C2(new_n506), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  INV_X1    g125(.A(KEYINPUT75), .ZN(new_n551));
  NAND2_X1  g126(.A1(G78), .A2(G543), .ZN(new_n552));
  OAI21_X1  g127(.A(KEYINPUT74), .B1(new_n509), .B2(new_n508), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT5), .ZN(new_n554));
  INV_X1    g129(.A(G543), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT74), .ZN(new_n557));
  NAND2_X1  g132(.A1(KEYINPUT5), .A2(G543), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AND2_X1   g134(.A1(new_n553), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI211_X1 g136(.A(new_n551), .B(new_n552), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n561), .B1(new_n553), .B2(new_n559), .ZN(new_n563));
  INV_X1    g138(.A(new_n552), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT75), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n562), .A2(G651), .A3(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(G53), .ZN(new_n567));
  OR3_X1    g142(.A1(new_n514), .A2(KEYINPUT9), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g143(.A(KEYINPUT9), .B1(new_n514), .B2(new_n567), .ZN(new_n569));
  INV_X1    g144(.A(new_n512), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n568), .A2(new_n569), .B1(G91), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n566), .A2(new_n571), .ZN(G299));
  NAND2_X1  g147(.A1(new_n535), .A2(KEYINPUT76), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n574));
  OAI211_X1 g149(.A(new_n529), .B(new_n574), .C1(new_n533), .C2(new_n534), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G301));
  INV_X1    g152(.A(G168), .ZN(G286));
  INV_X1    g153(.A(G166), .ZN(G303));
  AND3_X1   g154(.A1(new_n504), .A2(new_n523), .A3(G87), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT77), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n504), .A2(G74), .ZN(new_n582));
  INV_X1    g157(.A(new_n514), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n582), .A2(G651), .B1(new_n583), .B2(G49), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n581), .A2(new_n584), .ZN(G288));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n522), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(G651), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(KEYINPUT78), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n588), .A2(new_n591), .A3(G651), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n570), .A2(G86), .B1(new_n583), .B2(G48), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n590), .A2(new_n592), .A3(new_n593), .ZN(G305));
  AOI22_X1  g169(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n595), .A2(new_n506), .ZN(new_n596));
  INV_X1    g171(.A(G85), .ZN(new_n597));
  INV_X1    g172(.A(G47), .ZN(new_n598));
  OAI22_X1  g173(.A1(new_n512), .A2(new_n597), .B1(new_n514), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G290));
  NAND3_X1  g176(.A1(new_n570), .A2(KEYINPUT10), .A3(G92), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  INV_X1    g178(.A(G92), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n512), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G66), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n607), .B1(new_n553), .B2(new_n559), .ZN(new_n608));
  AND2_X1   g183(.A1(G79), .A2(G543), .ZN(new_n609));
  OAI21_X1  g184(.A(G651), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n583), .A2(G54), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n606), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(new_n576), .B2(G868), .ZN(G284));
  AOI21_X1  g189(.A(new_n613), .B1(new_n576), .B2(G868), .ZN(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n568), .A2(new_n569), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n570), .A2(G91), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n563), .A2(new_n564), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n506), .B1(new_n620), .B2(new_n551), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n619), .B1(new_n621), .B2(new_n565), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n616), .B1(new_n622), .B2(G868), .ZN(G297));
  OAI21_X1  g198(.A(new_n616), .B1(new_n622), .B2(G868), .ZN(G280));
  INV_X1    g199(.A(new_n612), .ZN(new_n625));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G860), .ZN(G148));
  INV_X1    g202(.A(G868), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n544), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n612), .A2(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(new_n628), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g207(.A1(new_n478), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT12), .Z(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT79), .B(KEYINPUT13), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(KEYINPUT80), .B2(G2100), .ZN(new_n637));
  NAND2_X1  g212(.A1(KEYINPUT80), .A2(G2100), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n637), .B(new_n638), .Z(new_n639));
  NAND2_X1  g214(.A1(new_n489), .A2(G123), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n470), .A2(G135), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n642));
  INV_X1    g217(.A(G111), .ZN(new_n643));
  AOI22_X1  g218(.A1(new_n642), .A2(KEYINPUT81), .B1(new_n643), .B2(G2105), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(KEYINPUT81), .B2(new_n642), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n640), .A2(new_n641), .A3(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n646), .A2(G2096), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(G2096), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n639), .A2(new_n647), .A3(new_n648), .ZN(G156));
  XNOR2_X1  g224(.A(G2427), .B(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2430), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT15), .B(G2435), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(KEYINPUT14), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G1341), .B(G1348), .Z(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n655), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2451), .B(G2454), .Z(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n659), .A2(new_n662), .ZN(new_n664));
  AND3_X1   g239(.A1(new_n663), .A2(G14), .A3(new_n664), .ZN(G401));
  XNOR2_X1  g240(.A(G2072), .B(G2078), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT17), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT84), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n670), .A2(new_n666), .A3(new_n668), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT83), .B(KEYINPUT18), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n667), .A2(new_n668), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n666), .A2(new_n668), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n678), .A2(new_n670), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n673), .B(new_n676), .C1(new_n677), .C2(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G2096), .B(G2100), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(G227));
  XOR2_X1   g257(.A(G1991), .B(G1996), .Z(new_n683));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT19), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1956), .B(G2474), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1961), .B(G1966), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n687), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n685), .A2(KEYINPUT86), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n691), .B(new_n692), .Z(new_n693));
  NOR3_X1   g268(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT85), .B(KEYINPUT20), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n693), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n697), .B1(new_n693), .B2(new_n696), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n683), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n700), .ZN(new_n702));
  INV_X1    g277(.A(new_n683), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n702), .A2(new_n703), .A3(new_n698), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1981), .B(G1986), .ZN(new_n705));
  AND3_X1   g280(.A1(new_n701), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n705), .B1(new_n701), .B2(new_n704), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(G229));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G32), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n489), .A2(G129), .ZN(new_n711));
  INV_X1    g286(.A(G105), .ZN(new_n712));
  NOR3_X1   g287(.A1(new_n712), .A2(new_n466), .A3(G2105), .ZN(new_n713));
  NAND3_X1  g288(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT26), .ZN(new_n715));
  AOI211_X1 g290(.A(new_n713), .B(new_n715), .C1(new_n470), .C2(G141), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n710), .B1(new_n718), .B2(new_n709), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT27), .Z(new_n720));
  INV_X1    g295(.A(G1996), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n709), .A2(G26), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT28), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n489), .A2(G128), .ZN(new_n725));
  OAI21_X1  g300(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n726));
  INV_X1    g301(.A(G116), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n726), .B1(new_n727), .B2(G2105), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n470), .B2(G140), .ZN(new_n729));
  AND3_X1   g304(.A1(new_n725), .A2(KEYINPUT92), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(KEYINPUT92), .B1(new_n725), .B2(new_n729), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n724), .B1(new_n732), .B2(new_n709), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT93), .B(G2067), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n733), .B(new_n734), .Z(new_n735));
  NAND2_X1  g310(.A1(new_n722), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n709), .A2(G35), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G162), .B2(new_n709), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT29), .Z(new_n739));
  INV_X1    g314(.A(G2090), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT96), .ZN(new_n742));
  INV_X1    g317(.A(G16), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G20), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT23), .Z(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G299), .B2(G16), .ZN(new_n746));
  INV_X1    g321(.A(G1956), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n739), .B2(new_n740), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n709), .A2(G33), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n494), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n751), .A2(new_n478), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n478), .A2(G103), .A3(G2104), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT25), .Z(new_n754));
  INV_X1    g329(.A(G139), .ZN(new_n755));
  INV_X1    g330(.A(new_n470), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n752), .B(new_n754), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n750), .B1(new_n757), .B2(G29), .ZN(new_n758));
  INV_X1    g333(.A(G2072), .ZN(new_n759));
  OAI22_X1  g334(.A1(new_n758), .A2(new_n759), .B1(new_n646), .B2(new_n709), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n743), .A2(G21), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G168), .B2(new_n743), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT94), .B(G1966), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n762), .B(new_n763), .Z(new_n764));
  INV_X1    g339(.A(G34), .ZN(new_n765));
  AOI21_X1  g340(.A(G29), .B1(new_n765), .B2(KEYINPUT24), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(KEYINPUT24), .B2(new_n765), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n480), .B2(new_n709), .ZN(new_n768));
  INV_X1    g343(.A(G2084), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR3_X1   g345(.A1(new_n760), .A2(new_n764), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n545), .A2(G16), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G16), .B2(G19), .ZN(new_n773));
  INV_X1    g348(.A(G1341), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT30), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n777), .A2(G28), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n709), .B1(new_n777), .B2(G28), .ZN(new_n779));
  AND2_X1   g354(.A1(KEYINPUT31), .A2(G11), .ZN(new_n780));
  NOR2_X1   g355(.A1(KEYINPUT31), .A2(G11), .ZN(new_n781));
  OAI22_X1  g356(.A1(new_n778), .A2(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n775), .A2(new_n776), .A3(new_n782), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n758), .A2(new_n759), .B1(new_n769), .B2(new_n768), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n771), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n625), .A2(G16), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G4), .B2(G16), .ZN(new_n787));
  INV_X1    g362(.A(G1348), .ZN(new_n788));
  NOR2_X1   g363(.A1(G27), .A2(G29), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G164), .B2(G29), .ZN(new_n790));
  AOI22_X1  g365(.A1(new_n787), .A2(new_n788), .B1(G2078), .B2(new_n790), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n790), .A2(G2078), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n791), .B(new_n792), .C1(new_n788), .C2(new_n787), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n785), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n743), .A2(G5), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G171), .B2(new_n743), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT95), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1961), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n749), .A2(new_n794), .A3(new_n798), .ZN(new_n799));
  NOR3_X1   g374(.A1(new_n736), .A2(new_n742), .A3(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(G1976), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n743), .A2(G23), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n581), .A2(new_n584), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(new_n743), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n805), .A2(KEYINPUT90), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT33), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n805), .A2(KEYINPUT90), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n807), .B1(new_n806), .B2(new_n808), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n802), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT34), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n805), .B(KEYINPUT90), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(KEYINPUT33), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n815), .A2(new_n809), .A3(G1976), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n743), .A2(G22), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G166), .B2(new_n743), .ZN(new_n818));
  INV_X1    g393(.A(G1971), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  AND3_X1   g395(.A1(new_n590), .A2(new_n592), .A3(new_n593), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G16), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G6), .B2(G16), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT32), .B(G1981), .Z(new_n824));
  OAI21_X1  g399(.A(new_n820), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(new_n823), .B2(new_n824), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n812), .A2(new_n813), .A3(new_n816), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n709), .A2(G25), .ZN(new_n828));
  AND3_X1   g403(.A1(new_n487), .A2(G119), .A3(new_n488), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT87), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n830), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n834));
  INV_X1    g409(.A(G107), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n834), .B1(new_n835), .B2(G2105), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(G131), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n837), .B1(new_n756), .B2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n833), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT88), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n828), .B1(new_n842), .B2(new_n709), .ZN(new_n843));
  XOR2_X1   g418(.A(KEYINPUT35), .B(G1991), .Z(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n743), .A2(G24), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n600), .B2(new_n743), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT89), .ZN(new_n849));
  INV_X1    g424(.A(G1986), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(new_n843), .B2(new_n845), .ZN(new_n852));
  AND3_X1   g427(.A1(new_n827), .A2(new_n846), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n812), .A2(new_n816), .A3(new_n826), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT91), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n854), .A2(new_n855), .A3(KEYINPUT34), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n855), .B1(new_n854), .B2(KEYINPUT34), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n853), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(KEYINPUT36), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT36), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n853), .B(new_n861), .C1(new_n857), .C2(new_n858), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n801), .B1(new_n860), .B2(new_n862), .ZN(G311));
  INV_X1    g438(.A(new_n858), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(new_n856), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n861), .B1(new_n865), .B2(new_n853), .ZN(new_n866));
  INV_X1    g441(.A(new_n862), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n800), .B1(new_n866), .B2(new_n867), .ZN(G150));
  INV_X1    g443(.A(G93), .ZN(new_n869));
  INV_X1    g444(.A(G55), .ZN(new_n870));
  OAI22_X1  g445(.A1(new_n512), .A2(new_n869), .B1(new_n514), .B2(new_n870), .ZN(new_n871));
  AOI22_X1  g446(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n872));
  OAI21_X1  g447(.A(KEYINPUT98), .B1(new_n872), .B2(new_n506), .ZN(new_n873));
  OAI21_X1  g448(.A(G67), .B1(new_n509), .B2(new_n508), .ZN(new_n874));
  NAND2_X1  g449(.A1(G80), .A2(G543), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT98), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n876), .A2(new_n877), .A3(G651), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n871), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(G860), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT37), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n612), .A2(new_n626), .ZN(new_n883));
  XOR2_X1   g458(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n884));
  XNOR2_X1  g459(.A(new_n883), .B(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(G56), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n886), .B1(new_n556), .B2(new_n558), .ZN(new_n887));
  OAI21_X1  g462(.A(G651), .B1(new_n887), .B2(new_n542), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n888), .A2(KEYINPUT99), .A3(new_n537), .A4(new_n540), .ZN(new_n889));
  INV_X1    g464(.A(new_n871), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n877), .B1(new_n876), .B2(G651), .ZN(new_n891));
  AOI211_X1 g466(.A(KEYINPUT98), .B(new_n506), .C1(new_n874), .C2(new_n875), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n889), .B(new_n890), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT99), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT100), .ZN(new_n895));
  INV_X1    g470(.A(G81), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n538), .A2(new_n539), .ZN(new_n897));
  OAI22_X1  g472(.A1(new_n512), .A2(new_n896), .B1(new_n514), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(G56), .B1(new_n509), .B2(new_n508), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n506), .B1(new_n899), .B2(new_n541), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n894), .B(new_n895), .C1(new_n898), .C2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n895), .B1(new_n544), .B2(new_n894), .ZN(new_n903));
  NOR3_X1   g478(.A1(new_n893), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n894), .B1(new_n898), .B2(new_n900), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT100), .ZN(new_n906));
  AOI22_X1  g481(.A1(new_n906), .A2(new_n901), .B1(new_n879), .B2(new_n889), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n885), .B(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n910), .A2(KEYINPUT39), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n880), .B1(new_n910), .B2(KEYINPUT39), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n882), .B1(new_n911), .B2(new_n912), .ZN(G145));
  OR2_X1    g488(.A1(G106), .A2(G2105), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n914), .B(G2104), .C1(G118), .C2(new_n478), .ZN(new_n915));
  INV_X1    g490(.A(G142), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n915), .B1(new_n756), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n917), .B1(new_n489), .B2(G130), .ZN(new_n918));
  INV_X1    g493(.A(new_n634), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n919), .B1(new_n833), .B2(new_n840), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  AOI211_X1 g496(.A(new_n634), .B(new_n839), .C1(new_n831), .C2(new_n832), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n918), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n918), .ZN(new_n925));
  NOR3_X1   g500(.A1(new_n920), .A2(new_n922), .A3(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  OAI22_X1  g502(.A1(new_n730), .A2(new_n731), .B1(new_n496), .B2(new_n502), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n725), .A2(new_n729), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT92), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n725), .A2(KEYINPUT92), .A3(new_n729), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(G164), .A3(new_n932), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n928), .A2(new_n933), .A3(new_n757), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n757), .B1(new_n928), .B2(new_n933), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n717), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n928), .A2(new_n933), .ZN(new_n937));
  INV_X1    g512(.A(new_n757), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n928), .A2(new_n933), .A3(new_n757), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n939), .A2(new_n718), .A3(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n927), .A2(new_n936), .A3(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n646), .B(new_n480), .ZN(new_n943));
  XOR2_X1   g518(.A(new_n943), .B(G162), .Z(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n936), .A2(new_n941), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n947), .B1(new_n926), .B2(new_n924), .ZN(new_n948));
  AOI21_X1  g523(.A(G37), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT101), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n942), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n948), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n947), .B(new_n951), .C1(new_n926), .C2(new_n924), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n945), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n950), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n953), .A2(new_n954), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n944), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n956), .B1(new_n960), .B2(new_n949), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n958), .A2(new_n961), .ZN(G395));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n821), .A2(G166), .ZN(new_n964));
  NAND2_X1  g539(.A1(G303), .A2(G305), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT106), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT106), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n964), .A2(new_n968), .A3(new_n965), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT105), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n581), .A2(new_n970), .A3(new_n584), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n970), .B1(new_n581), .B2(new_n584), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n972), .A2(new_n973), .A3(new_n600), .ZN(new_n974));
  NAND2_X1  g549(.A1(G288), .A2(KEYINPUT105), .ZN(new_n975));
  AOI21_X1  g550(.A(G290), .B1(new_n975), .B2(new_n971), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n967), .B(new_n969), .C1(new_n974), .C2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n600), .B1(new_n972), .B2(new_n973), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n975), .A2(G290), .A3(new_n971), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n978), .A2(new_n979), .A3(KEYINPUT106), .A4(new_n966), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT107), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n982), .B(KEYINPUT42), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n908), .B(new_n630), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n612), .A2(new_n566), .A3(new_n571), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT103), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n987), .B1(new_n622), .B2(new_n612), .ZN(new_n988));
  NAND3_X1  g563(.A1(G299), .A2(new_n625), .A3(KEYINPUT103), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n986), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n984), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(G299), .A2(new_n625), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n985), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT41), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT104), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT104), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n994), .A2(new_n998), .A3(new_n995), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n988), .A2(new_n989), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n986), .A2(new_n995), .ZN(new_n1001));
  AOI22_X1  g576(.A1(new_n997), .A2(new_n999), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n992), .B1(new_n1002), .B2(new_n984), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n983), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT42), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n982), .B(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n1003), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(G868), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n879), .A2(G868), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n963), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n628), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1014));
  NOR3_X1   g589(.A1(new_n1014), .A2(KEYINPUT108), .A3(new_n1011), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1013), .A2(new_n1015), .ZN(G295));
  NAND2_X1  g591(.A1(new_n1010), .A2(new_n1012), .ZN(G331));
  INV_X1    g592(.A(KEYINPUT44), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT43), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n998), .B1(new_n994), .B2(new_n995), .ZN(new_n1021));
  AOI211_X1 g596(.A(KEYINPUT104), .B(KEYINPUT41), .C1(new_n993), .C2(new_n985), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1020), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT109), .B1(new_n904), .B2(new_n907), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n530), .A2(new_n531), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT72), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(G168), .B1(new_n1028), .B2(new_n529), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1029), .B1(new_n576), .B2(G168), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n893), .B1(new_n902), .B2(new_n903), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n906), .A2(new_n879), .A3(new_n889), .A4(new_n901), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT109), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1024), .A2(new_n1030), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n574), .B1(new_n1028), .B2(new_n529), .ZN(new_n1036));
  INV_X1    g611(.A(new_n575), .ZN(new_n1037));
  OAI21_X1  g612(.A(G168), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1029), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1031), .A2(new_n1033), .A3(new_n1032), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1033), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1040), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1023), .A2(new_n1035), .A3(new_n1043), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n977), .A2(new_n980), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1024), .A2(new_n1030), .A3(new_n1034), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1030), .B1(new_n1024), .B2(new_n1034), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n991), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1044), .A2(KEYINPUT111), .A3(new_n1045), .A4(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(G37), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n990), .B1(new_n1043), .B2(new_n1035), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1052), .B1(new_n1023), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT111), .B1(new_n1054), .B2(new_n1045), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1051), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1044), .A2(new_n1048), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT110), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT110), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1054), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1058), .A2(new_n1060), .A3(new_n981), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1019), .B1(new_n1056), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1043), .A2(new_n1035), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1048), .B(new_n1045), .C1(new_n1002), .C2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT111), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1066), .A2(new_n1050), .A3(new_n1049), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT112), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n994), .B2(new_n995), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n993), .A2(KEYINPUT112), .A3(KEYINPUT41), .A4(new_n985), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1069), .B(new_n1070), .C1(new_n990), .C2(KEYINPUT41), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1048), .A2(KEYINPUT113), .B1(new_n1053), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT113), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1052), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1045), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n1067), .A2(KEYINPUT43), .A3(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1018), .B1(new_n1062), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT114), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1078), .B1(new_n1067), .B2(new_n1075), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1053), .A2(new_n1071), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(new_n1073), .B2(new_n1052), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1074), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n981), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1080), .A2(new_n1084), .A3(KEYINPUT114), .A4(new_n1066), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1079), .A2(KEYINPUT43), .A3(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1056), .A2(new_n1019), .A3(new_n1061), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT44), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1077), .B1(new_n1086), .B2(new_n1088), .ZN(G397));
  INV_X1    g664(.A(G1384), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n496), .B2(new_n502), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT45), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n471), .A2(new_n477), .A3(G40), .A4(new_n479), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n732), .B(G2067), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n717), .B(new_n721), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n841), .B(new_n845), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1095), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n1100), .A2(KEYINPUT126), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(KEYINPUT126), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1095), .A2(new_n850), .A3(new_n600), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1103), .B(KEYINPUT48), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1101), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1095), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n842), .A2(new_n844), .ZN(new_n1107));
  OR2_X1    g682(.A1(new_n1107), .A2(KEYINPUT125), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1098), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(KEYINPUT125), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(G2067), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n732), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1106), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1095), .A2(new_n721), .ZN(new_n1115));
  XOR2_X1   g690(.A(new_n1115), .B(KEYINPUT46), .Z(new_n1116));
  NAND2_X1  g691(.A1(new_n1096), .A2(new_n718), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1116), .B1(new_n1117), .B2(new_n1095), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1118), .B(KEYINPUT47), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1105), .A2(new_n1114), .A3(new_n1119), .ZN(new_n1120));
  OR2_X1    g695(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1121));
  INV_X1    g696(.A(G2078), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1094), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .A4(new_n1093), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1124), .B(KEYINPUT53), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT50), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1127), .B(new_n1090), .C1(new_n496), .C2(new_n502), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n1128), .B(KEYINPUT115), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT121), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1094), .B1(KEYINPUT50), .B2(new_n1091), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1130), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1133), .A2(G1961), .A3(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n576), .B1(new_n1126), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(KEYINPUT123), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1138), .B(new_n576), .C1(new_n1126), .C2(new_n1135), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1129), .A2(new_n769), .A3(new_n1131), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1121), .A2(new_n1123), .A3(new_n1093), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n763), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(G8), .B1(new_n1144), .B2(G286), .ZN(new_n1145));
  AOI21_X1  g720(.A(G168), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT51), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT51), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1148), .B(G8), .C1(new_n1144), .C2(G286), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(KEYINPUT62), .ZN(new_n1151));
  OR2_X1    g726(.A1(new_n1094), .A2(new_n1091), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1152), .B(G8), .C1(new_n802), .C2(G288), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT52), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT52), .ZN(new_n1155));
  XOR2_X1   g730(.A(KEYINPUT117), .B(G1976), .Z(new_n1156));
  OAI21_X1  g731(.A(new_n1155), .B1(new_n804), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1154), .B1(new_n1153), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT118), .ZN(new_n1159));
  INV_X1    g734(.A(G1981), .ZN(new_n1160));
  XNOR2_X1  g735(.A(G305), .B(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1159), .B1(new_n1161), .B2(KEYINPUT49), .ZN(new_n1162));
  XNOR2_X1  g737(.A(G305), .B(G1981), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT49), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1163), .A2(KEYINPUT118), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1152), .A2(G8), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1167), .B1(new_n1161), .B2(KEYINPUT49), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1158), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1142), .A2(new_n819), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1131), .A2(new_n1128), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1170), .B1(G2090), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(G8), .ZN(new_n1173));
  AND2_X1   g748(.A1(G303), .A2(G8), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT55), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1175), .B1(KEYINPUT116), .B2(new_n1176), .ZN(new_n1177));
  XOR2_X1   g752(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n1178));
  NAND2_X1  g753(.A1(new_n1174), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1173), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1129), .A2(new_n740), .A3(new_n1131), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1183), .A2(new_n1170), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1180), .A2(new_n1184), .A3(G8), .ZN(new_n1185));
  AND3_X1   g760(.A1(new_n1169), .A2(new_n1182), .A3(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT62), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1147), .A2(new_n1187), .A3(new_n1149), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1140), .A2(new_n1151), .A3(new_n1186), .A4(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1185), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1169), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1192));
  NOR2_X1   g767(.A1(G288), .A2(G1976), .ZN(new_n1193));
  AOI22_X1  g768(.A1(new_n1192), .A2(new_n1193), .B1(new_n1160), .B2(new_n821), .ZN(new_n1194));
  XOR2_X1   g769(.A(new_n1167), .B(KEYINPUT119), .Z(new_n1195));
  OAI21_X1  g770(.A(new_n1191), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  AND3_X1   g771(.A1(new_n1144), .A2(G8), .A3(G168), .ZN(new_n1197));
  NAND4_X1  g772(.A1(new_n1169), .A2(new_n1182), .A3(new_n1185), .A4(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT63), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  AND2_X1   g775(.A1(new_n1197), .A2(KEYINPUT63), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1184), .A2(G8), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1202), .A2(new_n1181), .ZN(new_n1203));
  NAND4_X1  g778(.A1(new_n1201), .A2(new_n1169), .A3(new_n1185), .A4(new_n1203), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1196), .B1(new_n1200), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1189), .A2(new_n1205), .ZN(new_n1206));
  XOR2_X1   g781(.A(KEYINPUT58), .B(G1341), .Z(new_n1207));
  NAND2_X1  g782(.A1(new_n1152), .A2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1208), .B1(new_n1142), .B2(G1996), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1209), .A2(new_n545), .ZN(new_n1210));
  XOR2_X1   g785(.A(new_n1210), .B(KEYINPUT59), .Z(new_n1211));
  AND3_X1   g786(.A1(new_n1121), .A2(new_n1123), .A3(new_n1093), .ZN(new_n1212));
  XNOR2_X1  g787(.A(KEYINPUT56), .B(G2072), .ZN(new_n1213));
  AOI22_X1  g788(.A1(new_n1212), .A2(new_n1213), .B1(new_n1171), .B2(new_n747), .ZN(new_n1214));
  AOI21_X1  g789(.A(KEYINPUT57), .B1(new_n617), .B2(KEYINPUT120), .ZN(new_n1215));
  XNOR2_X1  g790(.A(G299), .B(new_n1215), .ZN(new_n1216));
  OR2_X1    g791(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1219), .A2(KEYINPUT61), .ZN(new_n1220));
  INV_X1    g795(.A(KEYINPUT61), .ZN(new_n1221));
  NAND3_X1  g796(.A1(new_n1217), .A2(new_n1221), .A3(new_n1218), .ZN(new_n1222));
  AOI21_X1  g797(.A(new_n1211), .B1(new_n1220), .B2(new_n1222), .ZN(new_n1223));
  NOR3_X1   g798(.A1(new_n1133), .A2(G1348), .A3(new_n1134), .ZN(new_n1224));
  NOR2_X1   g799(.A1(new_n1152), .A2(G2067), .ZN(new_n1225));
  NOR2_X1   g800(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1226), .A2(KEYINPUT60), .ZN(new_n1227));
  INV_X1    g802(.A(KEYINPUT60), .ZN(new_n1228));
  OAI21_X1  g803(.A(new_n1228), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1229));
  NAND3_X1  g804(.A1(new_n1227), .A2(new_n625), .A3(new_n1229), .ZN(new_n1230));
  NAND3_X1  g805(.A1(new_n1226), .A2(KEYINPUT60), .A3(new_n612), .ZN(new_n1231));
  NAND3_X1  g806(.A1(new_n1223), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  NOR2_X1   g807(.A1(new_n1226), .A2(new_n612), .ZN(new_n1233));
  INV_X1    g808(.A(new_n1217), .ZN(new_n1234));
  OAI21_X1  g809(.A(new_n1218), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  INV_X1    g810(.A(KEYINPUT122), .ZN(new_n1236));
  NAND2_X1  g811(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  OAI211_X1 g812(.A(KEYINPUT122), .B(new_n1218), .C1(new_n1233), .C2(new_n1234), .ZN(new_n1238));
  NAND3_X1  g813(.A1(new_n1232), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  INV_X1    g814(.A(KEYINPUT124), .ZN(new_n1240));
  OAI21_X1  g815(.A(KEYINPUT53), .B1(new_n1142), .B2(new_n1240), .ZN(new_n1241));
  XNOR2_X1  g816(.A(new_n1241), .B(new_n1124), .ZN(new_n1242));
  OAI21_X1  g817(.A(G171), .B1(new_n1242), .B2(new_n1135), .ZN(new_n1243));
  OR3_X1    g818(.A1(new_n1133), .A2(G1961), .A3(new_n1134), .ZN(new_n1244));
  NAND3_X1  g819(.A1(new_n1244), .A2(G301), .A3(new_n1125), .ZN(new_n1245));
  NAND3_X1  g820(.A1(new_n1243), .A2(KEYINPUT54), .A3(new_n1245), .ZN(new_n1246));
  NAND3_X1  g821(.A1(new_n1246), .A2(new_n1150), .A3(new_n1186), .ZN(new_n1247));
  INV_X1    g822(.A(KEYINPUT54), .ZN(new_n1248));
  OR3_X1    g823(.A1(new_n1242), .A2(new_n1135), .A3(new_n576), .ZN(new_n1249));
  NAND3_X1  g824(.A1(new_n1249), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1250));
  AOI21_X1  g825(.A(new_n1247), .B1(new_n1248), .B2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g826(.A(new_n1206), .B1(new_n1239), .B2(new_n1251), .ZN(new_n1252));
  NOR2_X1   g827(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1253));
  XNOR2_X1  g828(.A(new_n600), .B(G1986), .ZN(new_n1254));
  AOI21_X1  g829(.A(new_n1106), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g830(.A(new_n1120), .B1(new_n1252), .B2(new_n1255), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g831(.A1(new_n1062), .A2(new_n1076), .ZN(new_n1258));
  NOR3_X1   g832(.A1(G401), .A2(new_n461), .A3(G227), .ZN(new_n1259));
  OAI21_X1  g833(.A(new_n1259), .B1(new_n706), .B2(new_n707), .ZN(new_n1260));
  INV_X1    g834(.A(KEYINPUT127), .ZN(new_n1261));
  XNOR2_X1  g835(.A(new_n1260), .B(new_n1261), .ZN(new_n1262));
  OAI21_X1  g836(.A(new_n1262), .B1(new_n950), .B2(new_n955), .ZN(new_n1263));
  NOR2_X1   g837(.A1(new_n1258), .A2(new_n1263), .ZN(G308));
  OAI221_X1 g838(.A(new_n1262), .B1(new_n950), .B2(new_n955), .C1(new_n1062), .C2(new_n1076), .ZN(G225));
endmodule


