

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791;

  XNOR2_X1 U371 ( .A(n376), .B(n537), .ZN(n469) );
  INV_X1 U372 ( .A(G953), .ZN(n494) );
  OR2_X1 U373 ( .A1(n602), .A2(n601), .ZN(n639) );
  XNOR2_X1 U374 ( .A(n406), .B(KEYINPUT104), .ZN(n681) );
  BUF_X2 U375 ( .A(n655), .Z(n656) );
  XNOR2_X2 U376 ( .A(n765), .B(n470), .ZN(n524) );
  XNOR2_X2 U377 ( .A(KEYINPUT78), .B(KEYINPUT79), .ZN(n377) );
  XNOR2_X2 U378 ( .A(n379), .B(n378), .ZN(n765) );
  XNOR2_X2 U379 ( .A(G104), .B(G101), .ZN(n379) );
  XNOR2_X2 U380 ( .A(G107), .B(G110), .ZN(n378) );
  INV_X1 U381 ( .A(n403), .ZN(n752) );
  XNOR2_X1 U382 ( .A(n727), .B(n435), .ZN(n585) );
  AND2_X1 U383 ( .A1(n428), .A2(n427), .ZN(n426) );
  INV_X1 U384 ( .A(n659), .ZN(n417) );
  AND2_X1 U385 ( .A1(n441), .A2(n440), .ZN(n439) );
  NAND2_X1 U386 ( .A1(n370), .A2(n408), .ZN(n667) );
  NAND2_X1 U387 ( .A1(n577), .A2(n576), .ZN(n406) );
  XNOR2_X1 U388 ( .A(n630), .B(n481), .ZN(n562) );
  NOR2_X1 U389 ( .A1(n426), .A2(n421), .ZN(n413) );
  NAND2_X2 U390 ( .A1(n426), .A2(n423), .ZN(n727) );
  XNOR2_X1 U391 ( .A(n674), .B(n676), .ZN(n677) );
  XNOR2_X1 U392 ( .A(n668), .B(KEYINPUT59), .ZN(n669) );
  XNOR2_X1 U393 ( .A(n471), .B(KEYINPUT4), .ZN(n482) );
  XNOR2_X1 U394 ( .A(n564), .B(n367), .ZN(n351) );
  XNOR2_X1 U395 ( .A(n564), .B(n367), .ZN(n566) );
  XNOR2_X1 U396 ( .A(n352), .B(n353), .ZN(n571) );
  NOR2_X1 U397 ( .A1(n691), .A2(G902), .ZN(n352) );
  XOR2_X1 U398 ( .A(n529), .B(G469), .Z(n353) );
  NAND2_X1 U399 ( .A1(n451), .A2(n457), .ZN(n354) );
  NAND2_X1 U400 ( .A1(n354), .A2(n355), .ZN(n661) );
  AND2_X1 U401 ( .A1(G472), .A2(n466), .ZN(n355) );
  BUF_X1 U402 ( .A(n765), .Z(n356) );
  BUF_X1 U403 ( .A(n687), .Z(n758) );
  XNOR2_X1 U404 ( .A(n779), .B(G146), .ZN(n528) );
  XNOR2_X1 U405 ( .A(n380), .B(n366), .ZN(n403) );
  NAND2_X1 U406 ( .A1(n381), .A2(n585), .ZN(n380) );
  XNOR2_X1 U407 ( .A(n593), .B(KEYINPUT105), .ZN(n381) );
  NAND2_X1 U408 ( .A1(n411), .A2(n426), .ZN(n410) );
  NOR2_X1 U409 ( .A1(n414), .A2(n413), .ZN(n412) );
  AND2_X1 U410 ( .A1(n423), .A2(KEYINPUT108), .ZN(n411) );
  OR2_X1 U411 ( .A1(n712), .A2(n359), .ZN(n604) );
  OR2_X1 U412 ( .A1(n789), .A2(n788), .ZN(n390) );
  INV_X1 U413 ( .A(KEYINPUT46), .ZN(n389) );
  INV_X1 U414 ( .A(KEYINPUT72), .ZN(n392) );
  XNOR2_X1 U415 ( .A(n484), .B(n539), .ZN(n779) );
  XNOR2_X1 U416 ( .A(n482), .B(G137), .ZN(n484) );
  XNOR2_X1 U417 ( .A(n431), .B(n430), .ZN(n534) );
  INV_X1 U418 ( .A(KEYINPUT8), .ZN(n430) );
  XOR2_X1 U419 ( .A(G131), .B(G140), .Z(n551) );
  INV_X1 U420 ( .A(KEYINPUT76), .ZN(n470) );
  XNOR2_X1 U421 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n473) );
  NAND2_X1 U422 ( .A1(n462), .A2(n461), .ZN(n460) );
  NAND2_X1 U423 ( .A1(n653), .A2(n464), .ZN(n461) );
  NAND2_X1 U424 ( .A1(n506), .A2(n463), .ZN(n462) );
  NAND2_X1 U425 ( .A1(n464), .A2(KEYINPUT2), .ZN(n463) );
  AND2_X1 U426 ( .A1(n409), .A2(KEYINPUT65), .ZN(n458) );
  AND2_X1 U427 ( .A1(n401), .A2(n399), .ZN(n398) );
  INV_X1 U428 ( .A(n612), .ZN(n434) );
  NAND2_X1 U429 ( .A1(n417), .A2(n415), .ZN(n423) );
  INV_X1 U430 ( .A(n424), .ZN(n415) );
  NAND2_X1 U431 ( .A1(G902), .A2(G472), .ZN(n427) );
  XNOR2_X1 U432 ( .A(n571), .B(n570), .ZN(n632) );
  XNOR2_X1 U433 ( .A(n377), .B(KEYINPUT16), .ZN(n376) );
  XNOR2_X1 U434 ( .A(G122), .B(G116), .ZN(n537) );
  INV_X1 U435 ( .A(n780), .ZN(n432) );
  NAND2_X1 U436 ( .A1(n455), .A2(n456), .ZN(n466) );
  XNOR2_X1 U437 ( .A(n654), .B(KEYINPUT87), .ZN(n456) );
  XNOR2_X1 U438 ( .A(n373), .B(G478), .ZN(n602) );
  NAND2_X1 U439 ( .A1(n759), .A2(n553), .ZN(n373) );
  BUF_X1 U440 ( .A(n632), .Z(n408) );
  NAND2_X1 U441 ( .A1(n734), .A2(n422), .ZN(n421) );
  INV_X1 U442 ( .A(KEYINPUT108), .ZN(n422) );
  NOR2_X1 U443 ( .A1(n421), .A2(n424), .ZN(n416) );
  INV_X1 U444 ( .A(KEYINPUT65), .ZN(n464) );
  NOR2_X1 U445 ( .A1(n600), .A2(KEYINPUT34), .ZN(n402) );
  NAND2_X1 U446 ( .A1(n420), .A2(n418), .ZN(n414) );
  NAND2_X1 U447 ( .A1(n419), .A2(KEYINPUT108), .ZN(n418) );
  NAND2_X1 U448 ( .A1(n417), .A2(n416), .ZN(n420) );
  INV_X1 U449 ( .A(n734), .ZN(n419) );
  INV_X1 U450 ( .A(KEYINPUT15), .ZN(n476) );
  NOR2_X1 U451 ( .A1(G237), .A2(G902), .ZN(n477) );
  NAND2_X1 U452 ( .A1(n425), .A2(n553), .ZN(n424) );
  INV_X1 U453 ( .A(G472), .ZN(n425) );
  XNOR2_X1 U454 ( .A(KEYINPUT5), .B(G131), .ZN(n485) );
  XOR2_X1 U455 ( .A(G101), .B(G116), .Z(n486) );
  INV_X1 U456 ( .A(KEYINPUT10), .ZN(n492) );
  INV_X1 U457 ( .A(KEYINPUT48), .ZN(n386) );
  XNOR2_X1 U458 ( .A(n390), .B(n389), .ZN(n388) );
  NAND2_X1 U459 ( .A1(n632), .A2(n596), .ZN(n593) );
  OR2_X1 U460 ( .A1(n584), .A2(n520), .ZN(n521) );
  AND2_X1 U461 ( .A1(n584), .A2(n583), .ZN(n596) );
  INV_X1 U462 ( .A(KEYINPUT6), .ZN(n435) );
  XNOR2_X1 U463 ( .A(n569), .B(n568), .ZN(n574) );
  XNOR2_X1 U464 ( .A(n567), .B(KEYINPUT66), .ZN(n568) );
  BUF_X1 U465 ( .A(n489), .Z(n405) );
  XNOR2_X1 U466 ( .A(KEYINPUT95), .B(KEYINPUT96), .ZN(n500) );
  XNOR2_X1 U467 ( .A(KEYINPUT24), .B(G140), .ZN(n501) );
  XNOR2_X1 U468 ( .A(n429), .B(n495), .ZN(n496) );
  XNOR2_X1 U469 ( .A(KEYINPUT23), .B(KEYINPUT75), .ZN(n495) );
  XNOR2_X1 U470 ( .A(G128), .B(G137), .ZN(n498) );
  XNOR2_X1 U471 ( .A(KEYINPUT100), .B(KEYINPUT99), .ZN(n544) );
  NOR2_X1 U472 ( .A1(G953), .A2(G237), .ZN(n547) );
  XNOR2_X1 U473 ( .A(n528), .B(n527), .ZN(n691) );
  XNOR2_X1 U474 ( .A(n385), .B(n384), .ZN(n673) );
  XNOR2_X1 U475 ( .A(n524), .B(n469), .ZN(n384) );
  AND2_X2 U476 ( .A1(n454), .A2(n466), .ZN(n687) );
  NAND2_X1 U477 ( .A1(n457), .A2(n451), .ZN(n454) );
  NAND2_X1 U478 ( .A1(G234), .A2(G237), .ZN(n516) );
  XNOR2_X1 U479 ( .A(n589), .B(n588), .ZN(n684) );
  NOR2_X1 U480 ( .A1(n613), .A2(n394), .ZN(n636) );
  XNOR2_X1 U481 ( .A(n396), .B(n395), .ZN(n394) );
  INV_X1 U482 ( .A(KEYINPUT81), .ZN(n395) );
  INV_X1 U483 ( .A(n596), .ZN(n720) );
  BUF_X1 U484 ( .A(n574), .Z(n581) );
  XNOR2_X1 U485 ( .A(n659), .B(n658), .ZN(n660) );
  BUF_X1 U486 ( .A(n494), .Z(n781) );
  XNOR2_X1 U487 ( .A(n374), .B(n541), .ZN(n759) );
  XNOR2_X1 U488 ( .A(n542), .B(n540), .ZN(n374) );
  AND2_X1 U489 ( .A1(n662), .A2(G953), .ZN(n763) );
  INV_X1 U490 ( .A(n466), .ZN(n718) );
  XNOR2_X1 U491 ( .A(n371), .B(n631), .ZN(n370) );
  BUF_X1 U492 ( .A(n684), .Z(n685) );
  INV_X1 U493 ( .A(n730), .ZN(n467) );
  BUF_X1 U494 ( .A(G110), .Z(n683) );
  AND2_X1 U495 ( .A1(n369), .A2(n364), .ZN(n357) );
  AND2_X1 U496 ( .A1(n652), .A2(KEYINPUT2), .ZN(n358) );
  NOR2_X1 U497 ( .A1(n600), .A2(n599), .ZN(n359) );
  XOR2_X1 U498 ( .A(G143), .B(G113), .Z(n360) );
  OR2_X1 U499 ( .A1(n480), .A2(n478), .ZN(n361) );
  AND2_X1 U500 ( .A1(n565), .A2(n583), .ZN(n362) );
  AND2_X1 U501 ( .A1(n596), .A2(n434), .ZN(n363) );
  AND2_X1 U502 ( .A1(n652), .A2(n465), .ZN(n364) );
  NOR2_X1 U503 ( .A1(n685), .A2(KEYINPUT44), .ZN(n365) );
  XOR2_X1 U504 ( .A(KEYINPUT93), .B(KEYINPUT33), .Z(n366) );
  XOR2_X1 U505 ( .A(n563), .B(KEYINPUT0), .Z(n367) );
  INV_X1 U506 ( .A(G902), .ZN(n553) );
  AND2_X1 U507 ( .A1(KEYINPUT44), .A2(KEYINPUT89), .ZN(n368) );
  NAND2_X1 U508 ( .A1(n369), .A2(n358), .ZN(n654) );
  NAND2_X1 U509 ( .A1(n369), .A2(n652), .ZN(n780) );
  XNOR2_X2 U510 ( .A(n387), .B(n386), .ZN(n369) );
  NAND2_X1 U511 ( .A1(n372), .A2(n630), .ZN(n371) );
  XNOR2_X1 U512 ( .A(n647), .B(KEYINPUT110), .ZN(n372) );
  NAND2_X1 U513 ( .A1(n562), .A2(n561), .ZN(n564) );
  XNOR2_X2 U514 ( .A(n375), .B(KEYINPUT91), .ZN(n630) );
  NAND2_X2 U515 ( .A1(n614), .A2(n734), .ZN(n375) );
  XNOR2_X1 U516 ( .A(n382), .B(G113), .ZN(n489) );
  XNOR2_X2 U517 ( .A(KEYINPUT3), .B(G119), .ZN(n382) );
  XNOR2_X2 U518 ( .A(n383), .B(n361), .ZN(n614) );
  NOR2_X2 U519 ( .A1(n673), .A2(n506), .ZN(n383) );
  XNOR2_X1 U520 ( .A(n447), .B(n449), .ZN(n385) );
  NAND2_X1 U521 ( .A1(n391), .A2(n388), .ZN(n387) );
  XNOR2_X1 U522 ( .A(n393), .B(n392), .ZN(n391) );
  NAND2_X1 U523 ( .A1(n633), .A2(n634), .ZN(n393) );
  NAND2_X1 U524 ( .A1(n531), .A2(n363), .ZN(n396) );
  NAND2_X1 U525 ( .A1(n398), .A2(n397), .ZN(n589) );
  NAND2_X1 U526 ( .A1(n752), .A2(KEYINPUT34), .ZN(n397) );
  AND2_X1 U527 ( .A1(n400), .A2(n616), .ZN(n399) );
  NAND2_X1 U528 ( .A1(n600), .A2(KEYINPUT34), .ZN(n400) );
  NAND2_X1 U529 ( .A1(n403), .A2(n402), .ZN(n401) );
  NAND2_X1 U530 ( .A1(n609), .A2(n365), .ZN(n453) );
  AND2_X1 U531 ( .A1(n562), .A2(n533), .ZN(n704) );
  NAND2_X1 U532 ( .A1(n404), .A2(n708), .ZN(n620) );
  NAND2_X1 U533 ( .A1(n619), .A2(KEYINPUT47), .ZN(n404) );
  OR2_X2 U534 ( .A1(n532), .A2(n530), .ZN(n642) );
  OR2_X2 U535 ( .A1(n688), .A2(G902), .ZN(n513) );
  NAND2_X1 U536 ( .A1(n433), .A2(n432), .ZN(n459) );
  XNOR2_X2 U537 ( .A(n629), .B(KEYINPUT107), .ZN(n647) );
  XNOR2_X1 U538 ( .A(n407), .B(n546), .ZN(n549) );
  XNOR2_X1 U539 ( .A(n543), .B(n360), .ZN(n407) );
  NAND2_X1 U540 ( .A1(n459), .A2(n458), .ZN(n457) );
  NAND2_X1 U541 ( .A1(n574), .A2(n721), .ZN(n575) );
  NAND2_X1 U542 ( .A1(n445), .A2(KEYINPUT89), .ZN(n441) );
  INV_X1 U543 ( .A(n655), .ZN(n436) );
  XNOR2_X2 U544 ( .A(n437), .B(n610), .ZN(n655) );
  INV_X1 U545 ( .A(KEYINPUT2), .ZN(n409) );
  NAND2_X1 U546 ( .A1(n412), .A2(n410), .ZN(n611) );
  NAND2_X1 U547 ( .A1(n659), .A2(G472), .ZN(n428) );
  NAND2_X1 U548 ( .A1(n534), .A2(G221), .ZN(n429) );
  NAND2_X1 U549 ( .A1(n494), .A2(G234), .ZN(n431) );
  AND2_X1 U550 ( .A1(n459), .A2(n409), .ZN(n717) );
  INV_X1 U551 ( .A(n655), .ZN(n433) );
  XNOR2_X2 U552 ( .A(n513), .B(n512), .ZN(n584) );
  INV_X1 U553 ( .A(n585), .ZN(n628) );
  NAND2_X1 U554 ( .A1(n468), .A2(n585), .ZN(n629) );
  NAND2_X1 U555 ( .A1(n450), .A2(n453), .ZN(n437) );
  NAND2_X1 U556 ( .A1(n436), .A2(n357), .ZN(n452) );
  INV_X1 U557 ( .A(n656), .ZN(n455) );
  NOR2_X1 U558 ( .A1(n656), .A2(G953), .ZN(n773) );
  NAND2_X1 U559 ( .A1(n438), .A2(n608), .ZN(n445) );
  NAND2_X1 U560 ( .A1(n592), .A2(n591), .ZN(n438) );
  NAND2_X1 U561 ( .A1(n442), .A2(n439), .ZN(n450) );
  NAND2_X1 U562 ( .A1(n446), .A2(n368), .ZN(n440) );
  NAND2_X1 U563 ( .A1(n444), .A2(n443), .ZN(n442) );
  NAND2_X1 U564 ( .A1(n446), .A2(KEYINPUT44), .ZN(n443) );
  NOR2_X1 U565 ( .A1(n445), .A2(KEYINPUT89), .ZN(n444) );
  NAND2_X1 U566 ( .A1(n609), .A2(n590), .ZN(n446) );
  XNOR2_X1 U567 ( .A(n405), .B(n469), .ZN(n764) );
  XNOR2_X1 U568 ( .A(n448), .B(n474), .ZN(n447) );
  INV_X1 U569 ( .A(n489), .ZN(n448) );
  XNOR2_X1 U570 ( .A(n482), .B(n475), .ZN(n449) );
  AND2_X2 U571 ( .A1(n452), .A2(n460), .ZN(n451) );
  XNOR2_X2 U572 ( .A(G143), .B(G128), .ZN(n483) );
  NAND2_X1 U573 ( .A1(n566), .A2(n362), .ZN(n569) );
  NOR2_X2 U574 ( .A1(n679), .A2(n763), .ZN(n680) );
  NOR2_X2 U575 ( .A1(n671), .A2(n763), .ZN(n672) );
  NOR2_X2 U576 ( .A1(n663), .A2(n763), .ZN(n665) );
  NOR2_X1 U577 ( .A1(n653), .A2(KEYINPUT65), .ZN(n465) );
  INV_X1 U578 ( .A(n351), .ZN(n600) );
  NAND2_X1 U579 ( .A1(n351), .A2(n467), .ZN(n595) );
  AND2_X1 U580 ( .A1(n709), .A2(n627), .ZN(n468) );
  INV_X1 U581 ( .A(KEYINPUT7), .ZN(n540) );
  XNOR2_X2 U582 ( .A(KEYINPUT64), .B(KEYINPUT71), .ZN(n471) );
  NAND2_X1 U583 ( .A1(n494), .A2(G224), .ZN(n472) );
  XNOR2_X1 U584 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X2 U585 ( .A(G125), .B(G146), .ZN(n493) );
  XNOR2_X1 U586 ( .A(n493), .B(n483), .ZN(n475) );
  XNOR2_X1 U587 ( .A(n476), .B(G902), .ZN(n506) );
  XNOR2_X1 U588 ( .A(n477), .B(KEYINPUT80), .ZN(n480) );
  INV_X1 U589 ( .A(G210), .ZN(n478) );
  INV_X1 U590 ( .A(G214), .ZN(n479) );
  OR2_X1 U591 ( .A1(n480), .A2(n479), .ZN(n734) );
  XOR2_X1 U592 ( .A(KEYINPUT68), .B(KEYINPUT19), .Z(n481) );
  XNOR2_X1 U593 ( .A(n483), .B(G134), .ZN(n539) );
  XNOR2_X1 U594 ( .A(n486), .B(n485), .ZN(n488) );
  NAND2_X1 U595 ( .A1(n547), .A2(G210), .ZN(n487) );
  XNOR2_X1 U596 ( .A(n488), .B(n487), .ZN(n490) );
  XNOR2_X1 U597 ( .A(n405), .B(n490), .ZN(n491) );
  XNOR2_X1 U598 ( .A(n528), .B(n491), .ZN(n659) );
  XNOR2_X1 U599 ( .A(n493), .B(n492), .ZN(n550) );
  INV_X1 U600 ( .A(n550), .ZN(n497) );
  XNOR2_X1 U601 ( .A(n497), .B(n496), .ZN(n505) );
  XNOR2_X1 U602 ( .A(n683), .B(G119), .ZN(n499) );
  XNOR2_X1 U603 ( .A(n499), .B(n498), .ZN(n503) );
  XNOR2_X1 U604 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U605 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U606 ( .A(n505), .B(n504), .ZN(n688) );
  XOR2_X1 U607 ( .A(KEYINPUT97), .B(KEYINPUT20), .Z(n508) );
  INV_X1 U608 ( .A(n506), .ZN(n653) );
  NAND2_X1 U609 ( .A1(n653), .A2(G234), .ZN(n507) );
  XNOR2_X1 U610 ( .A(n508), .B(n507), .ZN(n514) );
  AND2_X1 U611 ( .A1(n514), .A2(G217), .ZN(n511) );
  XNOR2_X1 U612 ( .A(KEYINPUT82), .B(KEYINPUT98), .ZN(n509) );
  XNOR2_X1 U613 ( .A(n509), .B(KEYINPUT25), .ZN(n510) );
  XNOR2_X1 U614 ( .A(n511), .B(n510), .ZN(n512) );
  NAND2_X1 U615 ( .A1(n514), .A2(G221), .ZN(n515) );
  XNOR2_X1 U616 ( .A(n515), .B(KEYINPUT21), .ZN(n723) );
  XNOR2_X1 U617 ( .A(n516), .B(KEYINPUT14), .ZN(n748) );
  NOR2_X1 U618 ( .A1(G900), .A2(n781), .ZN(n517) );
  NAND2_X1 U619 ( .A1(n517), .A2(G902), .ZN(n518) );
  NAND2_X1 U620 ( .A1(G952), .A2(n781), .ZN(n558) );
  NAND2_X1 U621 ( .A1(n518), .A2(n558), .ZN(n519) );
  NAND2_X1 U622 ( .A1(n748), .A2(n519), .ZN(n612) );
  OR2_X1 U623 ( .A1(n723), .A2(n612), .ZN(n520) );
  XNOR2_X1 U624 ( .A(n521), .B(KEYINPUT73), .ZN(n627) );
  NAND2_X1 U625 ( .A1(n727), .A2(n627), .ZN(n522) );
  XNOR2_X1 U626 ( .A(n522), .B(KEYINPUT28), .ZN(n532) );
  NAND2_X1 U627 ( .A1(G227), .A2(n781), .ZN(n523) );
  XNOR2_X1 U628 ( .A(n551), .B(n523), .ZN(n526) );
  BUF_X1 U629 ( .A(n524), .Z(n525) );
  XNOR2_X1 U630 ( .A(n526), .B(n525), .ZN(n527) );
  INV_X1 U631 ( .A(KEYINPUT74), .ZN(n529) );
  BUF_X1 U632 ( .A(n571), .Z(n530) );
  INV_X1 U633 ( .A(n530), .ZN(n531) );
  INV_X1 U634 ( .A(n642), .ZN(n533) );
  XOR2_X1 U635 ( .A(KEYINPUT9), .B(KEYINPUT101), .Z(n536) );
  NAND2_X1 U636 ( .A1(n534), .A2(G217), .ZN(n535) );
  XNOR2_X1 U637 ( .A(n536), .B(n535), .ZN(n542) );
  XNOR2_X1 U638 ( .A(n537), .B(G107), .ZN(n538) );
  XNOR2_X1 U639 ( .A(n539), .B(n538), .ZN(n541) );
  XOR2_X1 U640 ( .A(G122), .B(G104), .Z(n543) );
  XOR2_X1 U641 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n545) );
  XNOR2_X1 U642 ( .A(n545), .B(n544), .ZN(n546) );
  NAND2_X1 U643 ( .A1(G214), .A2(n547), .ZN(n548) );
  XNOR2_X1 U644 ( .A(n549), .B(n548), .ZN(n552) );
  XNOR2_X1 U645 ( .A(n551), .B(n550), .ZN(n778) );
  XNOR2_X1 U646 ( .A(n552), .B(n778), .ZN(n668) );
  NAND2_X1 U647 ( .A1(n668), .A2(n553), .ZN(n555) );
  XNOR2_X1 U648 ( .A(KEYINPUT13), .B(G475), .ZN(n554) );
  XNOR2_X1 U649 ( .A(n555), .B(n554), .ZN(n601) );
  INV_X1 U650 ( .A(KEYINPUT106), .ZN(n556) );
  XNOR2_X2 U651 ( .A(n639), .B(n556), .ZN(n709) );
  NAND2_X1 U652 ( .A1(n704), .A2(n709), .ZN(n557) );
  XNOR2_X1 U653 ( .A(n557), .B(G146), .ZN(G48) );
  XNOR2_X1 U654 ( .A(KEYINPUT94), .B(G898), .ZN(n770) );
  NOR2_X1 U655 ( .A1(n781), .A2(n770), .ZN(n768) );
  NAND2_X1 U656 ( .A1(n768), .A2(G902), .ZN(n559) );
  NAND2_X1 U657 ( .A1(n559), .A2(n558), .ZN(n560) );
  AND2_X1 U658 ( .A1(n560), .A2(n748), .ZN(n561) );
  INV_X1 U659 ( .A(KEYINPUT69), .ZN(n563) );
  INV_X1 U660 ( .A(n601), .ZN(n586) );
  OR2_X1 U661 ( .A1(n586), .A2(n602), .ZN(n738) );
  INV_X1 U662 ( .A(n738), .ZN(n565) );
  INV_X1 U663 ( .A(n723), .ZN(n583) );
  XNOR2_X1 U664 ( .A(KEYINPUT77), .B(KEYINPUT22), .ZN(n567) );
  NAND2_X1 U665 ( .A1(n628), .A2(n584), .ZN(n572) );
  XNOR2_X1 U666 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n570) );
  NOR2_X1 U667 ( .A1(n572), .A2(n408), .ZN(n573) );
  NAND2_X1 U668 ( .A1(n581), .A2(n573), .ZN(n606) );
  XNOR2_X1 U669 ( .A(n606), .B(G101), .ZN(G3) );
  INV_X1 U670 ( .A(n408), .ZN(n721) );
  XNOR2_X1 U671 ( .A(n575), .B(KEYINPUT103), .ZN(n577) );
  NOR2_X1 U672 ( .A1(n727), .A2(n584), .ZN(n576) );
  XNOR2_X1 U673 ( .A(n628), .B(KEYINPUT84), .ZN(n579) );
  INV_X1 U674 ( .A(n584), .ZN(n724) );
  AND2_X1 U675 ( .A1(n408), .A2(n724), .ZN(n578) );
  AND2_X1 U676 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U677 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U678 ( .A(n582), .B(KEYINPUT32), .ZN(n790) );
  AND2_X2 U679 ( .A1(n681), .A2(n790), .ZN(n609) );
  AND2_X1 U680 ( .A1(n586), .A2(n602), .ZN(n616) );
  INV_X1 U681 ( .A(KEYINPUT83), .ZN(n587) );
  XNOR2_X1 U682 ( .A(n587), .B(KEYINPUT35), .ZN(n588) );
  NAND2_X1 U683 ( .A1(n684), .A2(KEYINPUT90), .ZN(n590) );
  NAND2_X1 U684 ( .A1(n684), .A2(KEYINPUT44), .ZN(n592) );
  INV_X1 U685 ( .A(KEYINPUT90), .ZN(n591) );
  INV_X1 U686 ( .A(n593), .ZN(n594) );
  NAND2_X1 U687 ( .A1(n594), .A2(n727), .ZN(n730) );
  XNOR2_X1 U688 ( .A(n595), .B(KEYINPUT31), .ZN(n712) );
  NOR2_X1 U689 ( .A1(n530), .A2(n720), .ZN(n598) );
  INV_X1 U690 ( .A(n727), .ZN(n597) );
  NAND2_X1 U691 ( .A1(n598), .A2(n597), .ZN(n599) );
  AND2_X1 U692 ( .A1(n601), .A2(n602), .ZN(n711) );
  INV_X1 U693 ( .A(n711), .ZN(n644) );
  AND2_X1 U694 ( .A1(n644), .A2(n639), .ZN(n740) );
  INV_X1 U695 ( .A(KEYINPUT86), .ZN(n603) );
  XNOR2_X1 U696 ( .A(n740), .B(n603), .ZN(n621) );
  NAND2_X1 U697 ( .A1(n604), .A2(n621), .ZN(n605) );
  XNOR2_X1 U698 ( .A(n605), .B(KEYINPUT102), .ZN(n607) );
  AND2_X1 U699 ( .A1(n607), .A2(n606), .ZN(n608) );
  INV_X1 U700 ( .A(KEYINPUT45), .ZN(n610) );
  XNOR2_X1 U701 ( .A(KEYINPUT30), .B(n611), .ZN(n613) );
  BUF_X1 U702 ( .A(n614), .Z(n649) );
  NAND2_X1 U703 ( .A1(n636), .A2(n649), .ZN(n615) );
  XNOR2_X1 U704 ( .A(n615), .B(KEYINPUT109), .ZN(n617) );
  NAND2_X1 U705 ( .A1(n617), .A2(n616), .ZN(n708) );
  INV_X1 U706 ( .A(n740), .ZN(n618) );
  NAND2_X1 U707 ( .A1(n704), .A2(n618), .ZN(n619) );
  XNOR2_X1 U708 ( .A(n620), .B(KEYINPUT85), .ZN(n626) );
  INV_X1 U709 ( .A(n621), .ZN(n623) );
  XNOR2_X1 U710 ( .A(KEYINPUT70), .B(KEYINPUT47), .ZN(n622) );
  NOR2_X1 U711 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U712 ( .A1(n624), .A2(n704), .ZN(n625) );
  AND2_X1 U713 ( .A1(n626), .A2(n625), .ZN(n634) );
  INV_X1 U714 ( .A(KEYINPUT36), .ZN(n631) );
  XNOR2_X1 U715 ( .A(n667), .B(KEYINPUT88), .ZN(n633) );
  INV_X1 U716 ( .A(KEYINPUT38), .ZN(n635) );
  XNOR2_X1 U717 ( .A(n649), .B(n635), .ZN(n735) );
  NAND2_X1 U718 ( .A1(n636), .A2(n735), .ZN(n638) );
  INV_X1 U719 ( .A(KEYINPUT39), .ZN(n637) );
  XNOR2_X1 U720 ( .A(n638), .B(n637), .ZN(n645) );
  NOR2_X1 U721 ( .A1(n645), .A2(n639), .ZN(n640) );
  XNOR2_X1 U722 ( .A(n640), .B(KEYINPUT40), .ZN(n789) );
  NAND2_X1 U723 ( .A1(n735), .A2(n734), .ZN(n739) );
  NOR2_X1 U724 ( .A1(n738), .A2(n739), .ZN(n641) );
  XNOR2_X1 U725 ( .A(KEYINPUT41), .B(n641), .ZN(n751) );
  NOR2_X1 U726 ( .A1(n751), .A2(n642), .ZN(n643) );
  XNOR2_X1 U727 ( .A(n643), .B(KEYINPUT42), .ZN(n788) );
  OR2_X1 U728 ( .A1(n645), .A2(n644), .ZN(n714) );
  AND2_X1 U729 ( .A1(n721), .A2(n734), .ZN(n646) );
  NAND2_X1 U730 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U731 ( .A(n648), .B(KEYINPUT43), .ZN(n651) );
  INV_X1 U732 ( .A(n649), .ZN(n650) );
  NAND2_X1 U733 ( .A1(n651), .A2(n650), .ZN(n715) );
  AND2_X1 U734 ( .A1(n714), .A2(n715), .ZN(n652) );
  XNOR2_X1 U735 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n657) );
  XOR2_X1 U736 ( .A(n657), .B(KEYINPUT62), .Z(n658) );
  XNOR2_X1 U737 ( .A(n661), .B(n660), .ZN(n663) );
  INV_X1 U738 ( .A(G952), .ZN(n662) );
  XNOR2_X1 U739 ( .A(KEYINPUT113), .B(KEYINPUT63), .ZN(n664) );
  XNOR2_X1 U740 ( .A(n665), .B(n664), .ZN(G57) );
  XOR2_X1 U741 ( .A(G125), .B(KEYINPUT37), .Z(n666) );
  XNOR2_X1 U742 ( .A(n667), .B(n666), .ZN(G27) );
  NAND2_X1 U743 ( .A1(n687), .A2(G475), .ZN(n670) );
  XNOR2_X1 U744 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U745 ( .A(n672), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U746 ( .A1(n687), .A2(G210), .ZN(n678) );
  BUF_X1 U747 ( .A(n673), .Z(n674) );
  XNOR2_X1 U748 ( .A(KEYINPUT92), .B(KEYINPUT54), .ZN(n675) );
  XOR2_X1 U749 ( .A(n675), .B(KEYINPUT55), .Z(n676) );
  XNOR2_X1 U750 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U751 ( .A(n680), .B(KEYINPUT56), .ZN(G51) );
  BUF_X1 U752 ( .A(n681), .Z(n682) );
  XNOR2_X1 U753 ( .A(n682), .B(n683), .ZN(G12) );
  XNOR2_X1 U754 ( .A(G122), .B(KEYINPUT126), .ZN(n686) );
  XOR2_X1 U755 ( .A(n686), .B(n685), .Z(G24) );
  NAND2_X1 U756 ( .A1(n758), .A2(G217), .ZN(n689) );
  XNOR2_X1 U757 ( .A(n689), .B(n688), .ZN(n690) );
  NOR2_X1 U758 ( .A1(n690), .A2(n763), .ZN(G66) );
  NAND2_X1 U759 ( .A1(n758), .A2(G469), .ZN(n697) );
  XNOR2_X1 U760 ( .A(n691), .B(KEYINPUT120), .ZN(n695) );
  XOR2_X1 U761 ( .A(KEYINPUT119), .B(KEYINPUT121), .Z(n693) );
  XNOR2_X1 U762 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n692) );
  XNOR2_X1 U763 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U764 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U765 ( .A(n697), .B(n696), .ZN(n698) );
  NOR2_X1 U766 ( .A1(n698), .A2(n763), .ZN(G54) );
  NAND2_X1 U767 ( .A1(n359), .A2(n709), .ZN(n699) );
  XNOR2_X1 U768 ( .A(n699), .B(G104), .ZN(G6) );
  XNOR2_X1 U769 ( .A(G107), .B(KEYINPUT27), .ZN(n703) );
  XOR2_X1 U770 ( .A(KEYINPUT114), .B(KEYINPUT26), .Z(n701) );
  NAND2_X1 U771 ( .A1(n359), .A2(n711), .ZN(n700) );
  XNOR2_X1 U772 ( .A(n701), .B(n700), .ZN(n702) );
  XNOR2_X1 U773 ( .A(n703), .B(n702), .ZN(G9) );
  NAND2_X1 U774 ( .A1(n704), .A2(n711), .ZN(n706) );
  XOR2_X1 U775 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n705) );
  XNOR2_X1 U776 ( .A(n706), .B(n705), .ZN(n707) );
  XOR2_X1 U777 ( .A(G128), .B(n707), .Z(G30) );
  XNOR2_X1 U778 ( .A(n708), .B(G143), .ZN(G45) );
  NAND2_X1 U779 ( .A1(n709), .A2(n712), .ZN(n710) );
  XNOR2_X1 U780 ( .A(n710), .B(G113), .ZN(G15) );
  NAND2_X1 U781 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U782 ( .A(n713), .B(G116), .ZN(G18) );
  XNOR2_X1 U783 ( .A(G134), .B(n714), .ZN(G36) );
  XNOR2_X1 U784 ( .A(n715), .B(G140), .ZN(n716) );
  XNOR2_X1 U785 ( .A(KEYINPUT116), .B(n716), .ZN(G42) );
  NOR2_X1 U786 ( .A1(n717), .A2(n718), .ZN(n719) );
  NOR2_X1 U787 ( .A1(n719), .A2(G953), .ZN(n756) );
  NAND2_X1 U788 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U789 ( .A(n722), .B(KEYINPUT50), .ZN(n729) );
  NAND2_X1 U790 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U791 ( .A(KEYINPUT49), .B(n725), .ZN(n726) );
  NOR2_X1 U792 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U793 ( .A1(n729), .A2(n728), .ZN(n731) );
  NAND2_X1 U794 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U795 ( .A(KEYINPUT51), .B(n732), .ZN(n733) );
  NOR2_X1 U796 ( .A1(n733), .A2(n751), .ZN(n745) );
  NOR2_X1 U797 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U798 ( .A(KEYINPUT117), .B(n736), .Z(n737) );
  NOR2_X1 U799 ( .A1(n738), .A2(n737), .ZN(n742) );
  NOR2_X1 U800 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U801 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U802 ( .A1(n752), .A2(n743), .ZN(n744) );
  NOR2_X1 U803 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U804 ( .A(n746), .B(KEYINPUT118), .ZN(n747) );
  XNOR2_X1 U805 ( .A(n747), .B(KEYINPUT52), .ZN(n750) );
  NAND2_X1 U806 ( .A1(n748), .A2(G952), .ZN(n749) );
  NOR2_X1 U807 ( .A1(n750), .A2(n749), .ZN(n754) );
  NOR2_X1 U808 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U809 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U810 ( .A1(n756), .A2(n755), .ZN(n757) );
  XOR2_X1 U811 ( .A(KEYINPUT53), .B(n757), .Z(G75) );
  NAND2_X1 U812 ( .A1(n758), .A2(G478), .ZN(n761) );
  XOR2_X1 U813 ( .A(n759), .B(KEYINPUT122), .Z(n760) );
  XNOR2_X1 U814 ( .A(n761), .B(n760), .ZN(n762) );
  NOR2_X1 U815 ( .A1(n763), .A2(n762), .ZN(G63) );
  XNOR2_X1 U816 ( .A(n356), .B(KEYINPUT125), .ZN(n766) );
  XNOR2_X1 U817 ( .A(n764), .B(n766), .ZN(n767) );
  NOR2_X1 U818 ( .A1(n768), .A2(n767), .ZN(n777) );
  NAND2_X1 U819 ( .A1(G953), .A2(G224), .ZN(n769) );
  XNOR2_X1 U820 ( .A(n769), .B(KEYINPUT61), .ZN(n771) );
  NAND2_X1 U821 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U822 ( .A(KEYINPUT123), .B(n772), .ZN(n775) );
  XNOR2_X1 U823 ( .A(n773), .B(KEYINPUT124), .ZN(n774) );
  NOR2_X1 U824 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U825 ( .A(n777), .B(n776), .Z(G69) );
  XNOR2_X1 U826 ( .A(n779), .B(n778), .ZN(n783) );
  XNOR2_X1 U827 ( .A(n780), .B(n783), .ZN(n782) );
  NAND2_X1 U828 ( .A1(n782), .A2(n781), .ZN(n787) );
  XNOR2_X1 U829 ( .A(G227), .B(n783), .ZN(n784) );
  NAND2_X1 U830 ( .A1(n784), .A2(G900), .ZN(n785) );
  NAND2_X1 U831 ( .A1(n785), .A2(G953), .ZN(n786) );
  NAND2_X1 U832 ( .A1(n787), .A2(n786), .ZN(G72) );
  XOR2_X1 U833 ( .A(G137), .B(n788), .Z(G39) );
  XOR2_X1 U834 ( .A(G131), .B(n789), .Z(G33) );
  XOR2_X1 U835 ( .A(G119), .B(n790), .Z(n791) );
  XNOR2_X1 U836 ( .A(KEYINPUT127), .B(n791), .ZN(G21) );
endmodule

