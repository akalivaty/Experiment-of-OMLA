

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738;

  XNOR2_X1 U369 ( .A(n605), .B(n411), .ZN(n723) );
  NAND2_X1 U370 ( .A1(n387), .A2(n386), .ZN(n533) );
  XNOR2_X2 U371 ( .A(n506), .B(n449), .ZN(n380) );
  INV_X1 U372 ( .A(G953), .ZN(n725) );
  NOR2_X1 U373 ( .A1(n731), .A2(n733), .ZN(n532) );
  AND2_X2 U374 ( .A1(n712), .A2(n448), .ZN(n391) );
  NOR2_X1 U375 ( .A1(n657), .A2(n656), .ZN(n539) );
  OR2_X1 U376 ( .A1(n401), .A2(n399), .ZN(n398) );
  XNOR2_X1 U377 ( .A(n562), .B(KEYINPUT107), .ZN(n732) );
  XNOR2_X1 U378 ( .A(n463), .B(KEYINPUT19), .ZN(n575) );
  XNOR2_X1 U379 ( .A(n422), .B(KEYINPUT101), .ZN(n631) );
  NOR2_X1 U380 ( .A1(n569), .A2(n568), .ZN(n588) );
  OR2_X1 U381 ( .A1(n542), .A2(n384), .ZN(n550) );
  XNOR2_X2 U382 ( .A(n390), .B(n347), .ZN(n601) );
  XNOR2_X1 U383 ( .A(n578), .B(n394), .ZN(n393) );
  INV_X1 U384 ( .A(KEYINPUT82), .ZN(n394) );
  XNOR2_X1 U385 ( .A(n475), .B(n407), .ZN(n717) );
  INV_X1 U386 ( .A(n491), .ZN(n407) );
  NAND2_X1 U387 ( .A1(n396), .A2(n412), .ZN(n605) );
  AND2_X1 U388 ( .A1(n729), .A2(n596), .ZN(n412) );
  OR2_X1 U389 ( .A1(G902), .A2(G237), .ZN(n462) );
  XNOR2_X1 U390 ( .A(n380), .B(n472), .ZN(n475) );
  XNOR2_X1 U391 ( .A(G131), .B(G134), .ZN(n472) );
  XNOR2_X1 U392 ( .A(n409), .B(G146), .ZN(n460) );
  INV_X1 U393 ( .A(G125), .ZN(n409) );
  OR2_X1 U394 ( .A1(n413), .A2(n397), .ZN(n364) );
  INV_X1 U395 ( .A(KEYINPUT87), .ZN(n377) );
  XOR2_X1 U396 ( .A(G140), .B(G137), .Z(n491) );
  XNOR2_X1 U397 ( .A(n460), .B(KEYINPUT10), .ZN(n485) );
  XNOR2_X1 U398 ( .A(G146), .B(G107), .ZN(n477) );
  INV_X1 U399 ( .A(KEYINPUT79), .ZN(n476) );
  XNOR2_X1 U400 ( .A(KEYINPUT6), .B(n542), .ZN(n589) );
  AND2_X1 U401 ( .A1(n521), .A2(n653), .ZN(n426) );
  INV_X1 U402 ( .A(KEYINPUT0), .ZN(n382) );
  NAND2_X1 U403 ( .A1(n575), .A2(n464), .ZN(n383) );
  INV_X1 U404 ( .A(KEYINPUT84), .ZN(n411) );
  XNOR2_X1 U405 ( .A(G119), .B(KEYINPUT93), .ZN(n488) );
  XNOR2_X1 U406 ( .A(n416), .B(n491), .ZN(n415) );
  XNOR2_X1 U407 ( .A(n492), .B(n486), .ZN(n416) );
  XNOR2_X1 U408 ( .A(G128), .B(G110), .ZN(n492) );
  XNOR2_X1 U409 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n486) );
  INV_X1 U410 ( .A(n485), .ZN(n718) );
  INV_X1 U411 ( .A(KEYINPUT97), .ZN(n510) );
  XNOR2_X1 U412 ( .A(KEYINPUT98), .B(KEYINPUT100), .ZN(n503) );
  XOR2_X1 U413 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n504) );
  INV_X1 U414 ( .A(KEYINPUT41), .ZN(n388) );
  INV_X1 U415 ( .A(KEYINPUT39), .ZN(n583) );
  NOR2_X1 U416 ( .A1(n582), .A2(n581), .ZN(n584) );
  INV_X1 U417 ( .A(n590), .ZN(n400) );
  NAND2_X1 U418 ( .A1(G214), .A2(n462), .ZN(n642) );
  XNOR2_X1 U419 ( .A(n359), .B(KEYINPUT104), .ZN(n401) );
  NAND2_X1 U420 ( .A1(n589), .A2(n360), .ZN(n359) );
  NOR2_X1 U421 ( .A1(n631), .A2(n361), .ZN(n360) );
  INV_X1 U422 ( .A(n588), .ZN(n361) );
  XNOR2_X1 U423 ( .A(n516), .B(n515), .ZN(n537) );
  INV_X1 U424 ( .A(G478), .ZN(n515) );
  XNOR2_X1 U425 ( .A(n502), .B(n423), .ZN(n538) );
  XNOR2_X1 U426 ( .A(n501), .B(n424), .ZN(n423) );
  INV_X1 U427 ( .A(G475), .ZN(n424) );
  INV_X1 U428 ( .A(n542), .ZN(n660) );
  OR2_X1 U429 ( .A1(n689), .A2(G902), .ZN(n379) );
  XNOR2_X1 U430 ( .A(n495), .B(n410), .ZN(n569) );
  XNOR2_X1 U431 ( .A(n494), .B(KEYINPUT25), .ZN(n410) );
  XNOR2_X1 U432 ( .A(n474), .B(n362), .ZN(n613) );
  XNOR2_X1 U433 ( .A(n475), .B(n473), .ZN(n362) );
  XOR2_X1 U434 ( .A(KEYINPUT88), .B(n609), .Z(n702) );
  AND2_X1 U435 ( .A1(n357), .A2(n350), .ZN(n678) );
  NAND2_X1 U436 ( .A1(n358), .A2(n349), .ZN(n357) );
  NOR2_X1 U437 ( .A1(n732), .A2(n564), .ZN(n566) );
  NOR2_X2 U438 ( .A1(n633), .A2(n635), .ZN(n648) );
  AND2_X1 U439 ( .A1(n371), .A2(n369), .ZN(n368) );
  NAND2_X1 U440 ( .A1(n370), .A2(n397), .ZN(n369) );
  NOR2_X1 U441 ( .A1(G953), .A2(G237), .ZN(n465) );
  INV_X1 U442 ( .A(KEYINPUT44), .ZN(n376) );
  XNOR2_X1 U443 ( .A(G140), .B(G122), .ZN(n437) );
  INV_X1 U444 ( .A(G131), .ZN(n420) );
  XOR2_X1 U445 ( .A(KEYINPUT12), .B(KEYINPUT95), .Z(n433) );
  INV_X1 U446 ( .A(KEYINPUT4), .ZN(n449) );
  XOR2_X1 U447 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n459) );
  NAND2_X1 U448 ( .A1(n538), .A2(n520), .ZN(n646) );
  NAND2_X1 U449 ( .A1(n588), .A2(n660), .ZN(n571) );
  XOR2_X1 U450 ( .A(G137), .B(KEYINPUT5), .Z(n467) );
  XNOR2_X1 U451 ( .A(n458), .B(n457), .ZN(n704) );
  XNOR2_X1 U452 ( .A(n421), .B(n418), .ZN(n500) );
  XNOR2_X1 U453 ( .A(n438), .B(n419), .ZN(n418) );
  XNOR2_X1 U454 ( .A(n436), .B(n485), .ZN(n421) );
  XNOR2_X1 U455 ( .A(n437), .B(n420), .ZN(n419) );
  XNOR2_X1 U456 ( .A(n717), .B(n406), .ZN(n689) );
  XNOR2_X1 U457 ( .A(n481), .B(n478), .ZN(n406) );
  XNOR2_X1 U458 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U459 ( .A(n428), .B(n704), .ZN(n683) );
  XNOR2_X1 U460 ( .A(n430), .B(n429), .ZN(n428) );
  XNOR2_X1 U461 ( .A(n480), .B(n461), .ZN(n429) );
  XNOR2_X1 U462 ( .A(n380), .B(n348), .ZN(n430) );
  NAND2_X1 U463 ( .A1(n673), .A2(n604), .ZN(n358) );
  OR2_X1 U464 ( .A1(n401), .A2(n384), .ZN(n597) );
  AND2_X1 U465 ( .A1(n559), .A2(n569), .ZN(n395) );
  NAND2_X1 U466 ( .A1(n601), .A2(n642), .ZN(n463) );
  XNOR2_X1 U467 ( .A(n522), .B(KEYINPUT73), .ZN(n523) );
  INV_X1 U468 ( .A(G472), .ZN(n402) );
  OR2_X1 U469 ( .A1(n613), .A2(G902), .ZN(n403) );
  XNOR2_X1 U470 ( .A(G110), .B(G104), .ZN(n706) );
  XNOR2_X1 U471 ( .A(n417), .B(n414), .ZN(n699) );
  XNOR2_X1 U472 ( .A(n490), .B(n431), .ZN(n417) );
  XNOR2_X1 U473 ( .A(n718), .B(n415), .ZN(n414) );
  XNOR2_X1 U474 ( .A(n513), .B(n385), .ZN(n696) );
  XNOR2_X1 U475 ( .A(n512), .B(n351), .ZN(n385) );
  XNOR2_X1 U476 ( .A(n580), .B(KEYINPUT42), .ZN(n736) );
  NAND2_X1 U477 ( .A1(n400), .A2(n642), .ZN(n399) );
  XNOR2_X1 U478 ( .A(n519), .B(n518), .ZN(n734) );
  XNOR2_X1 U479 ( .A(KEYINPUT80), .B(KEYINPUT35), .ZN(n518) );
  XOR2_X1 U480 ( .A(KEYINPUT102), .B(n529), .Z(n530) );
  NOR2_X1 U481 ( .A1(n538), .A2(n537), .ZN(n422) );
  AND2_X1 U482 ( .A1(n392), .A2(n657), .ZN(n534) );
  XOR2_X1 U483 ( .A(n613), .B(KEYINPUT62), .Z(n615) );
  NOR2_X1 U484 ( .A1(G953), .A2(n679), .ZN(n681) );
  AND2_X1 U485 ( .A1(G210), .A2(n462), .ZN(n347) );
  XOR2_X1 U486 ( .A(n460), .B(n459), .Z(n348) );
  NAND2_X1 U487 ( .A1(n712), .A2(n606), .ZN(n349) );
  OR2_X1 U488 ( .A1(n672), .A2(n671), .ZN(n350) );
  AND2_X1 U489 ( .A1(n514), .A2(G217), .ZN(n351) );
  AND2_X1 U490 ( .A1(n349), .A2(G475), .ZN(n352) );
  XOR2_X1 U491 ( .A(KEYINPUT1), .B(KEYINPUT66), .Z(n353) );
  INV_X1 U492 ( .A(n642), .ZN(n384) );
  XOR2_X1 U493 ( .A(n439), .B(KEYINPUT67), .Z(n354) );
  XOR2_X1 U494 ( .A(G902), .B(KEYINPUT15), .Z(n448) );
  INV_X1 U495 ( .A(KEYINPUT48), .ZN(n397) );
  XNOR2_X1 U496 ( .A(n355), .B(n376), .ZN(n378) );
  NAND2_X1 U497 ( .A1(n374), .A2(n375), .ZN(n355) );
  XNOR2_X1 U498 ( .A(n356), .B(KEYINPUT121), .ZN(G66) );
  NAND2_X1 U499 ( .A1(n703), .A2(n702), .ZN(n356) );
  NOR2_X1 U500 ( .A1(n638), .A2(n413), .ZN(n373) );
  AND2_X1 U501 ( .A1(n363), .A2(n372), .ZN(n367) );
  XNOR2_X1 U502 ( .A(n586), .B(n587), .ZN(n372) );
  NOR2_X1 U503 ( .A1(n638), .A2(n364), .ZN(n363) );
  NAND2_X1 U504 ( .A1(n365), .A2(n397), .ZN(n371) );
  INV_X1 U505 ( .A(n393), .ZN(n365) );
  NAND2_X1 U506 ( .A1(n368), .A2(n366), .ZN(n396) );
  NAND2_X1 U507 ( .A1(n393), .A2(n367), .ZN(n366) );
  NAND2_X1 U508 ( .A1(n373), .A2(n372), .ZN(n370) );
  XNOR2_X1 U509 ( .A(n532), .B(n377), .ZN(n374) );
  INV_X1 U510 ( .A(n734), .ZN(n375) );
  NAND2_X1 U511 ( .A1(n548), .A2(n378), .ZN(n549) );
  XNOR2_X2 U512 ( .A(n379), .B(G469), .ZN(n572) );
  AND2_X4 U513 ( .A1(n425), .A2(n349), .ZN(n381) );
  NAND2_X1 U514 ( .A1(n425), .A2(n352), .ZN(n607) );
  NAND2_X1 U515 ( .A1(n381), .A2(G217), .ZN(n701) );
  NAND2_X1 U516 ( .A1(n381), .A2(G210), .ZN(n685) );
  NAND2_X1 U517 ( .A1(n381), .A2(G472), .ZN(n614) );
  NAND2_X1 U518 ( .A1(n381), .A2(G469), .ZN(n692) );
  NAND2_X1 U519 ( .A1(n381), .A2(G478), .ZN(n695) );
  INV_X1 U520 ( .A(n427), .ZN(n541) );
  XNOR2_X2 U521 ( .A(n383), .B(n382), .ZN(n427) );
  XNOR2_X1 U522 ( .A(n614), .B(n615), .ZN(n616) );
  INV_X1 U523 ( .A(n589), .ZN(n386) );
  XNOR2_X1 U524 ( .A(n531), .B(KEYINPUT32), .ZN(n731) );
  NAND2_X1 U525 ( .A1(n552), .A2(n395), .ZN(n582) );
  NOR2_X1 U526 ( .A1(n533), .A2(n530), .ZN(n531) );
  INV_X1 U527 ( .A(n528), .ZN(n387) );
  XNOR2_X1 U528 ( .A(n389), .B(n388), .ZN(n652) );
  NOR2_X1 U529 ( .A1(n647), .A2(n646), .ZN(n389) );
  NAND2_X1 U530 ( .A1(n683), .A2(n603), .ZN(n390) );
  NAND2_X1 U531 ( .A1(n391), .A2(n723), .ZN(n405) );
  XNOR2_X1 U532 ( .A(n533), .B(KEYINPUT85), .ZN(n392) );
  XNOR2_X1 U533 ( .A(n398), .B(KEYINPUT36), .ZN(n591) );
  XNOR2_X2 U534 ( .A(n403), .B(n402), .ZN(n542) );
  XNOR2_X2 U535 ( .A(n404), .B(G143), .ZN(n506) );
  XNOR2_X2 U536 ( .A(G128), .B(KEYINPUT65), .ZN(n404) );
  NAND2_X2 U537 ( .A1(n405), .A2(n354), .ZN(n425) );
  INV_X1 U538 ( .A(n572), .ZN(n545) );
  NAND2_X1 U539 ( .A1(n539), .A2(n589), .ZN(n497) );
  XNOR2_X2 U540 ( .A(n572), .B(n353), .ZN(n657) );
  NAND2_X1 U541 ( .A1(n408), .A2(n652), .ZN(n580) );
  NAND2_X1 U542 ( .A1(n408), .A2(n575), .ZN(n630) );
  XNOR2_X1 U543 ( .A(n574), .B(KEYINPUT109), .ZN(n408) );
  NAND2_X1 U544 ( .A1(n723), .A2(n712), .ZN(n673) );
  XNOR2_X1 U545 ( .A(n594), .B(KEYINPUT76), .ZN(n413) );
  NAND2_X1 U546 ( .A1(n427), .A2(n426), .ZN(n524) );
  XOR2_X1 U547 ( .A(n489), .B(n488), .Z(n431) );
  INV_X1 U548 ( .A(KEYINPUT81), .ZN(n565) );
  INV_X1 U549 ( .A(n640), .ZN(n596) );
  INV_X1 U550 ( .A(n567), .ZN(n558) );
  XNOR2_X1 U551 ( .A(n509), .B(n456), .ZN(n457) );
  XNOR2_X1 U552 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U553 ( .A(n511), .B(n510), .ZN(n512) );
  NOR2_X1 U554 ( .A1(n541), .A2(n675), .ZN(n499) );
  XNOR2_X1 U555 ( .A(n585), .B(KEYINPUT40), .ZN(n737) );
  INV_X1 U556 ( .A(KEYINPUT60), .ZN(n611) );
  XNOR2_X1 U557 ( .A(G113), .B(G104), .ZN(n432) );
  XNOR2_X1 U558 ( .A(n433), .B(n432), .ZN(n438) );
  XOR2_X1 U559 ( .A(G143), .B(KEYINPUT11), .Z(n435) );
  NAND2_X1 U560 ( .A1(n465), .A2(G214), .ZN(n434) );
  XNOR2_X1 U561 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U562 ( .A(n500), .B(KEYINPUT59), .ZN(n608) );
  NAND2_X1 U563 ( .A1(n448), .A2(KEYINPUT2), .ZN(n439) );
  NAND2_X1 U564 ( .A1(G237), .A2(G234), .ZN(n440) );
  XNOR2_X1 U565 ( .A(n440), .B(KEYINPUT14), .ZN(n442) );
  NAND2_X1 U566 ( .A1(G952), .A2(n442), .ZN(n672) );
  NOR2_X1 U567 ( .A1(n672), .A2(G953), .ZN(n441) );
  XNOR2_X1 U568 ( .A(n441), .B(KEYINPUT89), .ZN(n555) );
  INV_X1 U569 ( .A(n555), .ZN(n446) );
  NAND2_X1 U570 ( .A1(G902), .A2(n442), .ZN(n553) );
  INV_X1 U571 ( .A(n553), .ZN(n443) );
  NOR2_X1 U572 ( .A1(G898), .A2(n725), .ZN(n707) );
  NAND2_X1 U573 ( .A1(n443), .A2(n707), .ZN(n444) );
  XOR2_X1 U574 ( .A(KEYINPUT90), .B(n444), .Z(n445) );
  NOR2_X1 U575 ( .A1(n446), .A2(n445), .ZN(n447) );
  XNOR2_X1 U576 ( .A(KEYINPUT91), .B(n447), .ZN(n464) );
  INV_X1 U577 ( .A(n448), .ZN(n603) );
  XNOR2_X1 U578 ( .A(G119), .B(G113), .ZN(n455) );
  INV_X1 U579 ( .A(G116), .ZN(n450) );
  NAND2_X1 U580 ( .A1(n450), .A2(KEYINPUT3), .ZN(n453) );
  INV_X1 U581 ( .A(KEYINPUT3), .ZN(n451) );
  NAND2_X1 U582 ( .A1(n451), .A2(G116), .ZN(n452) );
  NAND2_X1 U583 ( .A1(n453), .A2(n452), .ZN(n454) );
  XNOR2_X1 U584 ( .A(n455), .B(n454), .ZN(n473) );
  XNOR2_X1 U585 ( .A(n473), .B(KEYINPUT74), .ZN(n458) );
  XOR2_X1 U586 ( .A(G122), .B(G107), .Z(n509) );
  XNOR2_X1 U587 ( .A(KEYINPUT75), .B(KEYINPUT16), .ZN(n456) );
  XOR2_X1 U588 ( .A(KEYINPUT68), .B(G101), .Z(n468) );
  XNOR2_X1 U589 ( .A(n468), .B(n706), .ZN(n480) );
  NAND2_X1 U590 ( .A1(G224), .A2(n725), .ZN(n461) );
  NAND2_X1 U591 ( .A1(n465), .A2(G210), .ZN(n466) );
  XNOR2_X1 U592 ( .A(n467), .B(n466), .ZN(n471) );
  XNOR2_X1 U593 ( .A(G146), .B(n468), .ZN(n469) );
  XNOR2_X1 U594 ( .A(n469), .B(KEYINPUT78), .ZN(n470) );
  XOR2_X1 U595 ( .A(n471), .B(n470), .Z(n474) );
  NAND2_X1 U596 ( .A1(G227), .A2(n725), .ZN(n479) );
  XOR2_X1 U597 ( .A(KEYINPUT94), .B(KEYINPUT21), .Z(n484) );
  NAND2_X1 U598 ( .A1(n603), .A2(G234), .ZN(n482) );
  XNOR2_X1 U599 ( .A(n482), .B(KEYINPUT20), .ZN(n493) );
  NAND2_X1 U600 ( .A1(n493), .A2(G221), .ZN(n483) );
  XNOR2_X1 U601 ( .A(n484), .B(n483), .ZN(n653) );
  NAND2_X1 U602 ( .A1(G234), .A2(n725), .ZN(n487) );
  XOR2_X1 U603 ( .A(KEYINPUT8), .B(n487), .Z(n514) );
  NAND2_X1 U604 ( .A1(G221), .A2(n514), .ZN(n490) );
  XOR2_X1 U605 ( .A(KEYINPUT70), .B(KEYINPUT92), .Z(n489) );
  NOR2_X1 U606 ( .A1(n699), .A2(G902), .ZN(n495) );
  NAND2_X1 U607 ( .A1(n493), .A2(G217), .ZN(n494) );
  NAND2_X1 U608 ( .A1(n653), .A2(n569), .ZN(n656) );
  XNOR2_X1 U609 ( .A(KEYINPUT33), .B(KEYINPUT71), .ZN(n496) );
  XNOR2_X1 U610 ( .A(n497), .B(n496), .ZN(n675) );
  XNOR2_X1 U611 ( .A(KEYINPUT72), .B(KEYINPUT34), .ZN(n498) );
  XNOR2_X1 U612 ( .A(n499), .B(n498), .ZN(n517) );
  NOR2_X1 U613 ( .A1(G902), .A2(n500), .ZN(n502) );
  XNOR2_X1 U614 ( .A(KEYINPUT13), .B(KEYINPUT96), .ZN(n501) );
  XNOR2_X1 U615 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U616 ( .A(n505), .B(G134), .Z(n508) );
  XNOR2_X1 U617 ( .A(n506), .B(G116), .ZN(n507) );
  XNOR2_X1 U618 ( .A(n508), .B(n507), .ZN(n513) );
  XNOR2_X1 U619 ( .A(n509), .B(KEYINPUT99), .ZN(n511) );
  NOR2_X1 U620 ( .A1(G902), .A2(n696), .ZN(n516) );
  INV_X1 U621 ( .A(n537), .ZN(n520) );
  NOR2_X1 U622 ( .A1(n538), .A2(n520), .ZN(n561) );
  NAND2_X1 U623 ( .A1(n517), .A2(n561), .ZN(n519) );
  INV_X1 U624 ( .A(n646), .ZN(n521) );
  INV_X1 U625 ( .A(KEYINPUT22), .ZN(n522) );
  XNOR2_X1 U626 ( .A(n524), .B(n523), .ZN(n528) );
  NOR2_X1 U627 ( .A1(n528), .A2(n569), .ZN(n526) );
  INV_X1 U628 ( .A(n657), .ZN(n598) );
  NOR2_X1 U629 ( .A1(n598), .A2(n660), .ZN(n525) );
  NAND2_X1 U630 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U631 ( .A(KEYINPUT103), .B(n527), .ZN(n733) );
  NOR2_X1 U632 ( .A1(n657), .A2(n569), .ZN(n529) );
  INV_X1 U633 ( .A(n569), .ZN(n536) );
  XOR2_X1 U634 ( .A(KEYINPUT86), .B(n534), .Z(n535) );
  NOR2_X1 U635 ( .A1(n536), .A2(n535), .ZN(n618) );
  INV_X1 U636 ( .A(n631), .ZN(n633) );
  NAND2_X1 U637 ( .A1(n538), .A2(n537), .ZN(n626) );
  INV_X1 U638 ( .A(n626), .ZN(n635) );
  NAND2_X1 U639 ( .A1(n660), .A2(n539), .ZN(n663) );
  NOR2_X1 U640 ( .A1(n541), .A2(n663), .ZN(n540) );
  XOR2_X1 U641 ( .A(KEYINPUT31), .B(n540), .Z(n636) );
  NOR2_X1 U642 ( .A1(n541), .A2(n656), .ZN(n543) );
  NAND2_X1 U643 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X1 U644 ( .A1(n545), .A2(n544), .ZN(n623) );
  NOR2_X1 U645 ( .A1(n636), .A2(n623), .ZN(n546) );
  NOR2_X1 U646 ( .A1(n648), .A2(n546), .ZN(n547) );
  NOR2_X1 U647 ( .A1(n618), .A2(n547), .ZN(n548) );
  XNOR2_X2 U648 ( .A(n549), .B(KEYINPUT45), .ZN(n712) );
  INV_X1 U649 ( .A(n601), .ZN(n590) );
  XOR2_X1 U650 ( .A(KEYINPUT30), .B(KEYINPUT106), .Z(n551) );
  XNOR2_X1 U651 ( .A(n551), .B(n550), .ZN(n552) );
  NOR2_X1 U652 ( .A1(G900), .A2(n553), .ZN(n554) );
  NAND2_X1 U653 ( .A1(n554), .A2(G953), .ZN(n556) );
  NAND2_X1 U654 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U655 ( .A1(n557), .A2(n653), .ZN(n567) );
  AND2_X1 U656 ( .A1(n572), .A2(n558), .ZN(n559) );
  NOR2_X1 U657 ( .A1(n590), .A2(n582), .ZN(n560) );
  NAND2_X1 U658 ( .A1(n561), .A2(n560), .ZN(n562) );
  NAND2_X1 U659 ( .A1(KEYINPUT47), .A2(n648), .ZN(n563) );
  XNOR2_X1 U660 ( .A(KEYINPUT83), .B(n563), .ZN(n564) );
  XNOR2_X1 U661 ( .A(n566), .B(n565), .ZN(n577) );
  XOR2_X1 U662 ( .A(KEYINPUT69), .B(n567), .Z(n568) );
  XOR2_X1 U663 ( .A(KEYINPUT28), .B(KEYINPUT108), .Z(n570) );
  XNOR2_X1 U664 ( .A(n571), .B(n570), .ZN(n573) );
  NAND2_X1 U665 ( .A1(n573), .A2(n572), .ZN(n574) );
  NAND2_X1 U666 ( .A1(n630), .A2(KEYINPUT47), .ZN(n576) );
  NAND2_X1 U667 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U668 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n587) );
  INV_X1 U669 ( .A(KEYINPUT38), .ZN(n579) );
  XNOR2_X1 U670 ( .A(n400), .B(n579), .ZN(n643) );
  NAND2_X1 U671 ( .A1(n643), .A2(n642), .ZN(n647) );
  INV_X1 U672 ( .A(n643), .ZN(n581) );
  XNOR2_X1 U673 ( .A(n584), .B(n583), .ZN(n595) );
  NAND2_X1 U674 ( .A1(n595), .A2(n633), .ZN(n585) );
  NAND2_X1 U675 ( .A1(n736), .A2(n737), .ZN(n586) );
  NOR2_X1 U676 ( .A1(n657), .A2(n591), .ZN(n638) );
  NOR2_X1 U677 ( .A1(KEYINPUT47), .A2(n648), .ZN(n592) );
  XNOR2_X1 U678 ( .A(KEYINPUT77), .B(n592), .ZN(n593) );
  NOR2_X1 U679 ( .A1(n630), .A2(n593), .ZN(n594) );
  AND2_X1 U680 ( .A1(n595), .A2(n635), .ZN(n640) );
  NOR2_X1 U681 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U682 ( .A(n599), .B(KEYINPUT43), .ZN(n600) );
  NOR2_X1 U683 ( .A1(n400), .A2(n600), .ZN(n602) );
  XNOR2_X1 U684 ( .A(KEYINPUT105), .B(n602), .ZN(n729) );
  INV_X1 U685 ( .A(KEYINPUT2), .ZN(n604) );
  NOR2_X1 U686 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U687 ( .A(n608), .B(n607), .ZN(n610) );
  NOR2_X1 U688 ( .A1(G952), .A2(n725), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n610), .A2(n702), .ZN(n612) );
  XNOR2_X1 U690 ( .A(n612), .B(n611), .ZN(G60) );
  NAND2_X1 U691 ( .A1(n616), .A2(n702), .ZN(n617) );
  XNOR2_X1 U692 ( .A(n617), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U693 ( .A(n618), .B(G101), .Z(G3) );
  NAND2_X1 U694 ( .A1(n623), .A2(n633), .ZN(n619) );
  XNOR2_X1 U695 ( .A(n619), .B(G104), .ZN(G6) );
  XOR2_X1 U696 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n621) );
  XNOR2_X1 U697 ( .A(G107), .B(KEYINPUT26), .ZN(n620) );
  XNOR2_X1 U698 ( .A(n621), .B(n620), .ZN(n622) );
  XOR2_X1 U699 ( .A(KEYINPUT27), .B(n622), .Z(n625) );
  NAND2_X1 U700 ( .A1(n623), .A2(n635), .ZN(n624) );
  XNOR2_X1 U701 ( .A(n625), .B(n624), .ZN(G9) );
  NOR2_X1 U702 ( .A1(n626), .A2(n630), .ZN(n628) );
  XNOR2_X1 U703 ( .A(KEYINPUT29), .B(KEYINPUT112), .ZN(n627) );
  XNOR2_X1 U704 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U705 ( .A(G128), .B(n629), .ZN(G30) );
  NOR2_X1 U706 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U707 ( .A(G146), .B(n632), .Z(G48) );
  NAND2_X1 U708 ( .A1(n636), .A2(n633), .ZN(n634) );
  XNOR2_X1 U709 ( .A(n634), .B(G113), .ZN(G15) );
  NAND2_X1 U710 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U711 ( .A(n637), .B(G116), .ZN(G18) );
  XNOR2_X1 U712 ( .A(G125), .B(n638), .ZN(n639) );
  XNOR2_X1 U713 ( .A(n639), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U714 ( .A(G134), .B(n640), .ZN(n641) );
  XNOR2_X1 U715 ( .A(n641), .B(KEYINPUT113), .ZN(G36) );
  NOR2_X1 U716 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U717 ( .A(n644), .B(KEYINPUT116), .ZN(n645) );
  NOR2_X1 U718 ( .A1(n646), .A2(n645), .ZN(n650) );
  NOR2_X1 U719 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U720 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U721 ( .A1(n651), .A2(n675), .ZN(n669) );
  INV_X1 U722 ( .A(n652), .ZN(n674) );
  NOR2_X1 U723 ( .A1(n569), .A2(n653), .ZN(n654) );
  XNOR2_X1 U724 ( .A(n654), .B(KEYINPUT49), .ZN(n655) );
  XNOR2_X1 U725 ( .A(n655), .B(KEYINPUT114), .ZN(n662) );
  NAND2_X1 U726 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U727 ( .A(KEYINPUT50), .B(n658), .Z(n659) );
  NOR2_X1 U728 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U729 ( .A1(n662), .A2(n661), .ZN(n664) );
  NAND2_X1 U730 ( .A1(n664), .A2(n663), .ZN(n666) );
  XOR2_X1 U731 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n665) );
  XNOR2_X1 U732 ( .A(n666), .B(n665), .ZN(n667) );
  NOR2_X1 U733 ( .A1(n674), .A2(n667), .ZN(n668) );
  NOR2_X1 U734 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U735 ( .A(n670), .B(KEYINPUT52), .ZN(n671) );
  NOR2_X1 U736 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U737 ( .A(n676), .B(KEYINPUT117), .ZN(n677) );
  NAND2_X1 U738 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U739 ( .A(KEYINPUT118), .B(KEYINPUT53), .ZN(n680) );
  XNOR2_X1 U740 ( .A(n681), .B(n680), .ZN(G75) );
  XOR2_X1 U741 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n682) );
  XNOR2_X1 U742 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U743 ( .A(n685), .B(n684), .ZN(n686) );
  NAND2_X1 U744 ( .A1(n686), .A2(n702), .ZN(n688) );
  XNOR2_X1 U745 ( .A(KEYINPUT56), .B(KEYINPUT119), .ZN(n687) );
  XNOR2_X1 U746 ( .A(n688), .B(n687), .ZN(G51) );
  INV_X1 U747 ( .A(n702), .ZN(n698) );
  XNOR2_X1 U748 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n691) );
  XNOR2_X1 U749 ( .A(n689), .B(KEYINPUT57), .ZN(n690) );
  XNOR2_X1 U750 ( .A(n691), .B(n690), .ZN(n693) );
  XOR2_X1 U751 ( .A(n693), .B(n692), .Z(n694) );
  NOR2_X1 U752 ( .A1(n698), .A2(n694), .ZN(G54) );
  XNOR2_X1 U753 ( .A(n696), .B(n695), .ZN(n697) );
  NOR2_X1 U754 ( .A1(n698), .A2(n697), .ZN(G63) );
  INV_X1 U755 ( .A(n699), .ZN(n700) );
  XNOR2_X1 U756 ( .A(n701), .B(n700), .ZN(n703) );
  XOR2_X1 U757 ( .A(n704), .B(G101), .Z(n705) );
  XNOR2_X1 U758 ( .A(n706), .B(n705), .ZN(n708) );
  NOR2_X1 U759 ( .A1(n708), .A2(n707), .ZN(n716) );
  NAND2_X1 U760 ( .A1(G224), .A2(G953), .ZN(n709) );
  XNOR2_X1 U761 ( .A(n709), .B(KEYINPUT61), .ZN(n710) );
  XNOR2_X1 U762 ( .A(KEYINPUT122), .B(n710), .ZN(n711) );
  NAND2_X1 U763 ( .A1(G898), .A2(n711), .ZN(n714) );
  NAND2_X1 U764 ( .A1(n712), .A2(n725), .ZN(n713) );
  NAND2_X1 U765 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U766 ( .A(n716), .B(n715), .ZN(G69) );
  XNOR2_X1 U767 ( .A(n718), .B(n717), .ZN(n724) );
  XNOR2_X1 U768 ( .A(n724), .B(G227), .ZN(n719) );
  XNOR2_X1 U769 ( .A(n719), .B(KEYINPUT123), .ZN(n720) );
  NAND2_X1 U770 ( .A1(n720), .A2(G900), .ZN(n721) );
  NAND2_X1 U771 ( .A1(G953), .A2(n721), .ZN(n722) );
  XNOR2_X1 U772 ( .A(n722), .B(KEYINPUT124), .ZN(n728) );
  XNOR2_X1 U773 ( .A(n724), .B(n723), .ZN(n726) );
  NAND2_X1 U774 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U775 ( .A1(n728), .A2(n727), .ZN(G72) );
  XNOR2_X1 U776 ( .A(G140), .B(n729), .ZN(G42) );
  XOR2_X1 U777 ( .A(G119), .B(KEYINPUT126), .Z(n730) );
  XNOR2_X1 U778 ( .A(n731), .B(n730), .ZN(G21) );
  XOR2_X1 U779 ( .A(n732), .B(G143), .Z(G45) );
  XOR2_X1 U780 ( .A(G110), .B(n733), .Z(G12) );
  XNOR2_X1 U781 ( .A(G122), .B(KEYINPUT125), .ZN(n735) );
  XNOR2_X1 U782 ( .A(n735), .B(n734), .ZN(G24) );
  XNOR2_X1 U783 ( .A(G137), .B(n736), .ZN(G39) );
  XOR2_X1 U784 ( .A(G131), .B(n737), .Z(n738) );
  XNOR2_X1 U785 ( .A(KEYINPUT127), .B(n738), .ZN(G33) );
endmodule

