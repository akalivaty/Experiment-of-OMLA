

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590;

  XNOR2_X1 U323 ( .A(n417), .B(n416), .ZN(n533) );
  INV_X1 U324 ( .A(KEYINPUT117), .ZN(n415) );
  XNOR2_X1 U325 ( .A(n415), .B(KEYINPUT48), .ZN(n416) );
  XNOR2_X1 U326 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U327 ( .A(n340), .B(n339), .ZN(n347) );
  XOR2_X1 U328 ( .A(KEYINPUT81), .B(n561), .Z(n546) );
  XNOR2_X1 U329 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n457) );
  XNOR2_X1 U330 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  XOR2_X1 U331 ( .A(G176GAT), .B(G183GAT), .Z(n292) );
  XNOR2_X1 U332 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n291) );
  XNOR2_X1 U333 ( .A(n292), .B(n291), .ZN(n296) );
  XOR2_X1 U334 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n294) );
  XNOR2_X1 U335 ( .A(KEYINPUT89), .B(KEYINPUT88), .ZN(n293) );
  XNOR2_X1 U336 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U337 ( .A(n296), .B(n295), .Z(n427) );
  XOR2_X1 U338 ( .A(KEYINPUT90), .B(KEYINPUT66), .Z(n298) );
  XNOR2_X1 U339 ( .A(KEYINPUT86), .B(KEYINPUT20), .ZN(n297) );
  XNOR2_X1 U340 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U341 ( .A(n427), .B(n299), .ZN(n309) );
  XOR2_X1 U342 ( .A(G120GAT), .B(G71GAT), .Z(n373) );
  XOR2_X1 U343 ( .A(G99GAT), .B(n373), .Z(n301) );
  XOR2_X1 U344 ( .A(KEYINPUT0), .B(G127GAT), .Z(n446) );
  XNOR2_X1 U345 ( .A(G43GAT), .B(n446), .ZN(n300) );
  XNOR2_X1 U346 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U347 ( .A(KEYINPUT85), .B(KEYINPUT87), .Z(n303) );
  NAND2_X1 U348 ( .A1(G227GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U349 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U350 ( .A(n305), .B(n304), .Z(n307) );
  XOR2_X1 U351 ( .A(G113GAT), .B(G15GAT), .Z(n350) );
  XOR2_X1 U352 ( .A(G190GAT), .B(G134GAT), .Z(n336) );
  XNOR2_X1 U353 ( .A(n350), .B(n336), .ZN(n306) );
  XNOR2_X1 U354 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U355 ( .A(n309), .B(n308), .Z(n464) );
  INV_X1 U356 ( .A(n464), .ZN(n536) );
  XOR2_X1 U357 ( .A(KEYINPUT22), .B(KEYINPUT92), .Z(n311) );
  XNOR2_X1 U358 ( .A(KEYINPUT94), .B(KEYINPUT24), .ZN(n310) );
  XNOR2_X1 U359 ( .A(n311), .B(n310), .ZN(n325) );
  XOR2_X1 U360 ( .A(G148GAT), .B(G78GAT), .Z(n372) );
  XOR2_X1 U361 ( .A(G106GAT), .B(n372), .Z(n313) );
  XOR2_X1 U362 ( .A(G218GAT), .B(G162GAT), .Z(n335) );
  XNOR2_X1 U363 ( .A(G50GAT), .B(n335), .ZN(n312) );
  XNOR2_X1 U364 ( .A(n313), .B(n312), .ZN(n318) );
  XNOR2_X1 U365 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n314) );
  XNOR2_X1 U366 ( .A(n314), .B(KEYINPUT2), .ZN(n445) );
  XOR2_X1 U367 ( .A(KEYINPUT23), .B(n445), .Z(n316) );
  NAND2_X1 U368 ( .A1(G228GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U369 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U370 ( .A(n318), .B(n317), .Z(n323) );
  XOR2_X1 U371 ( .A(G141GAT), .B(G22GAT), .Z(n351) );
  XOR2_X1 U372 ( .A(KEYINPUT93), .B(G211GAT), .Z(n320) );
  XNOR2_X1 U373 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n319) );
  XNOR2_X1 U374 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U375 ( .A(G197GAT), .B(n321), .ZN(n428) );
  XOR2_X1 U376 ( .A(n351), .B(n428), .Z(n322) );
  XNOR2_X1 U377 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U378 ( .A(n325), .B(n324), .Z(n472) );
  XOR2_X1 U379 ( .A(KEYINPUT77), .B(KEYINPUT10), .Z(n327) );
  XNOR2_X1 U380 ( .A(KEYINPUT78), .B(KEYINPUT80), .ZN(n326) );
  XOR2_X1 U381 ( .A(n327), .B(n326), .Z(n332) );
  INV_X1 U382 ( .A(G106GAT), .ZN(n331) );
  XOR2_X1 U383 ( .A(KEYINPUT74), .B(G92GAT), .Z(n329) );
  XNOR2_X1 U384 ( .A(G99GAT), .B(G85GAT), .ZN(n328) );
  XNOR2_X1 U385 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U386 ( .A(n331), .B(n330), .ZN(n380) );
  XNOR2_X1 U387 ( .A(n332), .B(n380), .ZN(n340) );
  XOR2_X1 U388 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n334) );
  NAND2_X1 U389 ( .A1(G232GAT), .A2(G233GAT), .ZN(n333) );
  XOR2_X1 U390 ( .A(n334), .B(n333), .Z(n338) );
  XNOR2_X1 U391 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U392 ( .A(G43GAT), .B(G29GAT), .Z(n342) );
  XNOR2_X1 U393 ( .A(KEYINPUT68), .B(G50GAT), .ZN(n341) );
  XNOR2_X1 U394 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U395 ( .A(n343), .B(KEYINPUT7), .Z(n345) );
  XNOR2_X1 U396 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n344) );
  XNOR2_X1 U397 ( .A(n345), .B(n344), .ZN(n363) );
  XNOR2_X1 U398 ( .A(n363), .B(KEYINPUT79), .ZN(n346) );
  XNOR2_X1 U399 ( .A(n347), .B(n346), .ZN(n561) );
  XOR2_X1 U400 ( .A(KEYINPUT70), .B(KEYINPUT67), .Z(n349) );
  XNOR2_X1 U401 ( .A(KEYINPUT30), .B(KEYINPUT71), .ZN(n348) );
  XNOR2_X1 U402 ( .A(n349), .B(n348), .ZN(n355) );
  XOR2_X1 U403 ( .A(G197GAT), .B(n350), .Z(n353) );
  XNOR2_X1 U404 ( .A(G169GAT), .B(n351), .ZN(n352) );
  XNOR2_X1 U405 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U406 ( .A(n355), .B(n354), .Z(n357) );
  NAND2_X1 U407 ( .A1(G229GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U408 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U409 ( .A(n358), .B(KEYINPUT29), .Z(n361) );
  XNOR2_X1 U410 ( .A(G1GAT), .B(KEYINPUT69), .ZN(n359) );
  XNOR2_X1 U411 ( .A(n359), .B(G8GAT), .ZN(n390) );
  XNOR2_X1 U412 ( .A(n390), .B(KEYINPUT72), .ZN(n360) );
  XNOR2_X1 U413 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U414 ( .A(n363), .B(n362), .Z(n407) );
  INV_X1 U415 ( .A(KEYINPUT31), .ZN(n364) );
  NAND2_X1 U416 ( .A1(KEYINPUT76), .A2(n364), .ZN(n367) );
  INV_X1 U417 ( .A(KEYINPUT76), .ZN(n365) );
  NAND2_X1 U418 ( .A1(n365), .A2(KEYINPUT31), .ZN(n366) );
  NAND2_X1 U419 ( .A1(n367), .A2(n366), .ZN(n369) );
  XNOR2_X1 U420 ( .A(G176GAT), .B(G204GAT), .ZN(n368) );
  XNOR2_X1 U421 ( .A(n369), .B(n368), .ZN(n371) );
  XNOR2_X1 U422 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n370) );
  XNOR2_X1 U423 ( .A(n370), .B(G64GAT), .ZN(n389) );
  XOR2_X1 U424 ( .A(n371), .B(n389), .Z(n375) );
  XNOR2_X1 U425 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U426 ( .A(n375), .B(n374), .ZN(n379) );
  XOR2_X1 U427 ( .A(KEYINPUT75), .B(KEYINPUT32), .Z(n377) );
  NAND2_X1 U428 ( .A1(G230GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U429 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U430 ( .A(n379), .B(n378), .ZN(n382) );
  XOR2_X1 U431 ( .A(n380), .B(KEYINPUT33), .Z(n381) );
  XNOR2_X1 U432 ( .A(n382), .B(n381), .ZN(n580) );
  INV_X1 U433 ( .A(KEYINPUT64), .ZN(n383) );
  XNOR2_X1 U434 ( .A(n580), .B(n383), .ZN(n384) );
  XOR2_X1 U435 ( .A(KEYINPUT41), .B(n384), .Z(n566) );
  INV_X1 U436 ( .A(n566), .ZN(n555) );
  NOR2_X1 U437 ( .A1(n407), .A2(n555), .ZN(n385) );
  XNOR2_X1 U438 ( .A(n385), .B(KEYINPUT46), .ZN(n386) );
  NOR2_X1 U439 ( .A1(n561), .A2(n386), .ZN(n405) );
  XOR2_X1 U440 ( .A(KEYINPUT84), .B(KEYINPUT82), .Z(n388) );
  XNOR2_X1 U441 ( .A(KEYINPUT15), .B(KEYINPUT83), .ZN(n387) );
  XNOR2_X1 U442 ( .A(n388), .B(n387), .ZN(n396) );
  XNOR2_X1 U443 ( .A(n390), .B(n389), .ZN(n394) );
  XOR2_X1 U444 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n392) );
  XNOR2_X1 U445 ( .A(G15GAT), .B(G183GAT), .ZN(n391) );
  XNOR2_X1 U446 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U447 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U448 ( .A(n396), .B(n395), .ZN(n404) );
  NAND2_X1 U449 ( .A1(G231GAT), .A2(G233GAT), .ZN(n402) );
  XOR2_X1 U450 ( .A(G155GAT), .B(G71GAT), .Z(n398) );
  XNOR2_X1 U451 ( .A(G22GAT), .B(G127GAT), .ZN(n397) );
  XNOR2_X1 U452 ( .A(n398), .B(n397), .ZN(n400) );
  XOR2_X1 U453 ( .A(G211GAT), .B(G78GAT), .Z(n399) );
  XNOR2_X1 U454 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U455 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U456 ( .A(n404), .B(n403), .Z(n571) );
  INV_X1 U457 ( .A(n571), .ZN(n584) );
  NAND2_X1 U458 ( .A1(n405), .A2(n584), .ZN(n406) );
  XNOR2_X1 U459 ( .A(n406), .B(KEYINPUT47), .ZN(n414) );
  BUF_X1 U460 ( .A(n407), .Z(n576) );
  XNOR2_X1 U461 ( .A(n576), .B(KEYINPUT73), .ZN(n564) );
  INV_X1 U462 ( .A(KEYINPUT36), .ZN(n408) );
  XNOR2_X1 U463 ( .A(n408), .B(n546), .ZN(n588) );
  NOR2_X1 U464 ( .A1(n584), .A2(n588), .ZN(n410) );
  XNOR2_X1 U465 ( .A(KEYINPUT45), .B(KEYINPUT116), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n410), .B(n409), .ZN(n411) );
  NAND2_X1 U467 ( .A1(n411), .A2(n580), .ZN(n412) );
  NOR2_X1 U468 ( .A1(n564), .A2(n412), .ZN(n413) );
  NOR2_X1 U469 ( .A1(n414), .A2(n413), .ZN(n417) );
  XOR2_X1 U470 ( .A(KEYINPUT79), .B(G190GAT), .Z(n419) );
  XNOR2_X1 U471 ( .A(G36GAT), .B(G8GAT), .ZN(n418) );
  XNOR2_X1 U472 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U473 ( .A(KEYINPUT97), .B(G64GAT), .Z(n421) );
  XNOR2_X1 U474 ( .A(G218GAT), .B(G92GAT), .ZN(n420) );
  XNOR2_X1 U475 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U476 ( .A(n423), .B(n422), .Z(n425) );
  NAND2_X1 U477 ( .A1(G226GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U478 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U479 ( .A(n427), .B(n426), .ZN(n430) );
  INV_X1 U480 ( .A(n428), .ZN(n429) );
  XOR2_X1 U481 ( .A(n430), .B(n429), .Z(n525) );
  NOR2_X1 U482 ( .A1(n533), .A2(n525), .ZN(n431) );
  XNOR2_X1 U483 ( .A(n431), .B(KEYINPUT54), .ZN(n453) );
  XOR2_X1 U484 ( .A(KEYINPUT78), .B(G148GAT), .Z(n433) );
  XNOR2_X1 U485 ( .A(G29GAT), .B(G134GAT), .ZN(n432) );
  XNOR2_X1 U486 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U487 ( .A(KEYINPUT4), .B(G120GAT), .Z(n435) );
  XNOR2_X1 U488 ( .A(G141GAT), .B(G113GAT), .ZN(n434) );
  XNOR2_X1 U489 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U490 ( .A(n437), .B(n436), .Z(n442) );
  XOR2_X1 U491 ( .A(KEYINPUT6), .B(G57GAT), .Z(n439) );
  NAND2_X1 U492 ( .A1(G225GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U494 ( .A(KEYINPUT1), .B(n440), .ZN(n441) );
  XNOR2_X1 U495 ( .A(n442), .B(n441), .ZN(n452) );
  XOR2_X1 U496 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n444) );
  XNOR2_X1 U497 ( .A(G1GAT), .B(KEYINPUT95), .ZN(n443) );
  XNOR2_X1 U498 ( .A(n444), .B(n443), .ZN(n450) );
  XOR2_X1 U499 ( .A(G85GAT), .B(G162GAT), .Z(n448) );
  XNOR2_X1 U500 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U501 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U502 ( .A(n450), .B(n449), .Z(n451) );
  XNOR2_X1 U503 ( .A(n452), .B(n451), .ZN(n523) );
  NAND2_X1 U504 ( .A1(n453), .A2(n523), .ZN(n454) );
  XNOR2_X1 U505 ( .A(n454), .B(KEYINPUT65), .ZN(n575) );
  AND2_X1 U506 ( .A1(n472), .A2(n575), .ZN(n455) );
  XNOR2_X1 U507 ( .A(n455), .B(KEYINPUT55), .ZN(n456) );
  NOR2_X2 U508 ( .A1(n536), .A2(n456), .ZN(n572) );
  NAND2_X1 U509 ( .A1(n572), .A2(n546), .ZN(n458) );
  NAND2_X1 U510 ( .A1(n580), .A2(n564), .ZN(n497) );
  NOR2_X1 U511 ( .A1(n546), .A2(n584), .ZN(n459) );
  XNOR2_X1 U512 ( .A(n459), .B(KEYINPUT16), .ZN(n482) );
  INV_X1 U513 ( .A(n525), .ZN(n463) );
  XOR2_X1 U514 ( .A(KEYINPUT27), .B(KEYINPUT98), .Z(n460) );
  XOR2_X1 U515 ( .A(n463), .B(n460), .Z(n473) );
  NOR2_X1 U516 ( .A1(n472), .A2(n464), .ZN(n461) );
  XNOR2_X1 U517 ( .A(KEYINPUT26), .B(n461), .ZN(n574) );
  NAND2_X1 U518 ( .A1(n473), .A2(n574), .ZN(n462) );
  XNOR2_X1 U519 ( .A(KEYINPUT101), .B(n462), .ZN(n469) );
  NAND2_X1 U520 ( .A1(n464), .A2(n463), .ZN(n465) );
  NAND2_X1 U521 ( .A1(n465), .A2(n472), .ZN(n466) );
  XNOR2_X1 U522 ( .A(n466), .B(KEYINPUT102), .ZN(n467) );
  XNOR2_X1 U523 ( .A(n467), .B(KEYINPUT25), .ZN(n468) );
  NOR2_X1 U524 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U525 ( .A(n470), .B(KEYINPUT103), .ZN(n471) );
  NAND2_X1 U526 ( .A1(n471), .A2(n523), .ZN(n481) );
  XNOR2_X1 U527 ( .A(n472), .B(KEYINPUT28), .ZN(n534) );
  INV_X1 U528 ( .A(n534), .ZN(n476) );
  INV_X1 U529 ( .A(n473), .ZN(n474) );
  NOR2_X1 U530 ( .A1(n474), .A2(n523), .ZN(n475) );
  XNOR2_X1 U531 ( .A(n475), .B(KEYINPUT99), .ZN(n532) );
  NOR2_X1 U532 ( .A1(n476), .A2(n532), .ZN(n477) );
  XNOR2_X1 U533 ( .A(n477), .B(KEYINPUT100), .ZN(n479) );
  XOR2_X1 U534 ( .A(n536), .B(KEYINPUT91), .Z(n478) );
  NAND2_X1 U535 ( .A1(n479), .A2(n478), .ZN(n480) );
  NAND2_X1 U536 ( .A1(n481), .A2(n480), .ZN(n494) );
  NAND2_X1 U537 ( .A1(n482), .A2(n494), .ZN(n509) );
  OR2_X1 U538 ( .A1(n497), .A2(n509), .ZN(n490) );
  NOR2_X1 U539 ( .A1(n523), .A2(n490), .ZN(n484) );
  XNOR2_X1 U540 ( .A(KEYINPUT34), .B(KEYINPUT104), .ZN(n483) );
  XNOR2_X1 U541 ( .A(n484), .B(n483), .ZN(n485) );
  XOR2_X1 U542 ( .A(G1GAT), .B(n485), .Z(G1324GAT) );
  NOR2_X1 U543 ( .A1(n525), .A2(n490), .ZN(n486) );
  XOR2_X1 U544 ( .A(G8GAT), .B(n486), .Z(G1325GAT) );
  NOR2_X1 U545 ( .A1(n536), .A2(n490), .ZN(n488) );
  XNOR2_X1 U546 ( .A(KEYINPUT105), .B(KEYINPUT35), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U548 ( .A(G15GAT), .B(n489), .Z(G1326GAT) );
  NOR2_X1 U549 ( .A1(n534), .A2(n490), .ZN(n491) );
  XOR2_X1 U550 ( .A(KEYINPUT106), .B(n491), .Z(n492) );
  XNOR2_X1 U551 ( .A(G22GAT), .B(n492), .ZN(G1327GAT) );
  NOR2_X1 U552 ( .A1(n588), .A2(n571), .ZN(n493) );
  NAND2_X1 U553 ( .A1(n494), .A2(n493), .ZN(n495) );
  XNOR2_X1 U554 ( .A(KEYINPUT107), .B(n495), .ZN(n496) );
  XNOR2_X1 U555 ( .A(KEYINPUT37), .B(n496), .ZN(n521) );
  NOR2_X1 U556 ( .A1(n521), .A2(n497), .ZN(n498) );
  XOR2_X1 U557 ( .A(KEYINPUT108), .B(n498), .Z(n499) );
  XNOR2_X1 U558 ( .A(KEYINPUT38), .B(n499), .ZN(n507) );
  NOR2_X1 U559 ( .A1(n523), .A2(n507), .ZN(n501) );
  XNOR2_X1 U560 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n501), .B(n500), .ZN(G1328GAT) );
  NOR2_X1 U562 ( .A1(n525), .A2(n507), .ZN(n502) );
  XOR2_X1 U563 ( .A(G36GAT), .B(n502), .Z(G1329GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT110), .B(KEYINPUT40), .Z(n504) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(KEYINPUT109), .ZN(n503) );
  XNOR2_X1 U566 ( .A(n504), .B(n503), .ZN(n506) );
  NOR2_X1 U567 ( .A1(n536), .A2(n507), .ZN(n505) );
  XOR2_X1 U568 ( .A(n506), .B(n505), .Z(G1330GAT) );
  NOR2_X1 U569 ( .A1(n534), .A2(n507), .ZN(n508) );
  XOR2_X1 U570 ( .A(G50GAT), .B(n508), .Z(G1331GAT) );
  NAND2_X1 U571 ( .A1(n576), .A2(n566), .ZN(n520) );
  OR2_X1 U572 ( .A1(n520), .A2(n509), .ZN(n517) );
  NOR2_X1 U573 ( .A1(n523), .A2(n517), .ZN(n511) );
  XNOR2_X1 U574 ( .A(KEYINPUT111), .B(KEYINPUT42), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U576 ( .A(G57GAT), .B(n512), .ZN(G1332GAT) );
  NOR2_X1 U577 ( .A1(n525), .A2(n517), .ZN(n513) );
  XOR2_X1 U578 ( .A(KEYINPUT112), .B(n513), .Z(n514) );
  XNOR2_X1 U579 ( .A(G64GAT), .B(n514), .ZN(G1333GAT) );
  NOR2_X1 U580 ( .A1(n536), .A2(n517), .ZN(n516) );
  XNOR2_X1 U581 ( .A(G71GAT), .B(KEYINPUT113), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(G1334GAT) );
  NOR2_X1 U583 ( .A1(n534), .A2(n517), .ZN(n519) );
  XNOR2_X1 U584 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  NOR2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n522) );
  XOR2_X1 U587 ( .A(KEYINPUT114), .B(n522), .Z(n528) );
  NOR2_X1 U588 ( .A1(n528), .A2(n523), .ZN(n524) );
  XOR2_X1 U589 ( .A(G85GAT), .B(n524), .Z(G1336GAT) );
  NOR2_X1 U590 ( .A1(n528), .A2(n525), .ZN(n526) );
  XOR2_X1 U591 ( .A(G92GAT), .B(n526), .Z(G1337GAT) );
  NOR2_X1 U592 ( .A1(n536), .A2(n528), .ZN(n527) );
  XOR2_X1 U593 ( .A(G99GAT), .B(n527), .Z(G1338GAT) );
  NOR2_X1 U594 ( .A1(n528), .A2(n534), .ZN(n530) );
  XNOR2_X1 U595 ( .A(KEYINPUT115), .B(KEYINPUT44), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  NOR2_X1 U598 ( .A1(n533), .A2(n532), .ZN(n551) );
  NAND2_X1 U599 ( .A1(n551), .A2(n534), .ZN(n535) );
  NOR2_X1 U600 ( .A1(n536), .A2(n535), .ZN(n547) );
  NAND2_X1 U601 ( .A1(n547), .A2(n564), .ZN(n537) );
  XNOR2_X1 U602 ( .A(G113GAT), .B(n537), .ZN(G1340GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT49), .B(KEYINPUT119), .Z(n539) );
  NAND2_X1 U604 ( .A1(n547), .A2(n566), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(n541) );
  XOR2_X1 U606 ( .A(G120GAT), .B(KEYINPUT118), .Z(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  XNOR2_X1 U608 ( .A(G127GAT), .B(KEYINPUT121), .ZN(n545) );
  XOR2_X1 U609 ( .A(KEYINPUT50), .B(KEYINPUT120), .Z(n543) );
  NAND2_X1 U610 ( .A1(n547), .A2(n571), .ZN(n542) );
  XNOR2_X1 U611 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT51), .B(KEYINPUT122), .Z(n549) );
  NAND2_X1 U614 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U616 ( .A(G134GAT), .B(n550), .ZN(G1343GAT) );
  NAND2_X1 U617 ( .A1(n551), .A2(n574), .ZN(n560) );
  NOR2_X1 U618 ( .A1(n576), .A2(n560), .ZN(n553) );
  XNOR2_X1 U619 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(G141GAT), .B(n554), .ZN(G1344GAT) );
  NOR2_X1 U622 ( .A1(n555), .A2(n560), .ZN(n557) );
  XNOR2_X1 U623 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U625 ( .A(G148GAT), .B(n558), .ZN(G1345GAT) );
  NOR2_X1 U626 ( .A1(n584), .A2(n560), .ZN(n559) );
  XOR2_X1 U627 ( .A(G155GAT), .B(n559), .Z(G1346GAT) );
  INV_X1 U628 ( .A(n560), .ZN(n562) );
  NAND2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U631 ( .A1(n564), .A2(n572), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U633 ( .A1(n572), .A2(n566), .ZN(n568) );
  XOR2_X1 U634 ( .A(G176GAT), .B(KEYINPUT125), .Z(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n570) );
  XOR2_X1 U636 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(G1349GAT) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n587) );
  NOR2_X1 U641 ( .A1(n576), .A2(n587), .ZN(n578) );
  XNOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(n579), .ZN(G1352GAT) );
  NOR2_X1 U645 ( .A1(n580), .A2(n587), .ZN(n582) );
  XNOR2_X1 U646 ( .A(KEYINPUT126), .B(KEYINPUT61), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(n583), .ZN(G1353GAT) );
  NOR2_X1 U649 ( .A1(n584), .A2(n587), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1354GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U653 ( .A(KEYINPUT62), .B(n589), .Z(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

