//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 0 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 1 0 1 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1330, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1391, new_n1392, new_n1393, new_n1394, new_n1395,
    new_n1396, new_n1397;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  NOR3_X1   g0004(.A1(new_n202), .A2(G77), .A3(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n207), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT1), .ZN(new_n215));
  OR3_X1    g0015(.A1(new_n207), .A2(KEYINPUT65), .A3(G13), .ZN(new_n216));
  OAI21_X1  g0016(.A(KEYINPUT65), .B1(new_n207), .B2(G13), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT0), .Z(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n204), .A2(G50), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  AOI211_X1 g0025(.A(new_n215), .B(new_n220), .C1(new_n223), .C2(new_n225), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G232), .ZN(new_n228));
  XOR2_X1   g0028(.A(KEYINPUT2), .B(G226), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G264), .B(G270), .Z(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n230), .B(new_n233), .Z(G358));
  XOR2_X1   g0034(.A(G68), .B(G77), .Z(new_n235));
  XNOR2_X1  g0035(.A(G50), .B(G58), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G351));
  INV_X1    g0041(.A(G41), .ZN(new_n242));
  INV_X1    g0042(.A(G45), .ZN(new_n243));
  AOI21_X1  g0043(.A(G1), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g0044(.A1(G33), .A2(G41), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n245), .A2(G1), .A3(G13), .ZN(new_n246));
  AND3_X1   g0046(.A1(new_n244), .A2(new_n246), .A3(G274), .ZN(new_n247));
  AOI21_X1  g0047(.A(new_n221), .B1(G33), .B2(G41), .ZN(new_n248));
  AND2_X1   g0048(.A1(KEYINPUT66), .A2(G1), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT66), .A2(G1), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G41), .A2(G45), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n248), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n247), .B1(new_n254), .B2(G226), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT3), .B(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G1698), .ZN(new_n257));
  INV_X1    g0057(.A(G223), .ZN(new_n258));
  INV_X1    g0058(.A(G77), .ZN(new_n259));
  OAI22_X1  g0059(.A1(new_n257), .A2(new_n258), .B1(new_n259), .B2(new_n256), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT67), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n256), .A2(new_n261), .A3(G222), .A4(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n256), .A2(G222), .A3(new_n262), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT67), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n260), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n255), .B1(new_n266), .B2(new_n246), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G200), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n222), .B1(new_n201), .B2(new_n203), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT8), .B(G58), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n222), .A2(G33), .ZN(new_n271));
  INV_X1    g0071(.A(G150), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n222), .A2(new_n273), .ZN(new_n274));
  OAI22_X1  g0074(.A1(new_n270), .A2(new_n271), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n269), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n221), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  NOR3_X1   g0080(.A1(new_n249), .A2(new_n250), .A3(new_n222), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(new_n278), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G50), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT66), .ZN(new_n284));
  INV_X1    g0084(.A(G1), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(KEYINPUT66), .A2(G1), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n286), .A2(G13), .A3(G20), .A4(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n283), .B1(G50), .B2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n280), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(KEYINPUT9), .ZN(new_n291));
  OAI221_X1 g0091(.A(new_n283), .B1(G50), .B2(new_n288), .C1(new_n276), .C2(new_n279), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT9), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI211_X1 g0094(.A(G190), .B(new_n255), .C1(new_n266), .C2(new_n246), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n268), .A2(new_n291), .A3(new_n294), .A4(new_n295), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n296), .B(KEYINPUT10), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n267), .A2(G179), .ZN(new_n298));
  INV_X1    g0098(.A(G169), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n267), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n298), .A2(new_n292), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G274), .ZN(new_n303));
  AND2_X1   g0103(.A1(G1), .A2(G13), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n303), .B1(new_n304), .B2(new_n245), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n244), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n286), .A2(new_n287), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n246), .B1(new_n307), .B2(new_n252), .ZN(new_n308));
  INV_X1    g0108(.A(G244), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n306), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n256), .A2(G232), .A3(new_n262), .ZN(new_n311));
  INV_X1    g0111(.A(G107), .ZN(new_n312));
  INV_X1    g0112(.A(G238), .ZN(new_n313));
  OAI221_X1 g0113(.A(new_n311), .B1(new_n312), .B2(new_n256), .C1(new_n257), .C2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n310), .B1(new_n314), .B2(new_n248), .ZN(new_n315));
  INV_X1    g0115(.A(G179), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI22_X1  g0117(.A1(new_n270), .A2(new_n274), .B1(new_n222), .B2(new_n259), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT15), .B(G87), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n319), .A2(new_n271), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n278), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n288), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n259), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n282), .A2(G77), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n321), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n317), .B(new_n325), .C1(G169), .C2(new_n315), .ZN(new_n326));
  INV_X1    g0126(.A(G200), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n315), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n315), .A2(G190), .ZN(new_n329));
  INV_X1    g0129(.A(new_n325), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n326), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n302), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT16), .ZN(new_n334));
  INV_X1    g0134(.A(G68), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT7), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n336), .B1(new_n256), .B2(G20), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT3), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n338), .A2(G33), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n273), .A2(KEYINPUT3), .ZN(new_n340));
  OAI211_X1 g0140(.A(KEYINPUT7), .B(new_n222), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n335), .B1(new_n337), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G58), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n343), .A2(new_n335), .ZN(new_n344));
  OAI21_X1  g0144(.A(G20), .B1(new_n344), .B2(new_n203), .ZN(new_n345));
  INV_X1    g0145(.A(new_n274), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G159), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n334), .B1(new_n342), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT71), .ZN(new_n350));
  INV_X1    g0150(.A(new_n348), .ZN(new_n351));
  AND3_X1   g0151(.A1(new_n337), .A2(KEYINPUT70), .A3(new_n341), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT70), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n353), .B(new_n336), .C1(new_n256), .C2(G20), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G68), .ZN(new_n355));
  OAI211_X1 g0155(.A(KEYINPUT16), .B(new_n351), .C1(new_n352), .C2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT71), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n357), .B(new_n334), .C1(new_n342), .C2(new_n348), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n350), .A2(new_n278), .A3(new_n356), .A4(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n288), .A2(new_n270), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(new_n282), .B2(new_n270), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n273), .A2(KEYINPUT3), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n338), .A2(G33), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n363), .A2(new_n364), .A3(G226), .A4(G1698), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n363), .A2(new_n364), .A3(G223), .A4(new_n262), .ZN(new_n366));
  NAND2_X1  g0166(.A1(G33), .A2(G87), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n248), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT72), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT72), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n368), .A2(new_n371), .A3(new_n248), .ZN(new_n372));
  OAI211_X1 g0172(.A(G232), .B(new_n246), .C1(new_n307), .C2(new_n252), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n373), .A2(new_n316), .A3(new_n306), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n370), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n368), .A2(new_n248), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n373), .A2(new_n306), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n299), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n362), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT18), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n377), .A2(G190), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n383), .A2(new_n370), .A3(new_n372), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n327), .B1(new_n376), .B2(new_n377), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n359), .A2(new_n386), .A3(new_n361), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT17), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n379), .B1(new_n359), .B2(new_n361), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT18), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n359), .A2(new_n386), .A3(new_n361), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT17), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n382), .A2(new_n388), .A3(new_n391), .A4(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n335), .A2(G20), .ZN(new_n397));
  INV_X1    g0197(.A(G50), .ZN(new_n398));
  OAI221_X1 g0198(.A(new_n397), .B1(new_n271), .B2(new_n259), .C1(new_n398), .C2(new_n274), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n278), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT11), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT11), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n399), .A2(new_n402), .A3(new_n278), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n288), .A2(G68), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT12), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n405), .B(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n282), .A2(G68), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n404), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n363), .A2(new_n364), .A3(G232), .A4(G1698), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n363), .A2(new_n364), .A3(G226), .A4(new_n262), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G33), .A2(G97), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n413), .A2(new_n248), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n306), .B1(new_n308), .B2(new_n313), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT13), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n247), .B1(new_n254), .B2(G238), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT13), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n413), .A2(new_n248), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n409), .B1(G200), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT69), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n416), .A2(KEYINPUT68), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n418), .B1(new_n417), .B2(new_n419), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT68), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n424), .A2(new_n427), .A3(G190), .A4(new_n420), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n422), .A2(new_n423), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n423), .B1(new_n422), .B2(new_n428), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n431));
  OAI21_X1  g0231(.A(G169), .B1(new_n431), .B2(new_n425), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT14), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n421), .A2(KEYINPUT14), .A3(G169), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n425), .A2(new_n426), .ZN(new_n436));
  AOI211_X1 g0236(.A(KEYINPUT68), .B(new_n418), .C1(new_n417), .C2(new_n419), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n431), .A2(new_n316), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n434), .A2(new_n435), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n404), .A2(new_n407), .A3(new_n408), .ZN(new_n441));
  OAI22_X1  g0241(.A1(new_n429), .A2(new_n430), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n333), .A2(new_n396), .A3(new_n443), .ZN(new_n444));
  XNOR2_X1  g0244(.A(KEYINPUT5), .B(G41), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n305), .A2(new_n251), .A3(new_n445), .A4(G45), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n286), .A2(G45), .A3(new_n287), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n242), .A2(KEYINPUT5), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT5), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(G41), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g0251(.A(G264), .B(new_n246), .C1(new_n447), .C2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT84), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n251), .A2(new_n445), .A3(G45), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n455), .A2(KEYINPUT84), .A3(G264), .A4(new_n246), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT85), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n363), .A2(new_n364), .A3(G257), .A4(G1698), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n363), .A2(new_n364), .A3(G250), .A4(new_n262), .ZN(new_n460));
  INV_X1    g0260(.A(G294), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n459), .B(new_n460), .C1(new_n273), .C2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n248), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n457), .A2(new_n458), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n458), .B1(new_n457), .B2(new_n463), .ZN(new_n465));
  OAI211_X1 g0265(.A(G179), .B(new_n446), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n463), .A2(KEYINPUT83), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT83), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n462), .A2(new_n468), .A3(new_n248), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n467), .A2(new_n457), .A3(new_n446), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G169), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n312), .A2(G20), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT80), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n473), .A2(new_n474), .A3(KEYINPUT23), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G33), .A2(G116), .ZN(new_n477));
  OAI22_X1  g0277(.A1(new_n473), .A2(KEYINPUT23), .B1(G20), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n474), .B1(new_n473), .B2(KEYINPUT23), .ZN(new_n479));
  NOR3_X1   g0279(.A1(new_n476), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n363), .A2(new_n364), .A3(new_n222), .A4(G87), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT22), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT22), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n256), .A2(new_n483), .A3(new_n222), .A4(G87), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  XOR2_X1   g0285(.A(KEYINPUT79), .B(KEYINPUT24), .Z(new_n486));
  AND3_X1   g0286(.A1(new_n480), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n486), .B1(new_n480), .B2(new_n485), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n278), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT81), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT81), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n491), .B(new_n278), .C1(new_n487), .C2(new_n488), .ZN(new_n492));
  XNOR2_X1  g0292(.A(KEYINPUT82), .B(KEYINPUT25), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n322), .A2(new_n312), .A3(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT82), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n495), .B(KEYINPUT25), .C1(new_n288), .C2(G107), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n286), .A2(G33), .A3(new_n287), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n288), .A2(new_n279), .A3(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT74), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n288), .A2(new_n279), .A3(new_n498), .A4(KEYINPUT74), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n497), .B1(new_n503), .B2(G107), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n490), .A2(new_n492), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n472), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n470), .A2(G190), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n446), .B1(new_n464), .B2(new_n465), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n507), .B1(new_n508), .B2(new_n327), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n506), .B1(new_n505), .B2(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(G270), .B(new_n246), .C1(new_n447), .C2(new_n451), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n446), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(G303), .B1(new_n339), .B2(new_n340), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n363), .A2(new_n364), .A3(G264), .A4(G1698), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n363), .A2(new_n364), .A3(G257), .A4(new_n262), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n248), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n299), .B1(new_n513), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n281), .A2(G13), .B1(new_n498), .B2(G116), .ZN(new_n520));
  INV_X1    g0320(.A(G116), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n521), .B1(new_n288), .B2(new_n279), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n277), .A2(new_n221), .B1(G20), .B2(new_n521), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G283), .ZN(new_n524));
  INV_X1    g0324(.A(G97), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n524), .B(new_n222), .C1(G33), .C2(new_n525), .ZN(new_n526));
  AND3_X1   g0326(.A1(new_n523), .A2(KEYINPUT20), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT20), .B1(new_n523), .B2(new_n526), .ZN(new_n528));
  OAI22_X1  g0328(.A1(new_n520), .A2(new_n522), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT78), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n288), .A2(new_n279), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G116), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n498), .A2(G116), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n288), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n523), .A2(new_n526), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT20), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n523), .A2(KEYINPUT20), .A3(new_n526), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT78), .B1(new_n536), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n519), .B1(new_n531), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT21), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n517), .A2(new_n248), .ZN(new_n546));
  OAI211_X1 g0346(.A(KEYINPUT21), .B(G169), .C1(new_n546), .C2(new_n512), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n518), .A2(G179), .A3(new_n446), .A4(new_n511), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n529), .A2(new_n530), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n536), .A2(KEYINPUT78), .A3(new_n541), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n513), .A2(new_n518), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(G200), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n513), .A2(G190), .A3(new_n518), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n555), .A2(new_n550), .A3(new_n556), .A4(new_n551), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n545), .A2(new_n553), .A3(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n363), .A2(new_n364), .A3(new_n222), .A4(G68), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT19), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n271), .B2(new_n525), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n222), .ZN(new_n564));
  NOR4_X1   g0364(.A1(KEYINPUT76), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT76), .ZN(new_n566));
  NOR2_X1   g0366(.A1(G87), .A2(G97), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n566), .B1(new_n567), .B2(new_n312), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n564), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT77), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n562), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(KEYINPUT77), .B(new_n564), .C1(new_n565), .C2(new_n568), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n279), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n319), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n574), .A2(new_n288), .ZN(new_n575));
  INV_X1    g0375(.A(G87), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n576), .B1(new_n501), .B2(new_n502), .ZN(new_n577));
  NOR3_X1   g0377(.A1(new_n573), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n447), .A2(G250), .A3(new_n246), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n305), .A2(G45), .A3(new_n251), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n313), .A2(new_n262), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n309), .A2(G1698), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n363), .A2(new_n582), .A3(new_n364), .A4(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n246), .B1(new_n584), .B2(new_n477), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(G190), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n581), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n579), .A2(new_n580), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n589), .A2(new_n585), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n588), .B1(new_n590), .B2(G200), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n559), .A2(new_n561), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n576), .A2(new_n525), .A3(new_n312), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT76), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n567), .A2(new_n566), .A3(new_n312), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n594), .A2(new_n595), .B1(new_n222), .B2(new_n563), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n592), .B1(new_n596), .B2(KEYINPUT77), .ZN(new_n597));
  INV_X1    g0397(.A(new_n572), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n278), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n575), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n503), .A2(new_n574), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(G169), .B1(new_n589), .B2(new_n585), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n581), .A2(new_n586), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n603), .B1(new_n604), .B2(new_n316), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n578), .A2(new_n591), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n337), .A2(new_n341), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(G107), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT6), .ZN(new_n609));
  AND2_X1   g0409(.A1(G97), .A2(G107), .ZN(new_n610));
  NOR2_X1   g0410(.A1(G97), .A2(G107), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n312), .A2(KEYINPUT6), .A3(G97), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n222), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n274), .A2(new_n259), .ZN(new_n615));
  OAI21_X1  g0415(.A(KEYINPUT73), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT73), .ZN(new_n617));
  INV_X1    g0417(.A(new_n615), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n312), .A2(KEYINPUT6), .A3(G97), .ZN(new_n619));
  XNOR2_X1  g0419(.A(G97), .B(G107), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n619), .B1(new_n620), .B2(new_n609), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n617), .B(new_n618), .C1(new_n621), .C2(new_n222), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n608), .A2(new_n616), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n288), .A2(new_n525), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n501), .A2(G97), .A3(new_n502), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n623), .A2(new_n278), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n363), .A2(new_n364), .A3(G244), .A4(new_n262), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT4), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n256), .A2(KEYINPUT4), .A3(G244), .A4(new_n262), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n256), .A2(G250), .A3(G1698), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n629), .A2(new_n630), .A3(new_n524), .A4(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n248), .ZN(new_n633));
  OAI211_X1 g0433(.A(G257), .B(new_n246), .C1(new_n447), .C2(new_n451), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n446), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT75), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(new_n638), .A3(G200), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n635), .B1(new_n248), .B2(new_n632), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT75), .B1(new_n640), .B2(new_n327), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(G190), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n626), .A2(new_n639), .A3(new_n641), .A4(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n623), .A2(new_n278), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n625), .A2(new_n624), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n637), .A2(new_n299), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n640), .A2(new_n316), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n606), .A2(new_n643), .A3(new_n649), .ZN(new_n650));
  NOR4_X1   g0450(.A1(new_n444), .A2(new_n510), .A3(new_n558), .A4(new_n650), .ZN(G372));
  INV_X1    g0451(.A(new_n301), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n392), .B(KEYINPUT17), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n420), .A2(G190), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n436), .A2(new_n437), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(G200), .B1(new_n431), .B2(new_n425), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n441), .ZN(new_n657));
  OAI21_X1  g0457(.A(KEYINPUT69), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n422), .A2(new_n423), .A3(new_n428), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n326), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n439), .A2(new_n424), .A3(new_n427), .ZN(new_n661));
  AOI21_X1  g0461(.A(KEYINPUT14), .B1(new_n421), .B2(G169), .ZN(new_n662));
  AOI211_X1 g0462(.A(new_n433), .B(new_n299), .C1(new_n416), .C2(new_n420), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n409), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n653), .B1(new_n660), .B2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n390), .B1(new_n362), .B2(new_n380), .ZN(new_n668));
  AOI211_X1 g0468(.A(KEYINPUT18), .B(new_n379), .C1(new_n359), .C2(new_n361), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n652), .B1(new_n671), .B2(new_n297), .ZN(new_n672));
  AOI21_X1  g0472(.A(KEYINPUT21), .B1(new_n552), .B2(new_n519), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n547), .A2(new_n548), .B1(new_n550), .B2(new_n551), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n506), .A2(new_n675), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n470), .A2(G190), .ZN(new_n677));
  INV_X1    g0477(.A(new_n446), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n457), .A2(new_n463), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(KEYINPUT85), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n457), .A2(new_n458), .A3(new_n463), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n678), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n677), .B1(new_n682), .B2(G200), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n490), .A2(new_n492), .A3(new_n504), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n578), .A2(new_n591), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n299), .B1(new_n581), .B2(new_n586), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n589), .A2(new_n585), .A3(new_n316), .ZN(new_n688));
  OAI21_X1  g0488(.A(KEYINPUT86), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT86), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n690), .B(new_n603), .C1(new_n604), .C2(new_n316), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n602), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n643), .A2(new_n649), .A3(new_n686), .A4(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n676), .A2(new_n685), .A3(new_n694), .ZN(new_n695));
  AND3_X1   g0495(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n606), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT26), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT26), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n696), .A2(new_n699), .A3(new_n686), .A4(new_n692), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n698), .A2(new_n692), .A3(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n695), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n672), .B1(new_n444), .B2(new_n702), .ZN(G369));
  INV_X1    g0503(.A(KEYINPUT89), .ZN(new_n704));
  INV_X1    g0504(.A(G13), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G20), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT27), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n706), .A2(new_n286), .A3(new_n707), .A4(new_n287), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT87), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n251), .A2(KEYINPUT87), .A3(new_n707), .A4(new_n706), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT88), .ZN(new_n713));
  INV_X1    g0513(.A(G213), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n251), .A2(new_n706), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n714), .B1(new_n715), .B2(KEYINPUT27), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n712), .A2(new_n713), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n713), .B1(new_n712), .B2(new_n716), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n704), .B1(new_n719), .B2(G343), .ZN(new_n720));
  INV_X1    g0520(.A(G343), .ZN(new_n721));
  NOR4_X1   g0521(.A1(new_n717), .A2(new_n718), .A3(KEYINPUT89), .A4(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n723), .B1(new_n550), .B2(new_n551), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n724), .B1(new_n673), .B2(new_n674), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(new_n558), .B2(new_n724), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G330), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n685), .B(new_n506), .C1(new_n684), .C2(new_n723), .ZN(new_n728));
  INV_X1    g0528(.A(new_n506), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n717), .A2(new_n718), .ZN(new_n730));
  OAI21_X1  g0530(.A(KEYINPUT89), .B1(new_n730), .B2(new_n721), .ZN(new_n731));
  INV_X1    g0531(.A(new_n722), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n727), .B1(new_n728), .B2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n733), .A2(new_n675), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(new_n685), .A3(new_n506), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n729), .A2(new_n723), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n736), .A2(new_n740), .ZN(G399));
  INV_X1    g0541(.A(new_n218), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n742), .A2(KEYINPUT90), .A3(G41), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT90), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n744), .B1(new_n218), .B2(new_n242), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n565), .A2(new_n568), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n521), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n747), .A2(G1), .A3(new_n750), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n751), .B(KEYINPUT91), .C1(new_n224), .C2(new_n747), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(KEYINPUT91), .B2(new_n751), .ZN(new_n753));
  XOR2_X1   g0553(.A(new_n753), .B(KEYINPUT28), .Z(new_n754));
  NAND2_X1  g0554(.A1(new_n692), .A2(new_n686), .ZN(new_n755));
  OAI21_X1  g0555(.A(KEYINPUT26), .B1(new_n755), .B2(new_n649), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n696), .A2(new_n606), .A3(new_n699), .ZN(new_n757));
  AND3_X1   g0557(.A1(new_n756), .A2(new_n692), .A3(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n676), .A2(new_n694), .A3(new_n685), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(KEYINPUT94), .B1(new_n760), .B2(new_n723), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT94), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n762), .B(new_n733), .C1(new_n758), .C2(new_n759), .ZN(new_n763));
  OAI21_X1  g0563(.A(KEYINPUT29), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n723), .B1(new_n695), .B2(new_n701), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT29), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n464), .A2(new_n465), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT92), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n548), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n513), .A2(KEYINPUT92), .A3(G179), .A4(new_n518), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n770), .A2(new_n590), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT30), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n637), .A2(new_n774), .ZN(new_n775));
  AND4_X1   g0575(.A1(new_n316), .A2(new_n637), .A3(new_n554), .A4(new_n604), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n773), .A2(new_n775), .B1(new_n508), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n680), .A2(new_n681), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n771), .A2(new_n590), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n778), .A2(new_n779), .A3(new_n770), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n774), .B1(new_n780), .B2(new_n637), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(KEYINPUT31), .B1(new_n782), .B2(new_n733), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(KEYINPUT93), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n509), .A2(new_n505), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n729), .A2(new_n785), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n650), .A2(new_n558), .A3(new_n733), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT31), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n723), .A2(new_n788), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n786), .A2(new_n787), .B1(new_n782), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT93), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n723), .B1(new_n777), .B2(new_n781), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n791), .B1(new_n792), .B2(KEYINPUT31), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n784), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n764), .A2(new_n767), .B1(G330), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n754), .B1(new_n795), .B2(G1), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT95), .ZN(G364));
  INV_X1    g0597(.A(new_n727), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n285), .B1(new_n706), .B2(G45), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n746), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(G330), .B2(new_n726), .ZN(new_n803));
  INV_X1    g0603(.A(new_n256), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n742), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G355), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(G116), .B2(new_n218), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT96), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n742), .A2(new_n256), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n237), .A2(new_n243), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n811), .B(new_n812), .C1(new_n243), .C2(new_n225), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n807), .A2(new_n808), .ZN(new_n814));
  NOR3_X1   g0614(.A1(new_n809), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(G13), .A2(G33), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(G20), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n221), .B1(G20), .B2(new_n299), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n801), .B1(new_n815), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n222), .A2(new_n316), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n823), .A2(G190), .A3(G200), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n824), .A2(KEYINPUT97), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n824), .A2(KEYINPUT97), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(G326), .ZN(new_n829));
  NOR2_X1   g0629(.A1(G190), .A2(G200), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n823), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G311), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n830), .A2(G20), .A3(new_n316), .ZN(new_n833));
  INV_X1    g0633(.A(G329), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n831), .A2(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n823), .ZN(new_n836));
  NOR3_X1   g0636(.A1(new_n836), .A2(new_n587), .A3(G200), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n256), .B(new_n835), .C1(G322), .C2(new_n837), .ZN(new_n838));
  NOR3_X1   g0638(.A1(new_n222), .A2(new_n327), .A3(G179), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(G190), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n839), .A2(new_n587), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n841), .A2(G303), .B1(new_n843), .B2(G283), .ZN(new_n844));
  NOR3_X1   g0644(.A1(new_n836), .A2(G190), .A3(new_n327), .ZN(new_n845));
  XNOR2_X1  g0645(.A(KEYINPUT33), .B(G317), .ZN(new_n846));
  NOR3_X1   g0646(.A1(new_n587), .A2(G179), .A3(G200), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n847), .A2(new_n222), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n845), .A2(new_n846), .B1(new_n849), .B2(G294), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n829), .A2(new_n838), .A3(new_n844), .A4(new_n850), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n576), .A2(new_n840), .B1(new_n842), .B2(new_n312), .ZN(new_n852));
  INV_X1    g0652(.A(new_n837), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n256), .B1(new_n259), .B2(new_n831), .C1(new_n853), .C2(new_n343), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n849), .A2(G97), .ZN(new_n855));
  INV_X1    g0655(.A(new_n845), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n855), .B1(new_n856), .B2(new_n335), .ZN(new_n857));
  INV_X1    g0657(.A(new_n833), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(G159), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT32), .ZN(new_n860));
  OR4_X1    g0660(.A1(new_n852), .A2(new_n854), .A3(new_n857), .A4(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n827), .A2(new_n398), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n851), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OR2_X1    g0663(.A1(new_n863), .A2(KEYINPUT98), .ZN(new_n864));
  INV_X1    g0664(.A(new_n819), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(new_n863), .B2(KEYINPUT98), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n822), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n818), .B(KEYINPUT99), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n867), .B1(new_n726), .B2(new_n868), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n803), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(G396));
  INV_X1    g0671(.A(new_n801), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n794), .A2(G330), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n331), .A2(new_n328), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(new_n733), .B2(new_n325), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT101), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n326), .B(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n723), .B(new_n879), .C1(new_n695), .C2(new_n701), .ZN(new_n880));
  INV_X1    g0680(.A(new_n701), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n733), .B1(new_n881), .B2(new_n759), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n723), .A2(new_n326), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n883), .B1(new_n875), .B2(new_n877), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n880), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n872), .B1(new_n873), .B2(new_n886), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n887), .A2(KEYINPUT102), .B1(new_n873), .B2(new_n886), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(KEYINPUT102), .B2(new_n887), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n865), .A2(new_n817), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n801), .B1(G77), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n831), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n837), .A2(G143), .B1(G159), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(G137), .ZN(new_n894));
  OAI221_X1 g0694(.A(new_n893), .B1(new_n272), .B2(new_n856), .C1(new_n827), .C2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(KEYINPUT34), .ZN(new_n897));
  INV_X1    g0697(.A(G132), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n256), .B1(new_n833), .B2(new_n898), .ZN(new_n899));
  OAI22_X1  g0699(.A1(new_n842), .A2(new_n335), .B1(new_n848), .B2(new_n343), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n899), .B(new_n900), .C1(G50), .C2(new_n841), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n897), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n896), .A2(KEYINPUT34), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n845), .A2(G283), .B1(G116), .B2(new_n892), .ZN(new_n904));
  INV_X1    g0704(.A(G303), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n904), .B1(new_n827), .B2(new_n905), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n906), .B(KEYINPUT100), .Z(new_n907));
  OAI221_X1 g0707(.A(new_n804), .B1(new_n833), .B2(new_n832), .C1(new_n853), .C2(new_n461), .ZN(new_n908));
  OAI221_X1 g0708(.A(new_n855), .B1(new_n840), .B2(new_n312), .C1(new_n576), .C2(new_n842), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI22_X1  g0710(.A1(new_n902), .A2(new_n903), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n891), .B1(new_n911), .B2(new_n819), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n885), .B2(new_n817), .ZN(new_n913));
  AND2_X1   g0713(.A1(new_n889), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(G384));
  AOI21_X1  g0715(.A(new_n444), .B1(new_n766), .B2(new_n765), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n764), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n672), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n918), .B(KEYINPUT107), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT38), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n387), .A2(new_n389), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n362), .A2(new_n719), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n921), .A2(KEYINPUT106), .A3(KEYINPUT37), .A4(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n381), .A2(new_n922), .A3(new_n392), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n730), .B1(new_n359), .B2(new_n361), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT37), .B1(new_n925), .B2(KEYINPUT106), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n922), .B1(new_n653), .B2(new_n670), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n920), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n356), .A2(new_n278), .ZN(new_n931));
  OAI211_X1 g0731(.A(G68), .B(new_n354), .C1(new_n607), .C2(new_n353), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT16), .B1(new_n932), .B2(new_n351), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n361), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n719), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n395), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n934), .A2(new_n380), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n935), .A2(new_n938), .A3(new_n392), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT37), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT37), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n381), .A2(new_n922), .A3(new_n941), .A4(new_n392), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n937), .A2(KEYINPUT38), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n930), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT39), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n666), .A2(new_n723), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT105), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n940), .A2(new_n942), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n935), .B1(new_n653), .B2(new_n670), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n920), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n952), .A2(KEYINPUT39), .A3(new_n944), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n947), .A2(new_n949), .A3(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n409), .B1(new_n720), .B2(new_n722), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT104), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI211_X1 g0757(.A(KEYINPUT104), .B(new_n409), .C1(new_n720), .C2(new_n722), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n664), .B1(new_n658), .B2(new_n659), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n442), .A2(new_n959), .B1(new_n960), .B2(new_n955), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n877), .A2(new_n733), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n962), .B1(new_n880), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n952), .A2(new_n944), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n730), .B1(new_n668), .B2(new_n669), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n954), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n919), .B(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT30), .B1(new_n773), .B2(new_n640), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n778), .A2(new_n779), .A3(new_n770), .A4(new_n775), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n508), .A2(new_n776), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n789), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n558), .A2(new_n733), .ZN(new_n976));
  AND3_X1   g0776(.A1(new_n606), .A2(new_n643), .A3(new_n649), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n975), .B1(new_n978), .B2(new_n510), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n961), .B(new_n885), .C1(new_n979), .C2(new_n783), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT108), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n945), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT40), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n952), .A2(new_n984), .A3(new_n944), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n440), .B1(new_n429), .B2(new_n430), .ZN(new_n986));
  INV_X1    g0786(.A(new_n955), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n658), .A2(new_n659), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n989), .A2(new_n665), .A3(new_n957), .A4(new_n958), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n884), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n976), .A2(new_n977), .A3(new_n685), .A4(new_n506), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n992), .B(new_n975), .C1(KEYINPUT31), .C2(new_n792), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n981), .A2(KEYINPUT40), .ZN(new_n994));
  AND3_X1   g0794(.A1(new_n991), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n983), .A2(KEYINPUT40), .B1(new_n985), .B2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n993), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n996), .B1(new_n444), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n995), .A2(new_n985), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n980), .A2(new_n981), .B1(new_n930), .B2(new_n944), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n999), .B1(new_n1000), .B2(new_n984), .ZN(new_n1001));
  NOR4_X1   g0801(.A1(new_n302), .A2(new_n395), .A3(new_n442), .A4(new_n332), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1001), .A2(new_n1002), .A3(new_n993), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n998), .A2(G330), .A3(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT109), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n970), .A2(new_n1005), .B1(new_n251), .B2(new_n706), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(new_n1005), .B2(new_n970), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n621), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1008), .A2(KEYINPUT35), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(KEYINPUT35), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1009), .A2(new_n1010), .A3(G116), .A4(new_n223), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(KEYINPUT103), .B(KEYINPUT36), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1011), .B(new_n1012), .ZN(new_n1013));
  OR3_X1    g0813(.A1(new_n224), .A2(new_n259), .A3(new_n344), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n201), .A2(G68), .ZN(new_n1015));
  AOI211_X1 g0815(.A(G13), .B(new_n251), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1016));
  OR3_X1    g0816(.A1(new_n1007), .A2(new_n1013), .A3(new_n1016), .ZN(G367));
  OAI221_X1 g0817(.A(new_n820), .B1(new_n218), .B2(new_n319), .C1(new_n811), .C2(new_n233), .ZN(new_n1018));
  AND2_X1   g0818(.A1(new_n1018), .A2(new_n801), .ZN(new_n1019));
  OR3_X1    g0819(.A1(new_n723), .A2(new_n578), .A3(new_n692), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n723), .A2(new_n578), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1020), .B1(new_n755), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n828), .A2(G143), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n201), .A2(new_n831), .B1(new_n833), .B2(new_n894), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n804), .B(new_n1024), .C1(G150), .C2(new_n837), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G159), .A2(new_n845), .B1(new_n843), .B2(G77), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n841), .A2(G58), .B1(new_n849), .B2(G68), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1023), .A2(new_n1025), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(G283), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n853), .A2(new_n905), .B1(new_n831), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G107), .B2(new_n849), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n841), .A2(G116), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT46), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1031), .B(new_n1033), .C1(new_n461), .C2(new_n856), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT111), .ZN(new_n1035));
  INV_X1    g0835(.A(G317), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n804), .B1(new_n1036), .B2(new_n833), .C1(new_n842), .C2(new_n525), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n828), .A2(G311), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1028), .B1(new_n1034), .B2(new_n1039), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT47), .Z(new_n1041));
  OAI221_X1 g0841(.A(new_n1019), .B1(new_n1022), .B2(new_n868), .C1(new_n865), .C2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT44), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n643), .B(new_n649), .C1(new_n723), .C2(new_n626), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n733), .A2(new_n696), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1043), .B1(new_n740), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n738), .A2(new_n739), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1046), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1048), .A2(new_n1049), .A3(KEYINPUT44), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n740), .A2(KEYINPUT45), .A3(new_n1046), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT45), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n1047), .A2(new_n1050), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT110), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n736), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1047), .A2(new_n1050), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1059), .A2(KEYINPUT110), .A3(new_n735), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1056), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n728), .A2(new_n734), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1062), .A2(new_n737), .ZN(new_n1063));
  AND3_X1   g0863(.A1(new_n1063), .A2(new_n727), .A3(new_n738), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n727), .B1(new_n1063), .B2(new_n738), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n795), .B1(new_n1061), .B2(new_n1066), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n746), .B(KEYINPUT41), .Z(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n800), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n786), .A2(new_n737), .A3(new_n1046), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1071), .A2(KEYINPUT42), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n649), .B1(new_n1044), .B2(new_n506), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1071), .A2(KEYINPUT42), .B1(new_n723), .B2(new_n1073), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n1072), .A2(new_n1074), .B1(KEYINPUT43), .B2(new_n1022), .ZN(new_n1075));
  OR3_X1    g0875(.A1(new_n1075), .A2(KEYINPUT43), .A3(new_n1022), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1075), .B1(KEYINPUT43), .B2(new_n1022), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n735), .A2(new_n1046), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1076), .A2(new_n735), .A3(new_n1046), .A4(new_n1077), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1042), .B1(new_n1070), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(KEYINPUT112), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT112), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1085), .B(new_n1042), .C1(new_n1070), .C2(new_n1082), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n1084), .A2(new_n1086), .ZN(G387));
  INV_X1    g0887(.A(new_n1066), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n1062), .A2(new_n868), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n837), .A2(G317), .B1(G303), .B2(new_n892), .ZN(new_n1090));
  INV_X1    g0890(.A(G322), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n1090), .B1(new_n832), .B2(new_n856), .C1(new_n827), .C2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT48), .ZN(new_n1093));
  OR2_X1    g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n841), .A2(G294), .B1(new_n849), .B2(G283), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT49), .ZN(new_n1098));
  OR2_X1    g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n842), .A2(new_n521), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n256), .B(new_n1101), .C1(G326), .C2(new_n858), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1099), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n853), .A2(new_n398), .B1(new_n831), .B2(new_n335), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n804), .B(new_n1104), .C1(G150), .C2(new_n858), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n828), .A2(G159), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n840), .A2(new_n259), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(G97), .B2(new_n843), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n270), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1109), .A2(new_n845), .B1(new_n849), .B2(new_n574), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1105), .A2(new_n1106), .A3(new_n1108), .A4(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n865), .B1(new_n1103), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n230), .A2(G45), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT114), .ZN(new_n1116));
  AOI21_X1  g0916(.A(KEYINPUT50), .B1(new_n1109), .B2(new_n398), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n1109), .A2(KEYINPUT50), .A3(new_n398), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n1115), .B1(new_n749), .B2(new_n1116), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n750), .A2(KEYINPUT114), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n810), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT115), .ZN(new_n1122));
  OR2_X1    g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1114), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n805), .A2(new_n749), .B1(new_n312), .B2(new_n742), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n821), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NOR3_X1   g0927(.A1(new_n1112), .A2(new_n872), .A3(new_n1127), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n1088), .A2(new_n800), .B1(new_n1089), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1088), .A2(new_n795), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n746), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1088), .A2(new_n795), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1129), .B1(new_n1131), .B2(new_n1132), .ZN(G393));
  XNOR2_X1  g0933(.A(new_n1059), .B(new_n735), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n1134), .A2(new_n799), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n820), .B1(new_n525), .B2(new_n218), .C1(new_n811), .C2(new_n240), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1136), .A2(new_n801), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n818), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n828), .A2(G150), .B1(G159), .B2(new_n837), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT51), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n804), .B1(new_n858), .B2(G143), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n270), .B2(new_n831), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n335), .A2(new_n840), .B1(new_n842), .B2(new_n576), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n856), .A2(new_n201), .B1(new_n259), .B2(new_n848), .ZN(new_n1144));
  NOR4_X1   g0944(.A1(new_n1140), .A2(new_n1142), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n827), .A2(new_n1036), .B1(new_n832), .B2(new_n853), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT52), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n856), .A2(new_n905), .B1(new_n312), .B2(new_n842), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n804), .B1(new_n833), .B2(new_n1091), .C1(new_n831), .C2(new_n461), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n840), .A2(new_n1029), .B1(new_n848), .B2(new_n521), .ZN(new_n1150));
  NOR3_X1   g0950(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1145), .B1(new_n1147), .B2(new_n1151), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1137), .B1(new_n1046), .B2(new_n1138), .C1(new_n1152), .C2(new_n865), .ZN(new_n1153));
  OR2_X1    g0953(.A1(new_n1130), .A2(new_n1061), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n746), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1130), .A2(new_n1134), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1135), .B(new_n1153), .C1(new_n1155), .C2(new_n1157), .ZN(G390));
  NAND2_X1  g0958(.A1(new_n947), .A2(new_n953), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n816), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n801), .B1(new_n1109), .B2(new_n890), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n853), .A2(new_n521), .B1(new_n831), .B2(new_n525), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n256), .B(new_n1162), .C1(G294), .C2(new_n858), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n828), .A2(G283), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n841), .A2(G87), .B1(new_n843), .B2(G68), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(G107), .A2(new_n845), .B1(new_n849), .B2(G77), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(G137), .A2(new_n845), .B1(new_n849), .B2(G159), .ZN(new_n1168));
  XOR2_X1   g0968(.A(KEYINPUT54), .B(G143), .Z(new_n1169));
  AOI22_X1  g0969(.A1(new_n837), .A2(G132), .B1(new_n892), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n804), .B1(new_n858), .B2(G125), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n843), .A2(new_n202), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1168), .A2(new_n1170), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n840), .A2(new_n272), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT53), .ZN(new_n1175));
  INV_X1    g0975(.A(G128), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1175), .B1(new_n1176), .B2(new_n827), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1167), .B1(new_n1173), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1161), .B1(new_n1178), .B2(new_n819), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1160), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n953), .ZN(new_n1181));
  AOI21_X1  g0981(.A(KEYINPUT39), .B1(new_n930), .B2(new_n944), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n1181), .A2(new_n1182), .B1(new_n965), .B2(new_n949), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n794), .A2(G330), .A3(new_n885), .A4(new_n961), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT116), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n961), .B(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n885), .B1(new_n761), .B2(new_n763), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1186), .B1(new_n1187), .B2(new_n964), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n949), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n945), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1183), .B(new_n1184), .C1(new_n1188), .C2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1186), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n756), .A2(new_n692), .A3(new_n757), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n785), .A2(new_n693), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1193), .B1(new_n676), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n762), .B1(new_n1195), .B2(new_n733), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n760), .A2(KEYINPUT94), .A3(new_n723), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n884), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1192), .B1(new_n1198), .B2(new_n963), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1190), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n963), .B1(new_n882), .B2(new_n879), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1189), .B1(new_n1201), .B2(new_n962), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1199), .A2(new_n1200), .B1(new_n1159), .B2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(G330), .B1(new_n979), .B2(new_n783), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n961), .A2(new_n885), .ZN(new_n1205));
  OAI21_X1  g1005(.A(KEYINPUT117), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT117), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n991), .A2(new_n993), .A3(new_n1207), .A4(G330), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n1206), .A2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1191), .B1(new_n1203), .B2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1180), .B1(new_n1210), .B2(new_n799), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1002), .A2(G330), .A3(new_n993), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n766), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n767), .A2(new_n1002), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n672), .B(new_n1212), .C1(new_n1213), .C2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT118), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n917), .A2(KEYINPUT118), .A3(new_n672), .A4(new_n1212), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n962), .B1(new_n873), .B2(new_n884), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1201), .B1(new_n1209), .B2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n993), .A2(G330), .A3(new_n885), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1186), .A2(new_n1221), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1222), .A2(new_n1187), .A3(new_n1184), .A4(new_n964), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1217), .B(new_n1218), .C1(new_n1220), .C2(new_n1224), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n1210), .A2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n747), .B1(new_n1210), .B2(new_n1225), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1211), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(G378));
  AND2_X1   g1029(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1220), .A2(new_n1224), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1230), .B1(new_n1210), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(G330), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n302), .A2(new_n292), .A3(new_n719), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n297), .B(new_n301), .C1(new_n290), .C2(new_n730), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1236));
  AND3_X1   g1036(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1236), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n930), .A2(new_n944), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT108), .B1(new_n991), .B2(new_n993), .ZN(new_n1241));
  OAI21_X1  g1041(.A(KEYINPUT40), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1233), .B(new_n1239), .C1(new_n1242), .C2(new_n999), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1239), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(new_n1001), .B2(G330), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n969), .B1(new_n1243), .B2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1239), .B1(new_n996), .B2(new_n1233), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n969), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1001), .A2(G330), .A3(new_n1244), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1246), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1232), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT57), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n747), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1253), .B1(new_n1246), .B2(new_n1250), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1232), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(KEYINPUT120), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT120), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1255), .A2(new_n1258), .A3(new_n1232), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1254), .A2(new_n1257), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1239), .A2(new_n816), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n801), .B1(new_n202), .B2(new_n890), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n856), .A2(new_n525), .B1(new_n343), .B2(new_n842), .ZN(new_n1263));
  AOI211_X1 g1063(.A(new_n1107), .B(new_n1263), .C1(G68), .C2(new_n849), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n804), .A2(new_n242), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n831), .A2(new_n319), .B1(new_n833), .B2(new_n1029), .ZN(new_n1266));
  AOI211_X1 g1066(.A(new_n1265), .B(new_n1266), .C1(G107), .C2(new_n837), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1264), .B(new_n1267), .C1(new_n521), .C2(new_n827), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT58), .ZN(new_n1269));
  AOI21_X1  g1069(.A(G50), .B1(new_n273), .B2(new_n242), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n1268), .A2(new_n1269), .B1(new_n1265), .B2(new_n1270), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n853), .A2(new_n1176), .B1(new_n831), .B2(new_n894), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(G150), .B2(new_n849), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n841), .A2(new_n1169), .ZN(new_n1274));
  XOR2_X1   g1074(.A(new_n1274), .B(KEYINPUT119), .Z(new_n1275));
  NAND2_X1  g1075(.A1(new_n828), .A2(G125), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n845), .A2(G132), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1273), .A2(new_n1275), .A3(new_n1276), .A4(new_n1277), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1278), .A2(KEYINPUT59), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(KEYINPUT59), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n843), .A2(G159), .ZN(new_n1281));
  AOI211_X1 g1081(.A(G33), .B(G41), .C1(new_n858), .C2(G124), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1280), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  OAI221_X1 g1083(.A(new_n1271), .B1(new_n1269), .B2(new_n1268), .C1(new_n1279), .C2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1262), .B1(new_n1284), .B2(new_n819), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(new_n1251), .A2(new_n800), .B1(new_n1261), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1260), .A2(new_n1286), .ZN(G375));
  OR3_X1    g1087(.A1(new_n1231), .A2(KEYINPUT121), .A3(new_n799), .ZN(new_n1288));
  OAI21_X1  g1088(.A(KEYINPUT121), .B1(new_n1231), .B2(new_n799), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n828), .A2(G132), .ZN(new_n1290));
  OAI22_X1  g1090(.A1(new_n831), .A2(new_n272), .B1(new_n833), .B2(new_n1176), .ZN(new_n1291));
  AOI211_X1 g1091(.A(new_n804), .B(new_n1291), .C1(G137), .C2(new_n837), .ZN(new_n1292));
  AOI22_X1  g1092(.A1(new_n845), .A2(new_n1169), .B1(new_n843), .B2(G58), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(new_n841), .A2(G159), .B1(new_n849), .B2(G50), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1290), .A2(new_n1292), .A3(new_n1293), .A4(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n804), .B1(new_n842), .B2(new_n259), .ZN(new_n1296));
  XOR2_X1   g1096(.A(new_n1296), .B(KEYINPUT122), .Z(new_n1297));
  OAI22_X1  g1097(.A1(new_n831), .A2(new_n312), .B1(new_n833), .B2(new_n905), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n840), .A2(new_n525), .ZN(new_n1299));
  AOI211_X1 g1099(.A(new_n1298), .B(new_n1299), .C1(G116), .C2(new_n845), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n1297), .B(new_n1300), .C1(new_n461), .C2(new_n827), .ZN(new_n1301));
  AOI22_X1  g1101(.A1(G283), .A2(new_n837), .B1(new_n849), .B2(new_n574), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(new_n1302), .B(KEYINPUT123), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1295), .B1(new_n1301), .B2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT124), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n865), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1306), .B1(new_n1305), .B2(new_n1304), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n801), .B1(G68), .B2(new_n890), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  OAI211_X1 g1109(.A(new_n1307), .B(new_n1309), .C1(new_n1192), .C2(new_n817), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1288), .A2(new_n1289), .A3(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1225), .A2(new_n1069), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1209), .A2(new_n1219), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1201), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1223), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1230), .A2(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1312), .B1(new_n1313), .B2(new_n1318), .ZN(G381));
  OR4_X1    g1119(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1320));
  NOR3_X1   g1120(.A1(new_n1320), .A2(G387), .A3(G381), .ZN(new_n1321));
  XOR2_X1   g1121(.A(new_n1321), .B(KEYINPUT125), .Z(new_n1322));
  INV_X1    g1122(.A(new_n1286), .ZN(new_n1323));
  AND3_X1   g1123(.A1(new_n1255), .A2(new_n1258), .A3(new_n1232), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1258), .B1(new_n1255), .B2(new_n1232), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1323), .B1(new_n1326), .B2(new_n1254), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(new_n1228), .ZN(new_n1328));
  OR2_X1    g1128(.A1(new_n1322), .A2(new_n1328), .ZN(G407));
  NAND3_X1  g1129(.A1(new_n1327), .A2(new_n721), .A3(new_n1228), .ZN(new_n1330));
  OAI211_X1 g1130(.A(G213), .B(new_n1330), .C1(new_n1322), .C2(new_n1328), .ZN(G409));
  NAND3_X1  g1131(.A1(new_n1232), .A2(new_n1251), .A3(new_n1069), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1228), .A2(new_n1286), .A3(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n721), .A2(G213), .ZN(new_n1334));
  AND2_X1   g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1335), .B1(new_n1327), .B2(new_n1228), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT126), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1225), .A2(new_n746), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1339));
  AOI21_X1  g1139(.A(KEYINPUT60), .B1(new_n1231), .B2(new_n1339), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1338), .A2(new_n1340), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1231), .A2(new_n1339), .A3(KEYINPUT60), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1337), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT60), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1344), .B1(new_n1230), .B2(new_n1317), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n747), .B1(new_n1230), .B2(new_n1317), .ZN(new_n1346));
  NAND4_X1  g1146(.A1(new_n1345), .A2(new_n1346), .A3(new_n1337), .A4(new_n1342), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1347), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1312), .B1(new_n1343), .B2(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1349), .A2(new_n914), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1345), .A2(new_n1346), .A3(new_n1342), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1351), .A2(KEYINPUT126), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1352), .A2(new_n1347), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1353), .A2(G384), .A3(new_n1312), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1350), .A2(new_n1354), .ZN(new_n1355));
  OAI21_X1  g1155(.A(KEYINPUT62), .B1(new_n1336), .B2(new_n1355), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n721), .A2(G213), .A3(G2897), .ZN(new_n1357));
  INV_X1    g1157(.A(new_n1357), .ZN(new_n1358));
  AOI21_X1  g1158(.A(G384), .B1(new_n1353), .B2(new_n1312), .ZN(new_n1359));
  AOI211_X1 g1159(.A(new_n914), .B(new_n1311), .C1(new_n1352), .C2(new_n1347), .ZN(new_n1360));
  OAI21_X1  g1160(.A(new_n1358), .B1(new_n1359), .B2(new_n1360), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1350), .A2(new_n1354), .A3(new_n1357), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1336), .A2(new_n1361), .A3(new_n1362), .ZN(new_n1363));
  INV_X1    g1163(.A(KEYINPUT61), .ZN(new_n1364));
  NOR2_X1   g1164(.A1(new_n1359), .A2(new_n1360), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(G375), .A2(G378), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT62), .ZN(new_n1367));
  NAND4_X1  g1167(.A1(new_n1365), .A2(new_n1366), .A3(new_n1367), .A4(new_n1335), .ZN(new_n1368));
  NAND4_X1  g1168(.A1(new_n1356), .A2(new_n1363), .A3(new_n1364), .A4(new_n1368), .ZN(new_n1369));
  XNOR2_X1  g1169(.A(G393), .B(G396), .ZN(new_n1370));
  OAI211_X1 g1170(.A(G390), .B(new_n1042), .C1(new_n1070), .C2(new_n1082), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1135), .A2(new_n1153), .ZN(new_n1372));
  INV_X1    g1172(.A(new_n1155), .ZN(new_n1373));
  AOI21_X1  g1173(.A(new_n1372), .B1(new_n1373), .B2(new_n1156), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1374), .A2(new_n1083), .ZN(new_n1375));
  AOI21_X1  g1175(.A(new_n1370), .B1(new_n1371), .B2(new_n1375), .ZN(new_n1376));
  NAND3_X1  g1176(.A1(new_n1084), .A2(new_n1374), .A3(new_n1086), .ZN(new_n1377));
  INV_X1    g1177(.A(KEYINPUT127), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1377), .A2(new_n1378), .ZN(new_n1379));
  NAND4_X1  g1179(.A1(new_n1084), .A2(new_n1374), .A3(KEYINPUT127), .A4(new_n1086), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1379), .A2(new_n1380), .ZN(new_n1381));
  AND2_X1   g1181(.A1(new_n1371), .A2(new_n1370), .ZN(new_n1382));
  AOI21_X1  g1182(.A(new_n1376), .B1(new_n1381), .B2(new_n1382), .ZN(new_n1383));
  NAND2_X1  g1183(.A1(new_n1369), .A2(new_n1383), .ZN(new_n1384));
  NAND3_X1  g1184(.A1(new_n1365), .A2(new_n1366), .A3(new_n1335), .ZN(new_n1385));
  INV_X1    g1185(.A(KEYINPUT63), .ZN(new_n1386));
  AOI21_X1  g1186(.A(new_n1383), .B1(new_n1385), .B2(new_n1386), .ZN(new_n1387));
  NAND4_X1  g1187(.A1(new_n1365), .A2(new_n1366), .A3(KEYINPUT63), .A4(new_n1335), .ZN(new_n1388));
  NAND4_X1  g1188(.A1(new_n1387), .A2(new_n1364), .A3(new_n1363), .A4(new_n1388), .ZN(new_n1389));
  NAND2_X1  g1189(.A1(new_n1384), .A2(new_n1389), .ZN(G405));
  NAND2_X1  g1190(.A1(new_n1328), .A2(new_n1366), .ZN(new_n1391));
  NAND2_X1  g1191(.A1(new_n1391), .A2(new_n1365), .ZN(new_n1392));
  NAND3_X1  g1192(.A1(new_n1355), .A2(new_n1328), .A3(new_n1366), .ZN(new_n1393));
  NAND2_X1  g1193(.A1(new_n1392), .A2(new_n1393), .ZN(new_n1394));
  AND2_X1   g1194(.A1(new_n1381), .A2(new_n1382), .ZN(new_n1395));
  OAI21_X1  g1195(.A(new_n1394), .B1(new_n1376), .B2(new_n1395), .ZN(new_n1396));
  NAND3_X1  g1196(.A1(new_n1392), .A2(new_n1383), .A3(new_n1393), .ZN(new_n1397));
  NAND2_X1  g1197(.A1(new_n1396), .A2(new_n1397), .ZN(G402));
endmodule


