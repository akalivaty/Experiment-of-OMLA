

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732;

  XNOR2_X1 U368 ( .A(n346), .B(n418), .ZN(n656) );
  NOR2_X1 U369 ( .A1(n558), .A2(n559), .ZN(n405) );
  AND2_X2 U370 ( .A1(n364), .A2(n362), .ZN(n359) );
  XNOR2_X2 U371 ( .A(n715), .B(G146), .ZN(n523) );
  XNOR2_X2 U372 ( .A(n505), .B(n462), .ZN(n715) );
  XNOR2_X2 U373 ( .A(n385), .B(n384), .ZN(n465) );
  NOR2_X1 U374 ( .A1(n728), .A2(n729), .ZN(n420) );
  NOR2_X2 U375 ( .A1(n661), .A2(n659), .ZN(n540) );
  BUF_X1 U376 ( .A(n359), .Z(n698) );
  NOR2_X1 U377 ( .A1(n595), .A2(n588), .ZN(n571) );
  NAND2_X1 U378 ( .A1(n535), .A2(n579), .ZN(n595) );
  INV_X1 U379 ( .A(KEYINPUT45), .ZN(n604) );
  NOR2_X1 U380 ( .A1(n726), .A2(n445), .ZN(n602) );
  AND2_X1 U381 ( .A1(n398), .A2(n397), .ZN(n561) );
  XNOR2_X1 U382 ( .A(n396), .B(KEYINPUT40), .ZN(n730) );
  XNOR2_X1 U383 ( .A(n405), .B(KEYINPUT77), .ZN(n629) );
  XNOR2_X1 U384 ( .A(n571), .B(KEYINPUT33), .ZN(n672) );
  NOR2_X1 U385 ( .A1(n581), .A2(n541), .ZN(n542) );
  XNOR2_X1 U386 ( .A(n399), .B(KEYINPUT105), .ZN(n619) );
  OR2_X1 U387 ( .A1(n556), .A2(n557), .ZN(n399) );
  XNOR2_X1 U388 ( .A(n534), .B(n426), .ZN(n579) );
  XNOR2_X1 U389 ( .A(n436), .B(n713), .ZN(n697) );
  XOR2_X1 U390 ( .A(n689), .B(KEYINPUT59), .Z(n691) );
  XNOR2_X1 U391 ( .A(n439), .B(n437), .ZN(n436) );
  XOR2_X1 U392 ( .A(G146), .B(G125), .Z(n473) );
  BUF_X1 U393 ( .A(n390), .Z(n346) );
  XNOR2_X1 U394 ( .A(n358), .B(n459), .ZN(n390) );
  NOR2_X1 U395 ( .A1(n370), .A2(n369), .ZN(n368) );
  XNOR2_X1 U396 ( .A(n376), .B(KEYINPUT82), .ZN(n677) );
  XOR2_X1 U397 ( .A(KEYINPUT4), .B(G131), .Z(n462) );
  XNOR2_X1 U398 ( .A(n430), .B(KEYINPUT68), .ZN(n475) );
  INV_X1 U399 ( .A(G137), .ZN(n430) );
  XNOR2_X1 U400 ( .A(n454), .B(n413), .ZN(n412) );
  XNOR2_X1 U401 ( .A(n449), .B(n414), .ZN(n413) );
  XNOR2_X1 U402 ( .A(n452), .B(n403), .ZN(n454) );
  XNOR2_X1 U403 ( .A(n503), .B(n434), .ZN(n713) );
  INV_X1 U404 ( .A(n475), .ZN(n434) );
  INV_X1 U405 ( .A(G110), .ZN(n384) );
  XNOR2_X1 U406 ( .A(G137), .B(G116), .ZN(n516) );
  XOR2_X1 U407 ( .A(KEYINPUT5), .B(KEYINPUT98), .Z(n517) );
  INV_X1 U408 ( .A(n677), .ZN(n360) );
  INV_X1 U409 ( .A(n682), .ZN(n362) );
  XNOR2_X1 U410 ( .A(n415), .B(n354), .ZN(n377) );
  INV_X1 U411 ( .A(KEYINPUT38), .ZN(n418) );
  OR2_X1 U412 ( .A1(G237), .A2(G902), .ZN(n527) );
  NOR2_X1 U413 ( .A1(G902), .A2(n612), .ZN(n524) );
  XNOR2_X1 U414 ( .A(n388), .B(n448), .ZN(n521) );
  XNOR2_X1 U415 ( .A(n447), .B(n446), .ZN(n388) );
  INV_X1 U416 ( .A(KEYINPUT3), .ZN(n446) );
  XNOR2_X1 U417 ( .A(G119), .B(G128), .ZN(n481) );
  XOR2_X1 U418 ( .A(KEYINPUT96), .B(G110), .Z(n482) );
  INV_X1 U419 ( .A(KEYINPUT23), .ZN(n438) );
  XNOR2_X1 U420 ( .A(n387), .B(n386), .ZN(n513) );
  XNOR2_X1 U421 ( .A(G116), .B(G107), .ZN(n387) );
  XNOR2_X1 U422 ( .A(n435), .B(n473), .ZN(n503) );
  XNOR2_X1 U423 ( .A(n474), .B(G140), .ZN(n435) );
  XOR2_X1 U424 ( .A(KEYINPUT67), .B(KEYINPUT10), .Z(n474) );
  AND2_X1 U425 ( .A1(n374), .A2(n577), .ZN(n531) );
  AND2_X1 U426 ( .A1(n619), .A2(n375), .ZN(n374) );
  INV_X1 U427 ( .A(n541), .ZN(n375) );
  XNOR2_X1 U428 ( .A(n531), .B(n373), .ZN(n372) );
  INV_X1 U429 ( .A(KEYINPUT113), .ZN(n373) );
  AND2_X1 U430 ( .A1(n576), .A2(n394), .ZN(n422) );
  INV_X1 U431 ( .A(KEYINPUT1), .ZN(n426) );
  NOR2_X1 U432 ( .A1(n697), .A2(G902), .ZN(n488) );
  XNOR2_X1 U433 ( .A(n429), .B(n427), .ZN(n466) );
  XNOR2_X1 U434 ( .A(n464), .B(n428), .ZN(n427) );
  NOR2_X1 U435 ( .A1(G952), .A2(n720), .ZN(n702) );
  NOR2_X1 U436 ( .A1(n681), .A2(n682), .ZN(n381) );
  NOR2_X1 U437 ( .A1(n662), .A2(n629), .ZN(n560) );
  XNOR2_X1 U438 ( .A(n453), .B(n404), .ZN(n403) );
  INV_X1 U439 ( .A(KEYINPUT90), .ZN(n404) );
  INV_X1 U440 ( .A(n473), .ZN(n414) );
  INV_X1 U441 ( .A(n461), .ZN(n449) );
  XNOR2_X1 U442 ( .A(G101), .B(G113), .ZN(n447) );
  INV_X1 U443 ( .A(G134), .ZN(n460) );
  NAND2_X1 U444 ( .A1(G234), .A2(G237), .ZN(n489) );
  NAND2_X1 U445 ( .A1(n656), .A2(n655), .ZN(n661) );
  XNOR2_X1 U446 ( .A(G902), .B(KEYINPUT15), .ZN(n457) );
  NOR2_X1 U447 ( .A1(n348), .A2(n655), .ZN(n369) );
  XNOR2_X1 U448 ( .A(n401), .B(n504), .ZN(n549) );
  XNOR2_X1 U449 ( .A(n468), .B(G469), .ZN(n534) );
  XNOR2_X1 U450 ( .A(n523), .B(n522), .ZN(n612) );
  BUF_X1 U451 ( .A(n677), .Z(n716) );
  XNOR2_X1 U452 ( .A(KEYINPUT103), .B(KEYINPUT102), .ZN(n506) );
  XOR2_X1 U453 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n507) );
  XNOR2_X1 U454 ( .A(G131), .B(KEYINPUT12), .ZN(n497) );
  NOR2_X1 U455 ( .A1(G953), .A2(G237), .ZN(n518) );
  XNOR2_X1 U456 ( .A(KEYINPUT73), .B(G140), .ZN(n428) );
  XNOR2_X1 U457 ( .A(n475), .B(n463), .ZN(n429) );
  AND2_X1 U458 ( .A1(n363), .A2(n609), .ZN(n682) );
  AND2_X1 U459 ( .A1(n377), .A2(n389), .ZN(n609) );
  XNOR2_X1 U460 ( .A(n431), .B(KEYINPUT39), .ZN(n563) );
  NAND2_X1 U461 ( .A1(n432), .A2(n552), .ZN(n431) );
  AND2_X1 U462 ( .A1(n656), .A2(n550), .ZN(n433) );
  XNOR2_X1 U463 ( .A(n393), .B(n392), .ZN(n425) );
  INV_X1 U464 ( .A(KEYINPUT34), .ZN(n392) );
  BUF_X1 U465 ( .A(n575), .Z(n596) );
  XNOR2_X1 U466 ( .A(n408), .B(n407), .ZN(n515) );
  INV_X1 U467 ( .A(G478), .ZN(n407) );
  XNOR2_X1 U468 ( .A(n596), .B(KEYINPUT93), .ZN(n411) );
  XNOR2_X1 U469 ( .A(n383), .B(n513), .ZN(n382) );
  XNOR2_X1 U470 ( .A(n465), .B(KEYINPUT16), .ZN(n383) );
  XNOR2_X1 U471 ( .A(n477), .B(n438), .ZN(n437) );
  XNOR2_X1 U472 ( .A(n480), .B(n483), .ZN(n439) );
  INV_X1 U473 ( .A(n702), .ZN(n441) );
  XNOR2_X1 U474 ( .A(n400), .B(KEYINPUT36), .ZN(n532) );
  XNOR2_X1 U475 ( .A(n694), .B(n391), .ZN(n696) );
  XNOR2_X1 U476 ( .A(n695), .B(KEYINPUT122), .ZN(n391) );
  XNOR2_X1 U477 ( .A(n687), .B(n686), .ZN(n688) );
  INV_X1 U478 ( .A(KEYINPUT53), .ZN(n378) );
  AND2_X1 U479 ( .A1(n683), .A2(n720), .ZN(n406) );
  NAND2_X1 U480 ( .A1(n646), .A2(n579), .ZN(n347) );
  XNOR2_X1 U481 ( .A(KEYINPUT71), .B(KEYINPUT19), .ZN(n348) );
  INV_X1 U482 ( .A(n579), .ZN(n642) );
  XNOR2_X1 U483 ( .A(KEYINPUT78), .B(n608), .ZN(n349) );
  XOR2_X1 U484 ( .A(G113), .B(G143), .Z(n350) );
  INV_X1 U485 ( .A(n389), .ZN(n640) );
  OR2_X1 U486 ( .A1(n577), .A2(n347), .ZN(n351) );
  AND2_X1 U487 ( .A1(n389), .A2(n639), .ZN(n352) );
  XNOR2_X1 U488 ( .A(n574), .B(KEYINPUT75), .ZN(n353) );
  XOR2_X1 U489 ( .A(KEYINPUT48), .B(KEYINPUT84), .Z(n354) );
  XOR2_X1 U490 ( .A(n546), .B(KEYINPUT85), .Z(n355) );
  XNOR2_X1 U491 ( .A(n382), .B(n521), .ZN(n703) );
  OR2_X1 U492 ( .A1(n678), .A2(n607), .ZN(n356) );
  XOR2_X1 U493 ( .A(n611), .B(KEYINPUT56), .Z(n357) );
  NOR2_X1 U494 ( .A1(n458), .A2(n469), .ZN(n358) );
  NAND2_X1 U495 ( .A1(n365), .A2(n356), .ZN(n364) );
  INV_X1 U496 ( .A(n536), .ZN(n581) );
  INV_X1 U497 ( .A(n644), .ZN(n592) );
  NAND2_X1 U498 ( .A1(n361), .A2(n360), .ZN(n365) );
  XNOR2_X1 U499 ( .A(n606), .B(KEYINPUT80), .ZN(n361) );
  NOR2_X1 U500 ( .A1(n705), .A2(n349), .ZN(n363) );
  AND2_X1 U501 ( .A1(n346), .A2(n655), .ZN(n371) );
  NAND2_X1 U502 ( .A1(n368), .A2(n366), .ZN(n569) );
  NAND2_X1 U503 ( .A1(n390), .A2(n367), .ZN(n366) );
  AND2_X1 U504 ( .A1(n655), .A2(n348), .ZN(n367) );
  NOR2_X1 U505 ( .A1(n390), .A2(n348), .ZN(n370) );
  XNOR2_X2 U506 ( .A(n461), .B(n460), .ZN(n505) );
  NAND2_X1 U507 ( .A1(n372), .A2(n371), .ZN(n400) );
  NAND2_X1 U508 ( .A1(n377), .A2(n352), .ZN(n376) );
  XNOR2_X1 U509 ( .A(n379), .B(n378), .ZN(G75) );
  NAND2_X1 U510 ( .A1(n380), .A2(n406), .ZN(n379) );
  XNOR2_X1 U511 ( .A(n381), .B(KEYINPUT81), .ZN(n380) );
  XNOR2_X2 U512 ( .A(G104), .B(KEYINPUT89), .ZN(n385) );
  INV_X1 U513 ( .A(G122), .ZN(n386) );
  NAND2_X1 U514 ( .A1(n554), .A2(n346), .ZN(n555) );
  OR2_X1 U515 ( .A1(n530), .A2(n346), .ZN(n389) );
  XNOR2_X1 U516 ( .A(n613), .B(n614), .ZN(n615) );
  NAND2_X1 U517 ( .A1(n410), .A2(n411), .ZN(n393) );
  AND2_X1 U518 ( .A1(n646), .A2(n394), .ZN(n495) );
  INV_X1 U519 ( .A(n647), .ZN(n394) );
  XNOR2_X2 U520 ( .A(n488), .B(n487), .ZN(n646) );
  XNOR2_X1 U521 ( .A(n421), .B(KEYINPUT22), .ZN(n580) );
  NAND2_X1 U522 ( .A1(n395), .A2(n586), .ZN(n603) );
  NAND2_X1 U523 ( .A1(n419), .A2(n409), .ZN(n395) );
  XNOR2_X1 U524 ( .A(n690), .B(n691), .ZN(n692) );
  NAND2_X1 U525 ( .A1(n423), .A2(n422), .ZN(n421) );
  NAND2_X1 U526 ( .A1(n359), .A2(G472), .ZN(n613) );
  NAND2_X1 U527 ( .A1(n563), .A2(n619), .ZN(n396) );
  XNOR2_X2 U528 ( .A(n592), .B(KEYINPUT108), .ZN(n536) );
  XNOR2_X1 U529 ( .A(n703), .B(n412), .ZN(n458) );
  NOR2_X2 U530 ( .A1(n615), .A2(n702), .ZN(n618) );
  XNOR2_X1 U531 ( .A(n420), .B(n585), .ZN(n419) );
  INV_X1 U532 ( .A(n628), .ZN(n397) );
  XNOR2_X1 U533 ( .A(n560), .B(KEYINPUT47), .ZN(n398) );
  AND2_X1 U534 ( .A1(n551), .A2(n433), .ZN(n432) );
  NOR2_X2 U535 ( .A1(n580), .A2(n579), .ZN(n587) );
  NOR2_X1 U536 ( .A1(n689), .A2(G902), .ZN(n401) );
  XNOR2_X1 U537 ( .A(n402), .B(n499), .ZN(n501) );
  XNOR2_X1 U538 ( .A(n496), .B(n350), .ZN(n402) );
  NOR2_X2 U539 ( .A1(n705), .A2(n607), .ZN(n606) );
  NOR2_X1 U540 ( .A1(n695), .A2(G902), .ZN(n408) );
  NOR2_X1 U541 ( .A1(n548), .A2(n637), .ZN(n417) );
  NAND2_X1 U542 ( .A1(n417), .A2(n416), .ZN(n415) );
  INV_X1 U543 ( .A(n672), .ZN(n410) );
  INV_X1 U544 ( .A(n725), .ZN(n409) );
  XNOR2_X2 U545 ( .A(n424), .B(n353), .ZN(n725) );
  NAND2_X1 U546 ( .A1(n411), .A2(n535), .ZN(n591) );
  XNOR2_X1 U547 ( .A(n561), .B(KEYINPUT70), .ZN(n416) );
  INV_X1 U548 ( .A(n575), .ZN(n423) );
  NAND2_X1 U549 ( .A1(n425), .A2(n573), .ZN(n424) );
  XNOR2_X1 U550 ( .A(n440), .B(n357), .ZN(G51) );
  NAND2_X1 U551 ( .A1(n442), .A2(n441), .ZN(n440) );
  XNOR2_X1 U552 ( .A(n443), .B(n610), .ZN(n442) );
  NAND2_X1 U553 ( .A1(n359), .A2(G210), .ZN(n443) );
  INV_X1 U554 ( .A(n596), .ZN(n597) );
  AND2_X1 U555 ( .A1(n518), .A2(G210), .ZN(n444) );
  AND2_X1 U556 ( .A1(n601), .A2(n600), .ZN(n445) );
  XNOR2_X1 U557 ( .A(n519), .B(n444), .ZN(n520) );
  XNOR2_X1 U558 ( .A(n570), .B(KEYINPUT0), .ZN(n575) );
  XNOR2_X1 U559 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U560 ( .A(n465), .B(n466), .ZN(n467) );
  INV_X1 U561 ( .A(n569), .ZN(n559) );
  XNOR2_X1 U562 ( .A(n523), .B(n467), .ZN(n685) );
  XNOR2_X1 U563 ( .A(n685), .B(n684), .ZN(n686) );
  XNOR2_X1 U564 ( .A(n616), .B(KEYINPUT63), .ZN(n617) );
  XNOR2_X1 U565 ( .A(n618), .B(n617), .ZN(G57) );
  INV_X2 U566 ( .A(G953), .ZN(n720) );
  XOR2_X1 U567 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n456) );
  XOR2_X1 U568 ( .A(KEYINPUT69), .B(G119), .Z(n448) );
  XOR2_X2 U569 ( .A(G143), .B(G128), .Z(n461) );
  XOR2_X1 U570 ( .A(KEYINPUT17), .B(KEYINPUT74), .Z(n451) );
  XNOR2_X1 U571 ( .A(KEYINPUT4), .B(KEYINPUT18), .ZN(n450) );
  XNOR2_X1 U572 ( .A(n451), .B(n450), .ZN(n452) );
  NAND2_X1 U573 ( .A1(G224), .A2(n720), .ZN(n453) );
  XNOR2_X1 U574 ( .A(n458), .B(KEYINPUT87), .ZN(n455) );
  XNOR2_X1 U575 ( .A(n456), .B(n455), .ZN(n610) );
  XOR2_X1 U576 ( .A(n457), .B(KEYINPUT88), .Z(n469) );
  NAND2_X1 U577 ( .A1(G210), .A2(n527), .ZN(n459) );
  XNOR2_X1 U578 ( .A(G101), .B(G107), .ZN(n463) );
  NAND2_X1 U579 ( .A1(G227), .A2(n720), .ZN(n464) );
  NOR2_X1 U580 ( .A1(G902), .A2(n685), .ZN(n468) );
  XOR2_X1 U581 ( .A(KEYINPUT97), .B(KEYINPUT21), .Z(n472) );
  INV_X1 U582 ( .A(n469), .ZN(n607) );
  NAND2_X1 U583 ( .A1(G234), .A2(n607), .ZN(n470) );
  XNOR2_X1 U584 ( .A(n470), .B(KEYINPUT20), .ZN(n484) );
  NAND2_X1 U585 ( .A1(G221), .A2(n484), .ZN(n471) );
  XNOR2_X1 U586 ( .A(n472), .B(n471), .ZN(n647) );
  XNOR2_X1 U587 ( .A(KEYINPUT24), .B(KEYINPUT94), .ZN(n476) );
  XNOR2_X1 U588 ( .A(n476), .B(KEYINPUT95), .ZN(n477) );
  XOR2_X1 U589 ( .A(KEYINPUT8), .B(KEYINPUT66), .Z(n479) );
  NAND2_X1 U590 ( .A1(G234), .A2(n720), .ZN(n478) );
  XNOR2_X1 U591 ( .A(n479), .B(n478), .ZN(n510) );
  NAND2_X1 U592 ( .A1(n510), .A2(G221), .ZN(n480) );
  XNOR2_X1 U593 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U594 ( .A(KEYINPUT25), .B(KEYINPUT72), .Z(n486) );
  NAND2_X1 U595 ( .A1(G217), .A2(n484), .ZN(n485) );
  XNOR2_X1 U596 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U597 ( .A(n489), .B(KEYINPUT14), .ZN(n491) );
  NAND2_X1 U598 ( .A1(G952), .A2(n491), .ZN(n671) );
  NOR2_X1 U599 ( .A1(n671), .A2(G953), .ZN(n490) );
  XNOR2_X1 U600 ( .A(n490), .B(KEYINPUT91), .ZN(n566) );
  NAND2_X1 U601 ( .A1(n491), .A2(G902), .ZN(n492) );
  XNOR2_X1 U602 ( .A(KEYINPUT92), .B(n492), .ZN(n564) );
  NOR2_X1 U603 ( .A1(G900), .A2(n564), .ZN(n493) );
  NAND2_X1 U604 ( .A1(G953), .A2(n493), .ZN(n494) );
  NAND2_X1 U605 ( .A1(n566), .A2(n494), .ZN(n550) );
  NAND2_X1 U606 ( .A1(n495), .A2(n550), .ZN(n541) );
  XNOR2_X1 U607 ( .A(KEYINPUT13), .B(G475), .ZN(n504) );
  XOR2_X1 U608 ( .A(G122), .B(G104), .Z(n496) );
  XOR2_X1 U609 ( .A(KEYINPUT100), .B(KEYINPUT11), .Z(n498) );
  XNOR2_X1 U610 ( .A(n498), .B(n497), .ZN(n499) );
  NAND2_X1 U611 ( .A1(G214), .A2(n518), .ZN(n500) );
  XNOR2_X1 U612 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U613 ( .A(n503), .B(n502), .Z(n689) );
  XNOR2_X1 U614 ( .A(n549), .B(KEYINPUT101), .ZN(n556) );
  INV_X1 U615 ( .A(n505), .ZN(n509) );
  XNOR2_X1 U616 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U617 ( .A(n509), .B(n508), .ZN(n512) );
  NAND2_X1 U618 ( .A1(G217), .A2(n510), .ZN(n511) );
  XNOR2_X1 U619 ( .A(n512), .B(n511), .ZN(n514) );
  XNOR2_X1 U620 ( .A(n514), .B(n513), .ZN(n695) );
  XNOR2_X1 U621 ( .A(KEYINPUT104), .B(n515), .ZN(n557) );
  XNOR2_X1 U622 ( .A(n517), .B(n516), .ZN(n519) );
  XNOR2_X2 U623 ( .A(n524), .B(G472), .ZN(n644) );
  XNOR2_X1 U624 ( .A(n644), .B(KEYINPUT106), .ZN(n526) );
  INV_X1 U625 ( .A(KEYINPUT6), .ZN(n525) );
  XNOR2_X1 U626 ( .A(n526), .B(n525), .ZN(n588) );
  INV_X1 U627 ( .A(n588), .ZN(n577) );
  NAND2_X1 U628 ( .A1(G214), .A2(n527), .ZN(n655) );
  NAND2_X1 U629 ( .A1(n531), .A2(n655), .ZN(n528) );
  NOR2_X1 U630 ( .A1(n579), .A2(n528), .ZN(n529) );
  XNOR2_X1 U631 ( .A(n529), .B(KEYINPUT43), .ZN(n530) );
  NOR2_X1 U632 ( .A1(n642), .A2(n532), .ZN(n637) );
  NOR2_X1 U633 ( .A1(n647), .A2(n646), .ZN(n533) );
  XNOR2_X1 U634 ( .A(n533), .B(KEYINPUT65), .ZN(n641) );
  INV_X1 U635 ( .A(n641), .ZN(n535) );
  INV_X1 U636 ( .A(n534), .ZN(n594) );
  AND2_X1 U637 ( .A1(n535), .A2(n594), .ZN(n552) );
  NAND2_X1 U638 ( .A1(n536), .A2(n655), .ZN(n538) );
  XOR2_X1 U639 ( .A(KEYINPUT30), .B(KEYINPUT110), .Z(n537) );
  XNOR2_X1 U640 ( .A(n538), .B(n537), .ZN(n551) );
  NOR2_X1 U641 ( .A1(n549), .A2(n557), .ZN(n576) );
  INV_X1 U642 ( .A(n576), .ZN(n659) );
  XNOR2_X1 U643 ( .A(KEYINPUT112), .B(KEYINPUT41), .ZN(n539) );
  XNOR2_X1 U644 ( .A(n540), .B(n539), .ZN(n673) );
  XNOR2_X1 U645 ( .A(n542), .B(KEYINPUT28), .ZN(n544) );
  XOR2_X1 U646 ( .A(n594), .B(KEYINPUT111), .Z(n543) );
  NAND2_X1 U647 ( .A1(n544), .A2(n543), .ZN(n558) );
  NOR2_X1 U648 ( .A1(n673), .A2(n558), .ZN(n545) );
  XOR2_X1 U649 ( .A(KEYINPUT42), .B(n545), .Z(n732) );
  NAND2_X1 U650 ( .A1(n730), .A2(n732), .ZN(n547) );
  XNOR2_X1 U651 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n546) );
  XNOR2_X1 U652 ( .A(n547), .B(n355), .ZN(n548) );
  NAND2_X1 U653 ( .A1(n549), .A2(n557), .ZN(n572) );
  AND2_X1 U654 ( .A1(n551), .A2(n550), .ZN(n553) );
  AND2_X1 U655 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U656 ( .A1(n572), .A2(n555), .ZN(n628) );
  NAND2_X1 U657 ( .A1(n557), .A2(n556), .ZN(n635) );
  INV_X1 U658 ( .A(n635), .ZN(n562) );
  NOR2_X1 U659 ( .A1(n619), .A2(n562), .ZN(n662) );
  NAND2_X1 U660 ( .A1(n563), .A2(n562), .ZN(n639) );
  INV_X1 U661 ( .A(KEYINPUT44), .ZN(n584) );
  INV_X1 U662 ( .A(n564), .ZN(n565) );
  NOR2_X1 U663 ( .A1(G898), .A2(n720), .ZN(n704) );
  NAND2_X1 U664 ( .A1(n565), .A2(n704), .ZN(n567) );
  NAND2_X1 U665 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U666 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U667 ( .A(n572), .B(KEYINPUT76), .Z(n573) );
  XNOR2_X1 U668 ( .A(KEYINPUT83), .B(KEYINPUT35), .ZN(n574) );
  NAND2_X1 U669 ( .A1(n584), .A2(n725), .ZN(n586) );
  NOR2_X1 U670 ( .A1(n580), .A2(n351), .ZN(n578) );
  XNOR2_X1 U671 ( .A(n578), .B(KEYINPUT32), .ZN(n729) );
  AND2_X1 U672 ( .A1(n646), .A2(n581), .ZN(n582) );
  NAND2_X1 U673 ( .A1(n587), .A2(n582), .ZN(n583) );
  XNOR2_X1 U674 ( .A(n583), .B(KEYINPUT109), .ZN(n728) );
  NAND2_X1 U675 ( .A1(n584), .A2(KEYINPUT86), .ZN(n585) );
  NAND2_X1 U676 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U677 ( .A1(n646), .A2(n589), .ZN(n590) );
  XOR2_X1 U678 ( .A(KEYINPUT107), .B(n590), .Z(n726) );
  NOR2_X1 U679 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U680 ( .A1(n594), .A2(n593), .ZN(n623) );
  XNOR2_X1 U681 ( .A(KEYINPUT99), .B(KEYINPUT31), .ZN(n599) );
  NOR2_X1 U682 ( .A1(n644), .A2(n595), .ZN(n652) );
  NAND2_X1 U683 ( .A1(n652), .A2(n597), .ZN(n598) );
  XNOR2_X1 U684 ( .A(n599), .B(n598), .ZN(n634) );
  NAND2_X1 U685 ( .A1(n623), .A2(n634), .ZN(n601) );
  INV_X1 U686 ( .A(n662), .ZN(n600) );
  NAND2_X1 U687 ( .A1(n603), .A2(n602), .ZN(n605) );
  XNOR2_X2 U688 ( .A(n605), .B(n604), .ZN(n705) );
  INV_X1 U689 ( .A(KEYINPUT2), .ZN(n678) );
  NAND2_X1 U690 ( .A1(KEYINPUT2), .A2(n639), .ZN(n608) );
  INV_X1 U691 ( .A(KEYINPUT121), .ZN(n611) );
  XNOR2_X1 U692 ( .A(n612), .B(KEYINPUT62), .ZN(n614) );
  INV_X1 U693 ( .A(KEYINPUT114), .ZN(n616) );
  INV_X1 U694 ( .A(n619), .ZN(n632) );
  NOR2_X1 U695 ( .A1(n632), .A2(n623), .ZN(n620) );
  XOR2_X1 U696 ( .A(G104), .B(n620), .Z(G6) );
  XOR2_X1 U697 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n622) );
  XNOR2_X1 U698 ( .A(G107), .B(KEYINPUT116), .ZN(n621) );
  XNOR2_X1 U699 ( .A(n622), .B(n621), .ZN(n625) );
  NOR2_X1 U700 ( .A1(n635), .A2(n623), .ZN(n624) );
  XOR2_X1 U701 ( .A(n625), .B(n624), .Z(G9) );
  NOR2_X1 U702 ( .A1(n635), .A2(n629), .ZN(n627) );
  XNOR2_X1 U703 ( .A(G128), .B(KEYINPUT29), .ZN(n626) );
  XNOR2_X1 U704 ( .A(n627), .B(n626), .ZN(G30) );
  XOR2_X1 U705 ( .A(G143), .B(n628), .Z(G45) );
  NOR2_X1 U706 ( .A1(n632), .A2(n629), .ZN(n631) );
  XNOR2_X1 U707 ( .A(G146), .B(KEYINPUT117), .ZN(n630) );
  XNOR2_X1 U708 ( .A(n631), .B(n630), .ZN(G48) );
  NOR2_X1 U709 ( .A1(n632), .A2(n634), .ZN(n633) );
  XOR2_X1 U710 ( .A(G113), .B(n633), .Z(G15) );
  NOR2_X1 U711 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U712 ( .A(G116), .B(n636), .Z(G18) );
  XNOR2_X1 U713 ( .A(G125), .B(n637), .ZN(n638) );
  XNOR2_X1 U714 ( .A(n638), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U715 ( .A(G134), .B(n639), .ZN(G36) );
  XOR2_X1 U716 ( .A(G140), .B(n640), .Z(G42) );
  NAND2_X1 U717 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U718 ( .A(n643), .B(KEYINPUT50), .ZN(n645) );
  NAND2_X1 U719 ( .A1(n645), .A2(n644), .ZN(n650) );
  NAND2_X1 U720 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U721 ( .A(KEYINPUT49), .B(n648), .ZN(n649) );
  NOR2_X1 U722 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U723 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U724 ( .A(KEYINPUT51), .B(n653), .Z(n654) );
  NOR2_X1 U725 ( .A1(n673), .A2(n654), .ZN(n668) );
  NOR2_X1 U726 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U727 ( .A(n657), .B(KEYINPUT118), .ZN(n658) );
  NOR2_X1 U728 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U729 ( .A(KEYINPUT119), .B(n660), .Z(n665) );
  NOR2_X1 U730 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U731 ( .A(KEYINPUT120), .B(n663), .ZN(n664) );
  NOR2_X1 U732 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U733 ( .A1(n666), .A2(n672), .ZN(n667) );
  NOR2_X1 U734 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U735 ( .A(n669), .B(KEYINPUT52), .ZN(n670) );
  NOR2_X1 U736 ( .A1(n671), .A2(n670), .ZN(n675) );
  NOR2_X1 U737 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U738 ( .A1(n675), .A2(n674), .ZN(n683) );
  NAND2_X1 U739 ( .A1(n705), .A2(n678), .ZN(n676) );
  XOR2_X1 U740 ( .A(n676), .B(KEYINPUT79), .Z(n680) );
  NAND2_X1 U741 ( .A1(n716), .A2(n678), .ZN(n679) );
  NAND2_X1 U742 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U743 ( .A1(n698), .A2(G469), .ZN(n687) );
  XOR2_X1 U744 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n684) );
  NOR2_X1 U745 ( .A1(n702), .A2(n688), .ZN(G54) );
  NAND2_X1 U746 ( .A1(n359), .A2(G475), .ZN(n690) );
  NOR2_X2 U747 ( .A1(n692), .A2(n702), .ZN(n693) );
  XNOR2_X1 U748 ( .A(n693), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U749 ( .A1(n698), .A2(G478), .ZN(n694) );
  NOR2_X1 U750 ( .A1(n702), .A2(n696), .ZN(G63) );
  XOR2_X1 U751 ( .A(n697), .B(KEYINPUT123), .Z(n700) );
  NAND2_X1 U752 ( .A1(n698), .A2(G217), .ZN(n699) );
  XNOR2_X1 U753 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U754 ( .A1(n702), .A2(n701), .ZN(G66) );
  NOR2_X1 U755 ( .A1(n703), .A2(n704), .ZN(n712) );
  OR2_X1 U756 ( .A1(G953), .A2(n705), .ZN(n709) );
  NAND2_X1 U757 ( .A1(G953), .A2(G224), .ZN(n706) );
  XNOR2_X1 U758 ( .A(KEYINPUT61), .B(n706), .ZN(n707) );
  NAND2_X1 U759 ( .A1(n707), .A2(G898), .ZN(n708) );
  NAND2_X1 U760 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U761 ( .A(n710), .B(KEYINPUT124), .ZN(n711) );
  XNOR2_X1 U762 ( .A(n712), .B(n711), .ZN(G69) );
  XOR2_X1 U763 ( .A(n713), .B(KEYINPUT125), .Z(n714) );
  XNOR2_X1 U764 ( .A(n715), .B(n714), .ZN(n718) );
  XNOR2_X1 U765 ( .A(n718), .B(n716), .ZN(n717) );
  NAND2_X1 U766 ( .A1(n717), .A2(n720), .ZN(n723) );
  XNOR2_X1 U767 ( .A(n718), .B(G227), .ZN(n719) );
  NOR2_X1 U768 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U769 ( .A1(G900), .A2(n721), .ZN(n722) );
  NAND2_X1 U770 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U771 ( .A(KEYINPUT126), .B(n724), .Z(G72) );
  XOR2_X1 U772 ( .A(G122), .B(n725), .Z(G24) );
  XNOR2_X1 U773 ( .A(G101), .B(n726), .ZN(n727) );
  XNOR2_X1 U774 ( .A(n727), .B(KEYINPUT115), .ZN(G3) );
  XOR2_X1 U775 ( .A(G110), .B(n728), .Z(G12) );
  XOR2_X1 U776 ( .A(G119), .B(n729), .Z(G21) );
  XOR2_X1 U777 ( .A(n730), .B(G131), .Z(n731) );
  XNOR2_X1 U778 ( .A(KEYINPUT127), .B(n731), .ZN(G33) );
  XNOR2_X1 U779 ( .A(G137), .B(n732), .ZN(G39) );
endmodule

