//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 0 0 0 0 1 0 0 1 0 0 1 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 1 1 0 1 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1 1 1 0 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n842,
    new_n843, new_n844, new_n845, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(G8gat), .ZN(new_n203));
  INV_X1    g002(.A(G1gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT16), .ZN(new_n205));
  INV_X1    g004(.A(G22gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G15gat), .ZN(new_n207));
  INV_X1    g006(.A(G15gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G22gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT88), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n207), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n210), .B1(new_n207), .B2(new_n209), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n205), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n208), .A2(G22gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n206), .A2(G15gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT88), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n217), .A2(new_n204), .A3(new_n211), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n203), .B1(new_n214), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n211), .ZN(new_n220));
  AOI21_X1  g019(.A(KEYINPUT89), .B1(new_n220), .B2(new_n205), .ZN(new_n221));
  XOR2_X1   g020(.A(KEYINPUT90), .B(G8gat), .Z(new_n222));
  NAND2_X1  g021(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n220), .A2(KEYINPUT89), .A3(new_n205), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n219), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  AND2_X1   g026(.A1(KEYINPUT85), .A2(G29gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(KEYINPUT85), .A2(G29gat), .ZN(new_n229));
  OAI21_X1  g028(.A(G36gat), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT86), .ZN(new_n231));
  XNOR2_X1  g030(.A(KEYINPUT85), .B(G29gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT86), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n232), .A2(new_n233), .A3(G36gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT14), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n235), .B1(G29gat), .B2(G36gat), .ZN(new_n236));
  INV_X1    g035(.A(G29gat), .ZN(new_n237));
  INV_X1    g036(.A(G36gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n237), .A2(new_n238), .A3(KEYINPUT14), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n231), .A2(new_n234), .A3(new_n236), .A4(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT15), .ZN(new_n241));
  OR2_X1    g040(.A1(G43gat), .A2(G50gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(G43gat), .A2(G50gat), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT87), .B(G50gat), .ZN(new_n245));
  INV_X1    g044(.A(G43gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n244), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n240), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n239), .A2(new_n236), .ZN(new_n251));
  INV_X1    g050(.A(new_n229), .ZN(new_n252));
  NAND2_X1  g051(.A1(KEYINPUT85), .A2(G29gat), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n238), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n251), .B1(new_n254), .B2(new_n233), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n244), .B1(new_n255), .B2(new_n231), .ZN(new_n256));
  OAI21_X1  g055(.A(KEYINPUT17), .B1(new_n250), .B2(new_n256), .ZN(new_n257));
  AND2_X1   g056(.A1(new_n247), .A2(new_n248), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n231), .B(new_n255), .C1(new_n258), .C2(new_n244), .ZN(new_n259));
  INV_X1    g058(.A(new_n244), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n240), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT17), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n259), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n227), .A2(new_n257), .A3(new_n263), .ZN(new_n264));
  NOR3_X1   g063(.A1(new_n212), .A2(new_n213), .A3(G1gat), .ZN(new_n265));
  INV_X1    g064(.A(new_n205), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n266), .B1(new_n217), .B2(new_n211), .ZN(new_n267));
  OAI21_X1  g066(.A(G8gat), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n218), .B(new_n222), .C1(new_n267), .C2(KEYINPUT89), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n268), .B1(new_n269), .B2(new_n225), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT91), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n250), .A2(new_n256), .ZN(new_n272));
  AND3_X1   g071(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n271), .B1(new_n270), .B2(new_n272), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n202), .B(new_n264), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT18), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(KEYINPUT92), .A3(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT93), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n278), .B1(new_n270), .B2(new_n272), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n259), .A2(new_n261), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n227), .A2(KEYINPUT93), .A3(new_n280), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n279), .B(new_n281), .C1(new_n273), .C2(new_n274), .ZN(new_n282));
  XOR2_X1   g081(.A(new_n202), .B(KEYINPUT13), .Z(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(KEYINPUT91), .B1(new_n227), .B2(new_n280), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n276), .A2(KEYINPUT92), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n287), .A2(new_n202), .A3(new_n264), .A4(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n277), .A2(new_n284), .A3(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G113gat), .B(G141gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G169gat), .B(G197gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n295), .B(KEYINPUT12), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n290), .A2(new_n297), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n277), .A2(new_n284), .A3(new_n289), .A4(new_n296), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT5), .ZN(new_n302));
  XNOR2_X1  g101(.A(G113gat), .B(G120gat), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT1), .B1(new_n303), .B2(KEYINPUT67), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n304), .B1(KEYINPUT67), .B2(new_n303), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT68), .ZN(new_n306));
  XNOR2_X1  g105(.A(G127gat), .B(G134gat), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  AND3_X1   g107(.A1(new_n305), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n306), .B1(new_n305), .B2(new_n308), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n308), .A2(KEYINPUT69), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT1), .ZN(new_n313));
  INV_X1    g112(.A(new_n303), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT69), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n307), .A2(new_n315), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n312), .A2(new_n313), .A3(new_n314), .A4(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT77), .B(KEYINPUT2), .ZN(new_n318));
  INV_X1    g117(.A(G141gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n319), .A2(G148gat), .ZN(new_n320));
  INV_X1    g119(.A(G148gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n321), .A2(G141gat), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n318), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G155gat), .A2(G162gat), .ZN(new_n324));
  INV_X1    g123(.A(G155gat), .ZN(new_n325));
  INV_X1    g124(.A(G162gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n323), .A2(new_n324), .A3(new_n327), .ZN(new_n328));
  XOR2_X1   g127(.A(KEYINPUT78), .B(G141gat), .Z(new_n329));
  AOI21_X1  g128(.A(new_n320), .B1(new_n329), .B2(G148gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n327), .A2(KEYINPUT2), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n331), .B1(G155gat), .B2(G162gat), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n317), .B(new_n328), .C1(new_n330), .C2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT79), .B1(new_n311), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n305), .A2(new_n308), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT68), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n305), .A2(new_n306), .A3(new_n308), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n333), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT79), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n317), .B1(new_n309), .B2(new_n310), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n328), .B1(new_n330), .B2(new_n332), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n334), .A2(new_n341), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(G225gat), .A2(G233gat), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n302), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT3), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n343), .B(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n347), .B1(new_n350), .B2(new_n342), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n338), .A2(new_n339), .A3(KEYINPUT4), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n334), .A2(new_n341), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n351), .B(new_n352), .C1(new_n353), .C2(KEYINPUT4), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n348), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(KEYINPUT4), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT4), .B1(new_n338), .B2(new_n339), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n356), .A2(new_n302), .A3(new_n351), .A4(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(G1gat), .B(G29gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(KEYINPUT0), .ZN(new_n362));
  XNOR2_X1  g161(.A(G57gat), .B(G85gat), .ZN(new_n363));
  XOR2_X1   g162(.A(new_n362), .B(new_n363), .Z(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n360), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n355), .A2(new_n364), .A3(new_n359), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT80), .B(KEYINPUT6), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT27), .ZN(new_n370));
  INV_X1    g169(.A(G183gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(KEYINPUT66), .B(G183gat), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n372), .B1(new_n373), .B2(new_n370), .ZN(new_n374));
  INV_X1    g173(.A(G190gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT28), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(KEYINPUT27), .B(G183gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n379), .A2(KEYINPUT28), .A3(new_n375), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(G169gat), .ZN(new_n382));
  INV_X1    g181(.A(G176gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OR2_X1    g183(.A1(new_n384), .A2(KEYINPUT26), .ZN(new_n385));
  NOR2_X1   g184(.A1(G169gat), .A2(G176gat), .ZN(new_n386));
  OR2_X1    g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI22_X1  g186(.A1(new_n386), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n381), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(G226gat), .ZN(new_n390));
  INV_X1    g189(.A(G233gat), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n384), .B1(KEYINPUT23), .B2(new_n386), .ZN(new_n394));
  OR2_X1    g193(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n395));
  NAND2_X1  g194(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n395), .B(new_n396), .C1(G169gat), .C2(G176gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n371), .A2(new_n375), .ZN(new_n399));
  OAI21_X1  g198(.A(KEYINPUT24), .B1(new_n371), .B2(new_n375), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT24), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n401), .A2(G183gat), .A3(G190gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n398), .A2(KEYINPUT65), .B1(new_n399), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT65), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n394), .A2(new_n405), .A3(new_n397), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT25), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  AOI22_X1  g206(.A1(new_n373), .A2(new_n375), .B1(new_n400), .B2(new_n402), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT25), .ZN(new_n409));
  NOR3_X1   g208(.A1(new_n398), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n389), .B(new_n393), .C1(new_n407), .C2(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n392), .A2(KEYINPUT29), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT65), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n403), .A2(new_n399), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(new_n406), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n410), .B1(new_n416), .B2(new_n409), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n387), .A2(new_n388), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n418), .B1(new_n378), .B2(new_n380), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n413), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n411), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT22), .ZN(new_n422));
  AOI22_X1  g221(.A1(new_n422), .A2(KEYINPUT73), .B1(G211gat), .B2(G218gat), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT73), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT22), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G197gat), .B(G204gat), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT74), .ZN(new_n428));
  XNOR2_X1  g227(.A(G211gat), .B(G218gat), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n426), .B(new_n427), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n428), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  OR2_X1    g232(.A1(new_n429), .A2(new_n428), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n434), .A2(new_n431), .A3(new_n426), .A4(new_n427), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT75), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n433), .A2(new_n435), .A3(KEYINPUT75), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(KEYINPUT76), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT76), .ZN(new_n440));
  INV_X1    g239(.A(new_n438), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n440), .B1(new_n441), .B2(new_n436), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n421), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n441), .A2(new_n436), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n411), .A2(new_n420), .A3(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n444), .A2(KEYINPUT37), .A3(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(G8gat), .B(G36gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(G64gat), .B(G92gat), .ZN(new_n449));
  XOR2_X1   g248(.A(new_n448), .B(new_n449), .Z(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n447), .A2(KEYINPUT82), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n444), .A2(new_n446), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT37), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT82), .B1(new_n447), .B2(new_n451), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT38), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AOI211_X1 g257(.A(KEYINPUT38), .B(new_n450), .C1(new_n453), .C2(new_n454), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n421), .B1(new_n441), .B2(new_n436), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n460), .B(KEYINPUT37), .C1(new_n421), .C2(new_n443), .ZN(new_n461));
  AOI22_X1  g260(.A1(new_n459), .A2(new_n461), .B1(new_n450), .B2(new_n453), .ZN(new_n462));
  INV_X1    g261(.A(new_n368), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n360), .A2(new_n365), .A3(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n369), .A2(new_n458), .A3(new_n462), .A4(new_n464), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n411), .A2(new_n420), .A3(new_n445), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n411), .A2(new_n420), .B1(new_n442), .B2(new_n439), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n450), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n444), .A2(new_n451), .A3(new_n446), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n468), .A2(new_n469), .A3(KEYINPUT30), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT30), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n453), .A2(new_n471), .A3(new_n450), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n364), .B1(new_n355), .B2(new_n359), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n350), .A2(new_n342), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n356), .A2(new_n476), .A3(new_n358), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT39), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(new_n478), .A3(new_n347), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n364), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT39), .B1(new_n345), .B2(new_n347), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n481), .B1(new_n477), .B2(new_n347), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n480), .A2(KEYINPUT40), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT40), .ZN(new_n484));
  INV_X1    g283(.A(new_n482), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n357), .B1(new_n353), .B2(KEYINPUT4), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n346), .B1(new_n486), .B2(new_n476), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n365), .B1(new_n487), .B2(new_n478), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n484), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n475), .B1(new_n483), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT29), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n491), .B1(new_n343), .B2(KEYINPUT3), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n439), .A2(new_n442), .A3(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(G228gat), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n433), .A2(new_n435), .A3(new_n491), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n349), .ZN(new_n496));
  AOI211_X1 g295(.A(new_n494), .B(new_n391), .C1(new_n496), .C2(new_n343), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n437), .A2(new_n438), .A3(new_n492), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n496), .A2(new_n343), .ZN(new_n500));
  OAI22_X1  g299(.A1(new_n499), .A2(new_n500), .B1(new_n494), .B2(new_n391), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n206), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n498), .A2(new_n501), .A3(new_n206), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(G78gat), .B(G106gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(KEYINPUT31), .B(G50gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n508), .B1(new_n502), .B2(KEYINPUT81), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n503), .A2(KEYINPUT81), .A3(new_n504), .A4(new_n508), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n465), .A2(new_n490), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n367), .A2(new_n368), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n464), .B1(new_n514), .B2(new_n474), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n473), .ZN(new_n516));
  INV_X1    g315(.A(new_n512), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT36), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n342), .B(new_n389), .C1(new_n407), .C2(new_n410), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n338), .B(new_n317), .C1(new_n417), .C2(new_n419), .ZN(new_n521));
  INV_X1    g320(.A(G227gat), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n522), .A2(new_n391), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n520), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT33), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT70), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT70), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n524), .A2(new_n528), .A3(new_n525), .ZN(new_n529));
  XNOR2_X1  g328(.A(G15gat), .B(G43gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(G71gat), .B(G99gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n532), .B1(new_n524), .B2(KEYINPUT32), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n527), .A2(new_n529), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n523), .B1(new_n520), .B2(new_n521), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT34), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI211_X1 g336(.A(KEYINPUT34), .B(new_n523), .C1(new_n520), .C2(new_n521), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT71), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n525), .B1(new_n532), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n541), .B1(new_n540), .B2(new_n532), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n524), .A2(KEYINPUT32), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n534), .A2(new_n539), .A3(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n539), .B1(new_n534), .B2(new_n543), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n519), .B1(new_n547), .B2(KEYINPUT72), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n534), .A2(new_n543), .ZN(new_n549));
  INV_X1    g348(.A(new_n539), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(new_n544), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT72), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n552), .A2(new_n553), .A3(KEYINPUT36), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n513), .A2(new_n518), .A3(new_n548), .A4(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n512), .A2(new_n551), .A3(new_n544), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT35), .B1(new_n516), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT83), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT35), .B1(new_n470), .B2(new_n472), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n515), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n558), .B1(new_n560), .B2(new_n556), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT35), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n473), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n563), .B1(new_n369), .B2(new_n464), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n564), .A2(KEYINPUT83), .A3(new_n512), .A4(new_n547), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n557), .A2(new_n561), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n301), .B1(new_n555), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(G71gat), .A2(G78gat), .ZN(new_n568));
  OR2_X1    g367(.A1(G71gat), .A2(G78gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(G57gat), .B(G64gat), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT9), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n568), .B(new_n569), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(G64gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(G57gat), .ZN(new_n574));
  INV_X1    g373(.A(G57gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(G64gat), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT94), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n575), .A2(G64gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT94), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n569), .A2(new_n568), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n578), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT95), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n572), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT21), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G231gat), .A2(G233gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(G127gat), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n227), .B1(new_n586), .B2(new_n585), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n591), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(new_n325), .ZN(new_n596));
  XNOR2_X1  g395(.A(G183gat), .B(G211gat), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n596), .B(new_n597), .Z(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n592), .A2(new_n593), .A3(new_n598), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G190gat), .B(G218gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(KEYINPUT97), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT41), .ZN(new_n605));
  INV_X1    g404(.A(G232gat), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n605), .B1(new_n606), .B2(new_n391), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n604), .B(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT96), .ZN(new_n610));
  NAND2_X1  g409(.A1(G85gat), .A2(G92gat), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT7), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT7), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n613), .A2(G85gat), .A3(G92gat), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(G99gat), .A2(G106gat), .ZN(new_n616));
  INV_X1    g415(.A(G85gat), .ZN(new_n617));
  INV_X1    g416(.A(G92gat), .ZN(new_n618));
  AOI22_X1  g417(.A1(KEYINPUT8), .A2(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G99gat), .B(G106gat), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n615), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n620), .B1(new_n615), .B2(new_n619), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n610), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n615), .A2(new_n619), .ZN(new_n625));
  INV_X1    g424(.A(new_n620), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n627), .A2(KEYINPUT96), .A3(new_n621), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n257), .A2(new_n263), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n630), .B(new_n631), .C1(new_n280), .C2(new_n629), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n603), .A2(KEYINPUT97), .ZN(new_n633));
  XNOR2_X1  g432(.A(G134gat), .B(G162gat), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n632), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n635), .B1(new_n632), .B2(new_n633), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n609), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n638), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n640), .A2(new_n608), .A3(new_n636), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n602), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n621), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n585), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT95), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n583), .B(new_n646), .ZN(new_n647));
  AOI22_X1  g446(.A1(KEYINPUT94), .A2(new_n579), .B1(new_n569), .B2(new_n568), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n647), .A2(new_n578), .A3(new_n648), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n649), .A2(new_n572), .A3(new_n621), .A4(new_n627), .ZN(new_n650));
  XOR2_X1   g449(.A(KEYINPUT98), .B(KEYINPUT10), .Z(new_n651));
  NAND3_X1  g450(.A1(new_n645), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n585), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n653), .A2(new_n624), .A3(new_n628), .A4(KEYINPUT10), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(G230gat), .A2(G233gat), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n645), .A2(new_n650), .ZN(new_n658));
  INV_X1    g457(.A(new_n656), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(G120gat), .B(G148gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT99), .ZN(new_n663));
  XNOR2_X1  g462(.A(G176gat), .B(G204gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n661), .A2(new_n665), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n643), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(KEYINPUT100), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT100), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n672), .B1(new_n643), .B2(new_n669), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n567), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n675), .A2(new_n515), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(new_n204), .ZN(G1324gat));
  NOR2_X1   g476(.A1(new_n675), .A2(new_n473), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT16), .B(G8gat), .Z(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT101), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n681), .A2(new_n682), .A3(KEYINPUT42), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT42), .B1(new_n678), .B2(new_n203), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n680), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n682), .B1(new_n681), .B2(KEYINPUT42), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n683), .B1(new_n685), .B2(new_n686), .ZN(G1325gat));
  INV_X1    g486(.A(new_n675), .ZN(new_n688));
  AOI21_X1  g487(.A(G15gat), .B1(new_n688), .B2(new_n547), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n548), .A2(new_n554), .ZN(new_n690));
  OR2_X1    g489(.A1(new_n690), .A2(KEYINPUT102), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(KEYINPUT102), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n693), .A2(new_n208), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT103), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n689), .B1(new_n695), .B2(new_n688), .ZN(G1326gat));
  OR3_X1    g495(.A1(new_n675), .A2(KEYINPUT104), .A3(new_n512), .ZN(new_n697));
  OAI21_X1  g496(.A(KEYINPUT104), .B1(new_n675), .B2(new_n512), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT43), .B(G22gat), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1327gat));
  INV_X1    g500(.A(new_n602), .ZN(new_n702));
  INV_X1    g501(.A(new_n669), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n704), .A2(new_n642), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n567), .A2(new_n705), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n706), .A2(new_n515), .A3(new_n232), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT45), .Z(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n555), .A2(new_n566), .ZN(new_n710));
  INV_X1    g509(.A(new_n642), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n713), .A2(KEYINPUT106), .ZN(new_n714));
  AOI211_X1 g513(.A(new_n642), .B(new_n714), .C1(new_n555), .C2(new_n566), .ZN(new_n715));
  OR2_X1    g514(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n298), .A2(KEYINPUT105), .A3(new_n299), .ZN(new_n717));
  AOI21_X1  g516(.A(KEYINPUT105), .B1(new_n298), .B2(new_n299), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n704), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n232), .B1(new_n721), .B2(new_n515), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n708), .A2(new_n722), .ZN(G1328gat));
  OAI21_X1  g522(.A(G36gat), .B1(new_n721), .B2(new_n473), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n706), .A2(G36gat), .A3(new_n473), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT46), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(G1329gat));
  NAND4_X1  g526(.A1(new_n567), .A2(new_n246), .A3(new_n547), .A4(new_n705), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n728), .A2(KEYINPUT108), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(KEYINPUT108), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n690), .B(new_n720), .C1(new_n712), .C2(new_n715), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(G43gat), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n731), .A2(new_n733), .A3(KEYINPUT47), .ZN(new_n734));
  INV_X1    g533(.A(new_n693), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n735), .B(new_n720), .C1(new_n712), .C2(new_n715), .ZN(new_n736));
  AOI22_X1  g535(.A1(new_n729), .A2(new_n730), .B1(new_n736), .B2(G43gat), .ZN(new_n737));
  XOR2_X1   g536(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n738));
  OAI21_X1  g537(.A(new_n734), .B1(new_n737), .B2(new_n738), .ZN(G1330gat));
  NOR2_X1   g538(.A1(new_n512), .A2(new_n245), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n720), .B(new_n740), .C1(new_n712), .C2(new_n715), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n245), .B1(new_n706), .B2(new_n512), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g543(.A(new_n719), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n745), .A2(new_n643), .A3(new_n703), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n710), .A2(new_n746), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n515), .B(KEYINPUT109), .Z(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g549(.A(new_n473), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT110), .ZN(new_n753));
  NOR2_X1   g552(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1333gat));
  NAND2_X1  g554(.A1(new_n747), .A2(new_n735), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n552), .A2(G71gat), .ZN(new_n757));
  AOI22_X1  g556(.A1(new_n756), .A2(G71gat), .B1(new_n747), .B2(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g558(.A1(new_n747), .A2(new_n517), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g560(.A1(new_n745), .A2(new_n602), .A3(new_n703), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n716), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(G85gat), .B1(new_n763), .B2(new_n515), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n642), .B1(new_n555), .B2(new_n566), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n745), .A2(new_n602), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n765), .A2(KEYINPUT51), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT51), .B1(new_n765), .B2(new_n766), .ZN(new_n768));
  OR2_X1    g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n515), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n769), .A2(new_n617), .A3(new_n770), .A4(new_n669), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n764), .A2(new_n771), .ZN(G1336gat));
  INV_X1    g571(.A(new_n473), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n773), .B(new_n762), .C1(new_n712), .C2(new_n715), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(G92gat), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n473), .A2(G92gat), .A3(new_n703), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(new_n767), .B2(new_n768), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g578(.A(G99gat), .B1(new_n763), .B2(new_n693), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n552), .A2(G99gat), .A3(new_n703), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n769), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(G1338gat));
  NOR3_X1   g582(.A1(new_n512), .A2(G106gat), .A3(new_n703), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(new_n767), .B2(new_n768), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT112), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n517), .B(new_n762), .C1(new_n712), .C2(new_n715), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n787), .A2(KEYINPUT111), .A3(G106gat), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT112), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n789), .B(new_n784), .C1(new_n767), .C2(new_n768), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n786), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT53), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n787), .A2(G106gat), .ZN(new_n793));
  NAND2_X1  g592(.A1(KEYINPUT111), .A2(KEYINPUT53), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n793), .B(new_n794), .C1(KEYINPUT53), .C2(new_n785), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n792), .A2(new_n795), .ZN(G1339gat));
  NAND3_X1  g595(.A1(new_n652), .A2(new_n654), .A3(new_n659), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(KEYINPUT113), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT113), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n652), .A2(new_n654), .A3(new_n799), .A4(new_n659), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n659), .B1(new_n652), .B2(new_n654), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(new_n665), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n806), .B1(new_n802), .B2(new_n803), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n805), .A2(KEYINPUT55), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n667), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n665), .B1(new_n657), .B2(KEYINPUT54), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n810), .B1(new_n801), .B2(new_n804), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n811), .A2(KEYINPUT55), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n813), .B1(new_n717), .B2(new_n718), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n282), .A2(new_n283), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n202), .B1(new_n287), .B2(new_n264), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n295), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n299), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n669), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n711), .B1(new_n814), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n666), .B1(new_n811), .B2(KEYINPUT55), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n807), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n299), .A2(new_n817), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n825), .A2(new_n642), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n702), .B1(new_n820), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n670), .A2(new_n719), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n556), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n748), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n831), .A2(new_n773), .ZN(new_n832));
  AOI21_X1  g631(.A(G113gat), .B1(new_n832), .B2(new_n745), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n770), .A2(new_n473), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n830), .A2(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n300), .A2(G113gat), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n833), .B1(new_n836), .B2(new_n837), .ZN(G1340gat));
  AOI21_X1  g637(.A(G120gat), .B1(new_n832), .B2(new_n669), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n669), .A2(G120gat), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n839), .B1(new_n836), .B2(new_n840), .ZN(G1341gat));
  INV_X1    g640(.A(new_n836), .ZN(new_n842));
  OAI21_X1  g641(.A(G127gat), .B1(new_n842), .B2(new_n702), .ZN(new_n843));
  INV_X1    g642(.A(G127gat), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n832), .A2(new_n844), .A3(new_n602), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(G1342gat));
  OAI21_X1  g645(.A(G134gat), .B1(new_n842), .B2(new_n642), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n773), .A2(new_n642), .ZN(new_n848));
  INV_X1    g647(.A(G134gat), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(KEYINPUT56), .B1(new_n831), .B2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT115), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n851), .A2(new_n852), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n831), .A2(KEYINPUT56), .A3(new_n850), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(KEYINPUT114), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n855), .A2(KEYINPUT114), .ZN(new_n857));
  OAI221_X1 g656(.A(new_n847), .B1(new_n853), .B2(new_n854), .C1(new_n856), .C2(new_n857), .ZN(G1343gat));
  NAND2_X1  g657(.A1(new_n828), .A2(new_n829), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n693), .A2(new_n517), .A3(new_n748), .A4(new_n859), .ZN(new_n860));
  NOR4_X1   g659(.A1(new_n860), .A2(G141gat), .A3(new_n301), .A4(new_n773), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(KEYINPUT58), .ZN(new_n862));
  INV_X1    g661(.A(new_n329), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n690), .A2(new_n834), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT57), .B1(new_n859), .B2(new_n517), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT57), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n512), .A2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n711), .A2(new_n813), .A3(new_n818), .ZN(new_n869));
  AOI22_X1  g668(.A1(new_n300), .A2(new_n813), .B1(new_n818), .B2(new_n669), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n869), .B1(new_n870), .B2(new_n711), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(KEYINPUT116), .A3(new_n702), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n872), .A2(new_n829), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT116), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n300), .A2(new_n813), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n819), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n827), .B1(new_n876), .B2(new_n642), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n874), .B1(new_n877), .B2(new_n602), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n868), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n864), .B1(new_n865), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n863), .B1(new_n880), .B2(new_n301), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n862), .A2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT105), .ZN(new_n883));
  INV_X1    g682(.A(new_n275), .ZN(new_n884));
  AOI22_X1  g683(.A1(new_n884), .A2(new_n288), .B1(new_n283), .B2(new_n282), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n296), .B1(new_n885), .B2(new_n277), .ZN(new_n886));
  INV_X1    g685(.A(new_n299), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n883), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n298), .A2(KEYINPUT105), .A3(new_n299), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n825), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n819), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n642), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n602), .B1(new_n892), .B2(new_n869), .ZN(new_n893));
  INV_X1    g692(.A(new_n829), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n517), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n878), .A2(new_n829), .A3(new_n872), .ZN(new_n896));
  AOI22_X1  g695(.A1(new_n895), .A2(new_n866), .B1(new_n867), .B2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n864), .ZN(new_n898));
  OAI21_X1  g697(.A(KEYINPUT117), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT117), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n900), .B(new_n864), .C1(new_n865), .C2(new_n879), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n899), .A2(new_n745), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n861), .B1(new_n902), .B2(new_n863), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT58), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n882), .B1(new_n903), .B2(new_n904), .ZN(G1344gat));
  NAND2_X1  g704(.A1(new_n859), .A2(new_n867), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT118), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n871), .A2(new_n907), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n869), .B(KEYINPUT118), .C1(new_n870), .C2(new_n711), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n909), .A3(new_n702), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n671), .A2(new_n301), .A3(new_n673), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n512), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n906), .B1(new_n912), .B2(KEYINPUT57), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n913), .A2(new_n669), .A3(new_n864), .ZN(new_n914));
  OAI21_X1  g713(.A(KEYINPUT59), .B1(new_n914), .B2(new_n321), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n899), .A2(new_n669), .A3(new_n901), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n321), .A2(KEYINPUT59), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n860), .A2(new_n773), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n321), .A3(new_n669), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1345gat));
  NAND3_X1  g720(.A1(new_n919), .A2(new_n325), .A3(new_n602), .ZN(new_n922));
  AND3_X1   g721(.A1(new_n899), .A2(new_n602), .A3(new_n901), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n923), .B2(new_n325), .ZN(G1346gat));
  NAND3_X1  g723(.A1(new_n899), .A2(new_n711), .A3(new_n901), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT119), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT119), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n899), .A2(new_n901), .A3(new_n927), .A4(new_n711), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n926), .A2(G162gat), .A3(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(new_n860), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n930), .A2(new_n326), .A3(new_n848), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(G1347gat));
  NOR2_X1   g731(.A1(new_n748), .A2(new_n473), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n830), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(G169gat), .B1(new_n934), .B2(new_n301), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT120), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n935), .A2(new_n936), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n770), .B1(new_n828), .B2(new_n829), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n939), .A2(new_n512), .A3(new_n773), .A4(new_n547), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n745), .A2(new_n382), .ZN(new_n941));
  OAI22_X1  g740(.A1(new_n937), .A2(new_n938), .B1(new_n940), .B2(new_n941), .ZN(G1348gat));
  OAI21_X1  g741(.A(G176gat), .B1(new_n934), .B2(new_n703), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n669), .A2(new_n383), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n940), .B2(new_n944), .ZN(G1349gat));
  NOR2_X1   g744(.A1(new_n934), .A2(new_n702), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n946), .A2(new_n373), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n602), .A2(new_n379), .ZN(new_n948));
  OR2_X1    g747(.A1(new_n940), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n947), .A2(KEYINPUT121), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(KEYINPUT60), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT60), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n947), .A2(KEYINPUT121), .A3(new_n952), .A4(new_n949), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n953), .ZN(G1350gat));
  NOR3_X1   g753(.A1(new_n940), .A2(G190gat), .A3(new_n642), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT122), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n375), .B1(KEYINPUT123), .B2(KEYINPUT61), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n957), .B1(new_n934), .B2(new_n642), .ZN(new_n958));
  NOR2_X1   g757(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n959));
  OR2_X1    g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n959), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n956), .A2(new_n960), .A3(new_n961), .ZN(G1351gat));
  AOI211_X1 g761(.A(new_n473), .B(new_n748), .C1(new_n691), .C2(new_n692), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n913), .A2(G197gat), .A3(new_n300), .A4(new_n963), .ZN(new_n964));
  INV_X1    g763(.A(G197gat), .ZN(new_n965));
  NAND4_X1  g764(.A1(new_n693), .A2(new_n939), .A3(new_n517), .A4(new_n773), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n965), .B1(new_n966), .B2(new_n719), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n964), .A2(new_n967), .ZN(G1352gat));
  NAND3_X1  g767(.A1(new_n913), .A2(new_n669), .A3(new_n963), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(G204gat), .ZN(new_n970));
  OR2_X1    g769(.A1(new_n703), .A2(G204gat), .ZN(new_n971));
  OR3_X1    g770(.A1(new_n966), .A2(KEYINPUT62), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g771(.A(KEYINPUT62), .B1(new_n966), .B2(new_n971), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n970), .A2(new_n972), .A3(new_n973), .ZN(G1353gat));
  NOR3_X1   g773(.A1(new_n966), .A2(G211gat), .A3(new_n702), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n913), .A2(new_n602), .A3(new_n963), .ZN(new_n976));
  AOI21_X1  g775(.A(KEYINPUT63), .B1(new_n976), .B2(G211gat), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT124), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n975), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n976), .A2(G211gat), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT63), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(KEYINPUT124), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n980), .A2(new_n981), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n979), .B1(new_n983), .B2(new_n984), .ZN(G1354gat));
  INV_X1    g784(.A(G218gat), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n986), .B1(new_n966), .B2(new_n642), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT125), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n913), .A2(new_n988), .A3(new_n963), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n711), .A2(G218gat), .ZN(new_n990));
  XNOR2_X1  g789(.A(new_n990), .B(KEYINPUT126), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n988), .B1(new_n913), .B2(new_n963), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n987), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT127), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI211_X1 g795(.A(KEYINPUT127), .B(new_n987), .C1(new_n992), .C2(new_n993), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n996), .A2(new_n997), .ZN(G1355gat));
endmodule


