//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 1 0 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n494, new_n495, new_n496, new_n497, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n583, new_n584, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n593, new_n594, new_n595, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n627, new_n630, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT66), .Z(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(new_n453), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(KEYINPUT3), .A3(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT69), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n465), .A2(KEYINPUT69), .A3(KEYINPUT3), .A4(new_n466), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(KEYINPUT70), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT70), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n476), .A2(new_n473), .A3(G2104), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n471), .A2(new_n472), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G137), .ZN(new_n481));
  AND2_X1   g056(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n482));
  NOR2_X1   g057(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G101), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT71), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n481), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(G113), .A2(G2104), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n474), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G125), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n495));
  XNOR2_X1  g070(.A(new_n494), .B(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n488), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G160));
  INV_X1    g073(.A(G136), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n472), .A2(G112), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n501));
  OAI22_X1  g076(.A1(new_n479), .A2(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n475), .A2(new_n477), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n503), .B1(new_n469), .B2(new_n470), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G2105), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT72), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n504), .A2(KEYINPUT72), .A3(G2105), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n502), .B1(new_n509), .B2(G124), .ZN(G162));
  NAND3_X1  g085(.A1(new_n504), .A2(G138), .A3(new_n472), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT4), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT3), .B(G2104), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT4), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n513), .A2(new_n514), .A3(G138), .A4(new_n472), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT75), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n515), .B(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  AND2_X1   g094(.A1(G126), .A2(G2105), .ZN(new_n520));
  AOI21_X1  g095(.A(KEYINPUT69), .B1(new_n484), .B2(KEYINPUT3), .ZN(new_n521));
  NOR4_X1   g096(.A1(new_n482), .A2(new_n483), .A3(new_n468), .A4(new_n473), .ZN(new_n522));
  OAI211_X1 g097(.A(new_n478), .B(new_n520), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT73), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n504), .A2(new_n525), .A3(new_n520), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g102(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n528));
  INV_X1    g103(.A(G114), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n528), .B1(new_n529), .B2(G2105), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g106(.A(KEYINPUT74), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT74), .ZN(new_n533));
  AOI211_X1 g108(.A(new_n533), .B(new_n530), .C1(new_n524), .C2(new_n526), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n519), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(G164));
  AND2_X1   g111(.A1(KEYINPUT6), .A2(G651), .ZN(new_n537));
  NOR2_X1   g112(.A1(KEYINPUT6), .A2(G651), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G50), .ZN(new_n542));
  AND2_X1   g117(.A1(KEYINPUT5), .A2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(KEYINPUT5), .A2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n539), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(G88), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n542), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n545), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n550), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G651), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n549), .A2(new_n553), .ZN(G166));
  NAND3_X1  g129(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT7), .ZN(new_n556));
  INV_X1    g131(.A(new_n539), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G51), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n556), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(G89), .ZN(new_n561));
  NAND2_X1  g136(.A1(G63), .A2(G651), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n545), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n560), .A2(new_n563), .ZN(G168));
  NAND2_X1  g139(.A1(G77), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G64), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n545), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT76), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n552), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n569), .B1(new_n568), .B2(new_n567), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n546), .A2(G90), .B1(new_n541), .B2(G52), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(G301));
  INV_X1    g147(.A(G301), .ZN(G171));
  NAND2_X1  g148(.A1(new_n546), .A2(G81), .ZN(new_n574));
  INV_X1    g149(.A(G43), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n575), .B2(new_n558), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n550), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n577), .A2(new_n552), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G860), .ZN(G153));
  NAND4_X1  g155(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n581));
  XOR2_X1   g156(.A(new_n581), .B(KEYINPUT77), .Z(G176));
  NAND2_X1  g157(.A1(G1), .A2(G3), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT8), .ZN(new_n584));
  NAND4_X1  g159(.A1(G319), .A2(G483), .A3(G661), .A4(new_n584), .ZN(G188));
  NAND2_X1  g160(.A1(new_n541), .A2(G53), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT9), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n550), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n588), .A2(new_n552), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n546), .A2(G91), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n587), .A2(new_n589), .A3(new_n590), .ZN(G299));
  INV_X1    g166(.A(G168), .ZN(G286));
  NAND2_X1  g167(.A1(G166), .A2(KEYINPUT78), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT78), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(new_n549), .B2(new_n553), .ZN(new_n595));
  AND2_X1   g170(.A1(new_n593), .A2(new_n595), .ZN(G303));
  NAND2_X1  g171(.A1(new_n546), .A2(G87), .ZN(new_n597));
  OAI21_X1  g172(.A(G651), .B1(new_n550), .B2(G74), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n541), .A2(G49), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(G288));
  INV_X1    g175(.A(G86), .ZN(new_n601));
  OAI21_X1  g176(.A(KEYINPUT79), .B1(new_n547), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(G73), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G61), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n545), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n605), .A2(G651), .B1(new_n541), .B2(G48), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT79), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n546), .A2(new_n607), .A3(G86), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n602), .A2(new_n606), .A3(new_n608), .ZN(G305));
  AOI22_X1  g184(.A1(new_n546), .A2(G85), .B1(new_n541), .B2(G47), .ZN(new_n610));
  AND2_X1   g185(.A1(new_n610), .A2(KEYINPUT80), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n610), .A2(KEYINPUT80), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n550), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n613));
  OAI22_X1  g188(.A1(new_n611), .A2(new_n612), .B1(new_n552), .B2(new_n613), .ZN(G290));
  NAND2_X1  g189(.A1(G301), .A2(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n546), .A2(G92), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT10), .Z(new_n617));
  NAND2_X1  g192(.A1(G79), .A2(G543), .ZN(new_n618));
  XOR2_X1   g193(.A(KEYINPUT81), .B(G66), .Z(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n545), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n620), .A2(G651), .B1(new_n541), .B2(G54), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n615), .B1(new_n623), .B2(G868), .ZN(G321));
  XOR2_X1   g199(.A(G321), .B(KEYINPUT82), .Z(G284));
  NAND2_X1  g200(.A1(G286), .A2(G868), .ZN(new_n626));
  AND3_X1   g201(.A1(new_n587), .A2(new_n589), .A3(new_n590), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(G868), .ZN(G297));
  OAI21_X1  g203(.A(new_n626), .B1(new_n627), .B2(G868), .ZN(G280));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n623), .B1(new_n630), .B2(G860), .ZN(G148));
  NAND2_X1  g206(.A1(new_n623), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G868), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(G868), .B2(new_n579), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g210(.A(new_n485), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n636), .A2(new_n491), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n637), .B(new_n638), .Z(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(KEYINPUT13), .ZN(new_n641));
  AOI22_X1  g216(.A1(new_n640), .A2(new_n641), .B1(KEYINPUT84), .B2(G2100), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(new_n641), .B2(new_n640), .ZN(new_n643));
  NOR2_X1   g218(.A1(KEYINPUT84), .A2(G2100), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  AND2_X1   g220(.A1(new_n509), .A2(G123), .ZN(new_n646));
  INV_X1    g221(.A(G135), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n472), .A2(G111), .ZN(new_n648));
  OAI21_X1  g223(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n649));
  OAI22_X1  g224(.A1(new_n479), .A2(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OR3_X1    g225(.A1(new_n646), .A2(G2096), .A3(new_n650), .ZN(new_n651));
  OAI21_X1  g226(.A(G2096), .B1(new_n646), .B2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n645), .A2(new_n651), .A3(new_n652), .ZN(G156));
  INV_X1    g228(.A(KEYINPUT14), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2427), .B(G2438), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2430), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT15), .B(G2435), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n654), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n658), .B1(new_n657), .B2(new_n656), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2451), .B(G2454), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1341), .B(G1348), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n659), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2443), .B(G2446), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  AND3_X1   g242(.A1(new_n666), .A2(G14), .A3(new_n667), .ZN(G401));
  INV_X1    g243(.A(KEYINPUT18), .ZN(new_n669));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(KEYINPUT17), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n670), .A2(new_n671), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n669), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G2100), .ZN(new_n676));
  XOR2_X1   g251(.A(G2072), .B(G2078), .Z(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(new_n672), .B2(KEYINPUT18), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G2096), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n676), .B(new_n679), .ZN(G227));
  XNOR2_X1  g255(.A(G1956), .B(G2474), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT85), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1961), .B(G1966), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1971), .B(G1976), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT20), .Z(new_n689));
  OR2_X1    g264(.A1(new_n682), .A2(new_n684), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n690), .A2(new_n687), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n690), .A2(new_n687), .A3(new_n685), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n689), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G1991), .B(G1996), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(G229));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(KEYINPUT24), .B2(G34), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(KEYINPUT24), .B2(G34), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n497), .B2(G29), .ZN(new_n704));
  INV_X1    g279(.A(G2084), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT93), .Z(new_n707));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G5), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G171), .B2(new_n708), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n509), .A2(G129), .ZN(new_n711));
  NAND3_X1  g286(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT26), .Z(new_n713));
  INV_X1    g288(.A(G105), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n636), .B2(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n480), .B2(G141), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n718), .A2(new_n701), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n701), .B2(G32), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT27), .B(G1996), .ZN(new_n721));
  OAI221_X1 g296(.A(new_n707), .B1(G1961), .B2(new_n710), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT94), .ZN(new_n723));
  AND2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n722), .A2(new_n723), .ZN(new_n725));
  NOR2_X1   g300(.A1(G29), .A2(G33), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT89), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT25), .Z(new_n729));
  INV_X1    g304(.A(G139), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(new_n479), .B2(new_n730), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n731), .A2(KEYINPUT90), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n731), .A2(KEYINPUT90), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n513), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n734));
  OAI22_X1  g309(.A1(new_n732), .A2(new_n733), .B1(new_n472), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT91), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n727), .B1(new_n736), .B2(new_n701), .ZN(new_n737));
  INV_X1    g312(.A(G2072), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n701), .A2(G26), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT28), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n509), .A2(G128), .ZN(new_n742));
  OAI21_X1  g317(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n743));
  INV_X1    g318(.A(G116), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(G2105), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n480), .B2(G140), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n741), .B1(new_n748), .B2(new_n701), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT88), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G2067), .ZN(new_n751));
  NOR4_X1   g326(.A1(new_n724), .A2(new_n725), .A3(new_n739), .A4(new_n751), .ZN(new_n752));
  MUX2_X1   g327(.A(G6), .B(G305), .S(G16), .Z(new_n753));
  XOR2_X1   g328(.A(KEYINPUT32), .B(G1981), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n708), .A2(KEYINPUT86), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n708), .A2(KEYINPUT86), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n758), .A2(G22), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G166), .B2(new_n758), .ZN(new_n760));
  INV_X1    g335(.A(G1971), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n708), .A2(G23), .ZN(new_n763));
  INV_X1    g338(.A(G288), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(new_n708), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT33), .B(G1976), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n755), .A2(new_n762), .A3(new_n767), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT34), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n701), .A2(G25), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n509), .A2(G119), .ZN(new_n771));
  OAI21_X1  g346(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n772));
  INV_X1    g347(.A(G107), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(G2105), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n480), .B2(G131), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n770), .B1(new_n777), .B2(new_n701), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT35), .B(G1991), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  MUX2_X1   g355(.A(G24), .B(G290), .S(new_n758), .Z(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(G1986), .Z(new_n782));
  NAND3_X1  g357(.A1(new_n769), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT36), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n701), .A2(G35), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G162), .B2(new_n701), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT29), .Z(new_n787));
  INV_X1    g362(.A(G2090), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n701), .A2(G27), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G164), .B2(new_n701), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n789), .B1(G2078), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G2078), .B2(new_n791), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n787), .A2(new_n788), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n758), .A2(G19), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n579), .B2(new_n758), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT87), .B(G1341), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n708), .A2(G4), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n623), .B2(new_n708), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1348), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n646), .A2(new_n650), .ZN(new_n802));
  AOI211_X1 g377(.A(new_n798), .B(new_n801), .C1(G29), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n720), .A2(new_n721), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n704), .A2(new_n705), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n756), .A2(G20), .A3(new_n757), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT23), .Z(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G299), .B2(G16), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G1956), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT31), .B(G11), .Z(new_n810));
  INV_X1    g385(.A(G28), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n811), .A2(KEYINPUT30), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT92), .Z(new_n813));
  AOI21_X1  g388(.A(G29), .B1(new_n811), .B2(KEYINPUT30), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n810), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n708), .A2(G21), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G168), .B2(new_n708), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n815), .B1(new_n817), .B2(G1966), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(G1966), .B2(new_n817), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n809), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(G1961), .B2(new_n710), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n803), .A2(new_n804), .A3(new_n805), .A4(new_n821), .ZN(new_n822));
  AOI211_X1 g397(.A(new_n794), .B(new_n822), .C1(new_n738), .C2(new_n737), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n752), .A2(new_n784), .A3(new_n793), .A4(new_n823), .ZN(G150));
  INV_X1    g399(.A(G150), .ZN(G311));
  NAND2_X1  g400(.A1(G80), .A2(G543), .ZN(new_n826));
  INV_X1    g401(.A(G67), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n545), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n552), .B1(new_n828), .B2(KEYINPUT95), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(KEYINPUT95), .B2(new_n828), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n546), .A2(G93), .B1(new_n541), .B2(G55), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(G860), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT37), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n623), .A2(G559), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT38), .ZN(new_n836));
  NOR3_X1   g411(.A1(new_n832), .A2(new_n578), .A3(new_n576), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n579), .B1(new_n830), .B2(new_n831), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n836), .B(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT96), .Z(new_n844));
  INV_X1    g419(.A(G860), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(new_n841), .B2(new_n842), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n834), .B1(new_n844), .B2(new_n846), .ZN(G145));
  NAND2_X1  g422(.A1(new_n480), .A2(G142), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT99), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n851));
  INV_X1    g426(.A(G118), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n851), .B1(new_n852), .B2(G2105), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(new_n509), .B2(G130), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(new_n777), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT100), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n850), .A2(new_n776), .A3(new_n854), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n857), .B1(new_n856), .B2(new_n858), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n640), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n861), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n863), .A2(new_n639), .A3(new_n859), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(KEYINPUT101), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT97), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n523), .A2(KEYINPUT73), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n525), .B1(new_n504), .B2(new_n520), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n531), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n517), .B1(new_n511), .B2(KEYINPUT4), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n867), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n530), .B1(new_n524), .B2(new_n526), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n519), .A2(KEYINPUT97), .A3(new_n873), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n748), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT98), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n736), .A2(new_n877), .A3(new_n717), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n717), .B1(new_n736), .B2(new_n877), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n876), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n880), .ZN(new_n882));
  INV_X1    g457(.A(new_n876), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(new_n878), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT101), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n862), .A2(new_n864), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n866), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n887), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n889), .A2(new_n884), .A3(new_n881), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n802), .B(G162), .Z(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(G160), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(G37), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n888), .A2(new_n890), .A3(new_n893), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g474(.A(G868), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n832), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(G290), .B(G305), .ZN(new_n902));
  XNOR2_X1  g477(.A(G166), .B(new_n764), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n902), .B(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT42), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n905), .A2(KEYINPUT104), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n632), .B(new_n839), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT102), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n627), .A2(new_n908), .ZN(new_n909));
  OAI211_X1 g484(.A(new_n617), .B(new_n621), .C1(G299), .C2(KEYINPUT102), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n623), .A2(new_n908), .A3(new_n627), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(KEYINPUT103), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n915), .B1(new_n911), .B2(new_n912), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n907), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n913), .A2(KEYINPUT41), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT41), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n919), .B1(new_n911), .B2(new_n912), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n917), .B1(new_n907), .B2(new_n921), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n906), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n906), .A2(new_n922), .ZN(new_n924));
  AOI22_X1  g499(.A1(new_n923), .A2(new_n924), .B1(KEYINPUT104), .B2(new_n905), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n901), .B1(new_n925), .B2(new_n900), .ZN(G295));
  NAND2_X1  g501(.A1(G295), .A2(KEYINPUT105), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT105), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n928), .B(new_n901), .C1(new_n925), .C2(new_n900), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(G331));
  INV_X1    g505(.A(new_n904), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n914), .A2(new_n916), .ZN(new_n932));
  NOR2_X1   g507(.A1(G171), .A2(G168), .ZN(new_n933));
  NOR2_X1   g508(.A1(G286), .A2(G301), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT107), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(new_n936), .A3(new_n839), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n839), .ZN(new_n938));
  OAI22_X1  g513(.A1(new_n933), .A2(new_n934), .B1(new_n837), .B2(new_n838), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(new_n939), .A3(KEYINPUT107), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n932), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n938), .A2(new_n939), .A3(new_n942), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n840), .B(KEYINPUT108), .C1(new_n933), .C2(new_n934), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n921), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n931), .B1(new_n941), .B2(new_n946), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n918), .A2(new_n920), .A3(new_n940), .A4(new_n937), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n945), .A2(new_n913), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(new_n949), .A3(new_n904), .ZN(new_n950));
  AOI21_X1  g525(.A(G37), .B1(new_n950), .B2(KEYINPUT109), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n948), .A2(new_n949), .A3(new_n952), .A4(new_n904), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n947), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n948), .A2(new_n949), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n931), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n951), .A2(new_n953), .A3(new_n957), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n955), .B(KEYINPUT44), .C1(KEYINPUT43), .C2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT43), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n947), .A2(new_n951), .A3(new_n961), .A4(new_n953), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n959), .B1(new_n963), .B2(new_n964), .ZN(G397));
  INV_X1    g540(.A(KEYINPUT119), .ZN(new_n966));
  INV_X1    g541(.A(G8), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT50), .ZN(new_n968));
  INV_X1    g543(.A(G1384), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n535), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n481), .A2(new_n496), .A3(G40), .A4(new_n487), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n519), .A2(new_n873), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n969), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n971), .B1(new_n973), .B2(KEYINPUT50), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n970), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT118), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n970), .A2(new_n974), .A3(KEYINPUT118), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(new_n788), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n535), .A2(new_n969), .ZN(new_n980));
  XNOR2_X1  g555(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n971), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n983), .A2(G1384), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n872), .A2(new_n874), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT112), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n872), .A2(new_n874), .A3(KEYINPUT112), .A4(new_n984), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n982), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n761), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n967), .B1(new_n979), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n593), .A2(G8), .A3(new_n595), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT55), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n966), .B1(new_n992), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n997), .B(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(G1971), .B1(new_n982), .B2(new_n989), .ZN(new_n1001));
  AOI21_X1  g576(.A(G1384), .B1(new_n519), .B2(new_n873), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n971), .B1(new_n1002), .B2(new_n968), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n870), .A2(new_n533), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n873), .A2(KEYINPUT74), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(G1384), .B1(new_n1006), .B2(new_n519), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1003), .B1(new_n1007), .B2(new_n968), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1008), .A2(G2090), .ZN(new_n1009));
  OAI211_X1 g584(.A(G8), .B(new_n1000), .C1(new_n1001), .C2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n973), .A2(new_n971), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1011), .A2(new_n967), .ZN(new_n1012));
  OR3_X1    g587(.A1(G305), .A2(KEYINPUT115), .A3(G1981), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT115), .B1(G305), .B2(G1981), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n606), .B1(new_n601), .B2(new_n547), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(G1981), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(KEYINPUT116), .A2(KEYINPUT49), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1015), .B(new_n1017), .C1(KEYINPUT116), .C2(KEYINPUT49), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1012), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n764), .A2(G1976), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1023), .B(KEYINPUT114), .ZN(new_n1024));
  INV_X1    g599(.A(G1976), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT52), .B1(G288), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1012), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1022), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1029), .B1(new_n1012), .B2(new_n1024), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n1010), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n968), .B1(new_n535), .B2(new_n969), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n972), .A2(new_n968), .A3(new_n969), .ZN(new_n1034));
  INV_X1    g609(.A(new_n971), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n1033), .A2(G2084), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n981), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n535), .A2(new_n969), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n971), .B1(new_n973), .B2(new_n983), .ZN(new_n1040));
  AOI21_X1  g615(.A(G1966), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(G8), .B1(new_n1037), .B2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1042), .A2(G286), .ZN(new_n1043));
  INV_X1    g618(.A(new_n997), .ZN(new_n1044));
  AOI21_X1  g619(.A(G2090), .B1(new_n975), .B2(new_n976), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n1045), .A2(new_n978), .B1(new_n990), .B2(new_n761), .ZN(new_n1046));
  OAI211_X1 g621(.A(KEYINPUT119), .B(new_n1044), .C1(new_n1046), .C2(new_n967), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n998), .A2(new_n1032), .A3(new_n1043), .A4(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT63), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(G8), .B1(new_n1001), .B2(new_n1009), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n1044), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n1042), .A2(new_n1049), .A3(G286), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1032), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT120), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1032), .A2(KEYINPUT120), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1050), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g633(.A(KEYINPUT56), .B(G2072), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n982), .A2(new_n989), .A3(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n627), .B(KEYINPUT57), .ZN(new_n1061));
  INV_X1    g636(.A(G1956), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n975), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1060), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n973), .A2(G2067), .A3(new_n971), .ZN(new_n1065));
  INV_X1    g640(.A(G1348), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1065), .B1(new_n1008), .B2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1067), .A2(new_n622), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1061), .B1(new_n1060), .B2(new_n1063), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1064), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT60), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1066), .B1(new_n1033), .B2(new_n1036), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1065), .ZN(new_n1073));
  AND4_X1   g648(.A1(new_n1071), .A2(new_n1072), .A3(new_n623), .A4(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1071), .B1(new_n1067), .B2(new_n623), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n622), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1074), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G1996), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n982), .A2(new_n989), .A3(new_n1079), .ZN(new_n1080));
  XOR2_X1   g655(.A(KEYINPUT58), .B(G1341), .Z(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(new_n973), .B2(new_n971), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n579), .ZN(new_n1084));
  OR2_X1    g659(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1085));
  NAND2_X1  g660(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1061), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1090), .A2(KEYINPUT61), .A3(new_n1064), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1083), .A2(KEYINPUT121), .A3(KEYINPUT59), .A4(new_n579), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1078), .A2(new_n1087), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1060), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1094), .A2(new_n1069), .A3(KEYINPUT122), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1088), .A2(KEYINPUT122), .A3(new_n1089), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT61), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1070), .B1(new_n1093), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n998), .A2(new_n1032), .A3(new_n1047), .ZN(new_n1101));
  INV_X1    g676(.A(G2078), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n982), .A2(new_n989), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT53), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1035), .B1(new_n1002), .B2(KEYINPUT45), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1106), .B1(new_n1007), .B2(new_n1038), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1107), .A2(KEYINPUT53), .A3(new_n1102), .ZN(new_n1108));
  INV_X1    g683(.A(G1961), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1008), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1105), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(G301), .B(KEYINPUT54), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1103), .A2(new_n1104), .B1(new_n1109), .B2(new_n1008), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1038), .B1(new_n875), .B2(new_n969), .ZN(new_n1114));
  OR2_X1    g689(.A1(new_n488), .A2(KEYINPUT124), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n488), .A2(KEYINPUT124), .ZN(new_n1116));
  AND4_X1   g691(.A1(KEYINPUT53), .A2(new_n494), .A3(G40), .A4(new_n1102), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1112), .B1(new_n1119), .B2(new_n989), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1111), .A2(new_n1112), .B1(new_n1113), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT51), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n705), .B(new_n1003), .C1(new_n1007), .C2(new_n968), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n1107), .B2(G1966), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1122), .B(G8), .C1(new_n1124), .C2(G286), .ZN(new_n1125));
  NOR2_X1   g700(.A1(G168), .A2(new_n967), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1042), .A2(KEYINPUT51), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT123), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1129), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1131));
  INV_X1    g706(.A(G1966), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  AOI211_X1 g708(.A(KEYINPUT123), .B(new_n1127), .C1(new_n1133), .C2(new_n1123), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1125), .B(new_n1128), .C1(new_n1130), .C2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1121), .A2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1101), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1100), .A2(new_n1137), .ZN(new_n1138));
  OR2_X1    g713(.A1(new_n1135), .A2(KEYINPUT62), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1111), .A2(G171), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1140), .B1(new_n1135), .B2(KEYINPUT62), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1032), .A2(new_n1047), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1139), .A2(new_n1141), .A3(new_n998), .A4(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(G288), .A2(G1976), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1022), .A2(new_n1144), .B1(new_n1014), .B2(new_n1013), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1145), .A2(KEYINPUT117), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n1146), .A2(new_n967), .A3(new_n1011), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(KEYINPUT117), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1010), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1147), .A2(new_n1148), .B1(new_n1149), .B2(new_n1031), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1058), .A2(new_n1138), .A3(new_n1143), .A4(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1114), .A2(new_n1035), .ZN(new_n1152));
  OR3_X1    g727(.A1(new_n1152), .A2(G1986), .A3(G290), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1152), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1154), .A2(G1986), .A3(G290), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1156), .B(KEYINPUT111), .ZN(new_n1157));
  XOR2_X1   g732(.A(new_n747), .B(G2067), .Z(new_n1158));
  XNOR2_X1  g733(.A(new_n717), .B(new_n1079), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n776), .B(new_n779), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1152), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1157), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1151), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n777), .A2(new_n779), .ZN(new_n1166));
  OAI22_X1  g741(.A1(new_n1160), .A2(new_n1166), .B1(G2067), .B2(new_n747), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(new_n1154), .ZN(new_n1168));
  OR2_X1    g743(.A1(new_n1168), .A2(KEYINPUT125), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(KEYINPUT125), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT48), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1163), .B1(new_n1171), .B2(new_n1153), .ZN(new_n1172));
  OR2_X1    g747(.A1(new_n1153), .A2(new_n1171), .ZN(new_n1173));
  AOI22_X1  g748(.A1(new_n1169), .A2(new_n1170), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1152), .B1(new_n718), .B2(new_n1158), .ZN(new_n1175));
  OR3_X1    g750(.A1(new_n1152), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1176));
  OAI21_X1  g751(.A(KEYINPUT46), .B1(new_n1152), .B2(G1996), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1175), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT47), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1174), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT126), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1182), .B(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1165), .A2(new_n1184), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g760(.A1(G401), .A2(new_n461), .A3(G227), .ZN(new_n1187));
  NAND2_X1  g761(.A1(new_n699), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g762(.A(new_n1188), .B1(new_n960), .B2(new_n962), .ZN(new_n1189));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n1190));
  AOI21_X1  g764(.A(new_n893), .B1(new_n888), .B2(new_n890), .ZN(new_n1191));
  NAND2_X1  g765(.A1(new_n897), .A2(new_n896), .ZN(new_n1192));
  OAI211_X1 g766(.A(new_n1189), .B(new_n1190), .C1(new_n1191), .C2(new_n1192), .ZN(new_n1193));
  INV_X1    g767(.A(new_n1193), .ZN(new_n1194));
  AOI21_X1  g768(.A(new_n1190), .B1(new_n898), .B2(new_n1189), .ZN(new_n1195));
  NOR2_X1   g769(.A1(new_n1194), .A2(new_n1195), .ZN(G308));
  NAND2_X1  g770(.A1(new_n898), .A2(new_n1189), .ZN(G225));
endmodule


