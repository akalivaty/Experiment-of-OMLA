//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 1 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n623,
    new_n626, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1211, new_n1212, new_n1213, new_n1214;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XNOR2_X1  g016(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(new_n454), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT70), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(KEYINPUT70), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n465), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(G101), .A2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(KEYINPUT71), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT71), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n474), .B(new_n464), .C1(new_n470), .C2(new_n471), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  AND2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NOR2_X1   g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  OAI21_X1  g053(.A(G125), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g056(.A(KEYINPUT68), .B(G125), .C1(new_n477), .C2(new_n478), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(G113), .A2(G2104), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n485), .A2(new_n486), .A3(G2105), .ZN(new_n487));
  INV_X1    g062(.A(new_n484), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(new_n481), .B2(new_n482), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT69), .B1(new_n489), .B2(new_n464), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n476), .B1(new_n487), .B2(new_n490), .ZN(G160));
  OR2_X1    g066(.A1(G100), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n493));
  AND3_X1   g068(.A1(KEYINPUT70), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n494));
  AOI21_X1  g069(.A(KEYINPUT3), .B1(KEYINPUT70), .B2(G2104), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT73), .ZN(new_n497));
  NOR3_X1   g072(.A1(new_n496), .A2(new_n497), .A3(new_n464), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n468), .A2(new_n469), .ZN(new_n499));
  AOI21_X1  g074(.A(KEYINPUT73), .B1(new_n499), .B2(G2105), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G124), .ZN(new_n502));
  INV_X1    g077(.A(G136), .ZN(new_n503));
  NOR3_X1   g078(.A1(new_n496), .A2(KEYINPUT72), .A3(G2105), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n505), .B1(new_n499), .B2(new_n464), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  OAI221_X1 g082(.A(new_n493), .B1(new_n501), .B2(new_n502), .C1(new_n503), .C2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G162));
  XNOR2_X1  g084(.A(KEYINPUT3), .B(G2104), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n510), .A2(G138), .A3(new_n464), .ZN(new_n511));
  OAI21_X1  g086(.A(G126), .B1(new_n494), .B2(new_n495), .ZN(new_n512));
  NAND2_X1  g087(.A1(G114), .A2(G2104), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n464), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT4), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n511), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OAI211_X1 g091(.A(KEYINPUT4), .B(G138), .C1(new_n494), .C2(new_n495), .ZN(new_n517));
  NAND2_X1  g092(.A1(G102), .A2(G2104), .ZN(new_n518));
  AOI21_X1  g093(.A(G2105), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(G164));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT5), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT5), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G62), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n523), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G651), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT74), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AND2_X1   g108(.A1(KEYINPUT6), .A2(G651), .ZN(new_n534));
  NOR2_X1   g109(.A1(KEYINPUT6), .A2(G651), .ZN(new_n535));
  OAI211_X1 g110(.A(G50), .B(G543), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  OAI211_X1 g111(.A(new_n525), .B(new_n527), .C1(new_n534), .C2(new_n535), .ZN(new_n537));
  INV_X1    g112(.A(G88), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n530), .A2(KEYINPUT74), .A3(G651), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n533), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT75), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n533), .A2(KEYINPUT75), .A3(new_n540), .A4(new_n541), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(G166));
  NAND3_X1  g121(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT76), .ZN(new_n548));
  XOR2_X1   g123(.A(new_n548), .B(KEYINPUT7), .Z(new_n549));
  NOR2_X1   g124(.A1(new_n534), .A2(new_n535), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n524), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G51), .ZN(new_n552));
  INV_X1    g127(.A(new_n550), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n553), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n552), .B1(new_n554), .B2(new_n528), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n549), .A2(new_n555), .ZN(G168));
  INV_X1    g131(.A(new_n528), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n557), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G651), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n553), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G52), .ZN(new_n562));
  INV_X1    g137(.A(G90), .ZN(new_n563));
  OAI22_X1  g138(.A1(new_n561), .A2(new_n562), .B1(new_n563), .B2(new_n537), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n560), .A2(new_n564), .ZN(G171));
  AOI22_X1  g140(.A1(new_n557), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n566), .A2(new_n559), .ZN(new_n567));
  INV_X1    g142(.A(G43), .ZN(new_n568));
  INV_X1    g143(.A(G81), .ZN(new_n569));
  OAI22_X1  g144(.A1(new_n561), .A2(new_n568), .B1(new_n569), .B2(new_n537), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G860), .ZN(G153));
  AND3_X1   g147(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G36), .ZN(G176));
  NAND2_X1  g149(.A1(G1), .A2(G3), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT77), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT8), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT78), .ZN(G188));
  NAND2_X1  g154(.A1(new_n551), .A2(G53), .ZN(new_n580));
  XOR2_X1   g155(.A(new_n580), .B(KEYINPUT9), .Z(new_n581));
  INV_X1    g156(.A(new_n537), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G91), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n557), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n584), .B2(new_n559), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n581), .A2(new_n585), .ZN(G299));
  INV_X1    g161(.A(G171), .ZN(G301));
  INV_X1    g162(.A(G168), .ZN(G286));
  INV_X1    g163(.A(G166), .ZN(G303));
  NAND2_X1  g164(.A1(new_n551), .A2(G49), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT79), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n557), .A2(G74), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n592), .A2(G651), .B1(G87), .B2(new_n582), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n591), .A2(new_n593), .ZN(G288));
  AOI22_X1  g169(.A1(new_n557), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n595), .A2(new_n559), .ZN(new_n596));
  INV_X1    g171(.A(G48), .ZN(new_n597));
  INV_X1    g172(.A(G86), .ZN(new_n598));
  OAI22_X1  g173(.A1(new_n561), .A2(new_n597), .B1(new_n598), .B2(new_n537), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G305));
  AOI22_X1  g176(.A1(new_n557), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(new_n559), .ZN(new_n603));
  INV_X1    g178(.A(G47), .ZN(new_n604));
  INV_X1    g179(.A(G85), .ZN(new_n605));
  OAI22_X1  g180(.A1(new_n561), .A2(new_n604), .B1(new_n605), .B2(new_n537), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(G290));
  NAND2_X1  g183(.A1(G301), .A2(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n528), .B2(new_n611), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT81), .Z(new_n613));
  AOI22_X1  g188(.A1(new_n613), .A2(G651), .B1(G54), .B2(new_n551), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n582), .A2(G92), .ZN(new_n615));
  XOR2_X1   g190(.A(KEYINPUT80), .B(KEYINPUT10), .Z(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n609), .B1(new_n619), .B2(G868), .ZN(G284));
  OAI21_X1  g195(.A(new_n609), .B1(new_n619), .B2(G868), .ZN(G321));
  NAND2_X1  g196(.A1(G286), .A2(G868), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n581), .A2(new_n585), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G868), .ZN(G297));
  OAI21_X1  g199(.A(new_n622), .B1(new_n623), .B2(G868), .ZN(G280));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n619), .B1(new_n626), .B2(G860), .ZN(G148));
  NAND2_X1  g202(.A1(new_n619), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G868), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(G868), .B2(new_n571), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g206(.A1(new_n498), .A2(new_n500), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G123), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n504), .A2(new_n506), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(G135), .ZN(new_n635));
  OR2_X1    g210(.A1(G99), .A2(G2105), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n636), .B(G2104), .C1(G111), .C2(new_n464), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n633), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT82), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2096), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT13), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2100), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n640), .A2(new_n644), .ZN(G156));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2435), .ZN(new_n647));
  XOR2_X1   g222(.A(G2427), .B(G2438), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(KEYINPUT14), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2451), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n652), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G1341), .B(G1348), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n659), .A2(KEYINPUT84), .ZN(new_n660));
  INV_X1    g235(.A(G14), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n656), .B2(new_n658), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n659), .A2(KEYINPUT84), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n660), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(G401));
  XOR2_X1   g240(.A(G2072), .B(G2078), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT85), .ZN(new_n667));
  XOR2_X1   g242(.A(G2067), .B(G2678), .Z(new_n668));
  XNOR2_X1  g243(.A(G2084), .B(G2090), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT18), .Z(new_n672));
  NAND2_X1  g247(.A1(new_n668), .A2(new_n669), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n667), .B(KEYINPUT86), .ZN(new_n674));
  INV_X1    g249(.A(new_n670), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(new_n673), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n667), .B(KEYINPUT17), .ZN(new_n677));
  OAI221_X1 g252(.A(new_n672), .B1(new_n673), .B2(new_n674), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G2096), .ZN(new_n679));
  INV_X1    g254(.A(G2100), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(G227));
  XOR2_X1   g256(.A(G1956), .B(G2474), .Z(new_n682));
  XOR2_X1   g257(.A(G1961), .B(G1966), .Z(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1971), .B(G1976), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n682), .A2(new_n683), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT20), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n688), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n685), .A2(new_n687), .A3(new_n689), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n692), .B(new_n693), .C1(new_n691), .C2(new_n690), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT21), .B(G1986), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1991), .B(G1996), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT22), .B(G1981), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n700), .B(new_n701), .Z(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(G229));
  NAND2_X1  g278(.A1(new_n634), .A2(G139), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT25), .Z(new_n706));
  AOI22_X1  g281(.A1(new_n510), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT98), .Z(new_n708));
  OAI211_X1 g283(.A(new_n704), .B(new_n706), .C1(new_n708), .C2(new_n464), .ZN(new_n709));
  MUX2_X1   g284(.A(G33), .B(new_n709), .S(G29), .Z(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT99), .Z(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G2072), .ZN(new_n712));
  INV_X1    g287(.A(G29), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n713), .A2(G35), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(new_n508), .B2(G29), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT29), .ZN(new_n716));
  INV_X1    g291(.A(G2090), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n712), .A2(new_n718), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n716), .A2(new_n717), .ZN(new_n720));
  INV_X1    g295(.A(G16), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G19), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(new_n571), .B2(new_n721), .ZN(new_n723));
  MUX2_X1   g298(.A(new_n722), .B(new_n723), .S(KEYINPUT95), .Z(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(G1341), .Z(new_n725));
  NOR2_X1   g300(.A1(G5), .A2(G16), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G171), .B2(G16), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G1961), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n634), .A2(G141), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n632), .A2(G129), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n464), .A2(G105), .A3(G2104), .ZN(new_n731));
  NAND3_X1  g306(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT26), .Z(new_n733));
  NAND4_X1  g308(.A1(new_n729), .A2(new_n730), .A3(new_n731), .A4(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G29), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G29), .B2(G32), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT27), .B(G1996), .ZN(new_n738));
  INV_X1    g313(.A(G1966), .ZN(new_n739));
  NAND2_X1  g314(.A1(G168), .A2(G16), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G16), .B2(G21), .ZN(new_n741));
  AOI22_X1  g316(.A1(new_n737), .A2(new_n738), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n720), .A2(new_n725), .A3(new_n728), .A4(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n741), .A2(new_n739), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT100), .ZN(new_n745));
  INV_X1    g320(.A(new_n638), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G29), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n745), .B(new_n747), .C1(new_n737), .C2(new_n738), .ZN(new_n748));
  NOR3_X1   g323(.A1(new_n719), .A2(new_n743), .A3(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT31), .B(G11), .ZN(new_n750));
  NOR2_X1   g325(.A1(G27), .A2(G29), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G164), .B2(G29), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G2078), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n721), .A2(KEYINPUT23), .A3(G20), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT23), .ZN(new_n755));
  INV_X1    g330(.A(G20), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n756), .B2(G16), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n754), .B(new_n757), .C1(new_n623), .C2(new_n721), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G1956), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT30), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n760), .A2(G28), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n760), .A2(G28), .ZN(new_n762));
  NOR3_X1   g337(.A1(new_n761), .A2(new_n762), .A3(G29), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT24), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n765), .A2(G34), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(G34), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n766), .A2(new_n767), .A3(new_n713), .ZN(new_n768));
  INV_X1    g343(.A(G160), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n769), .B2(new_n713), .ZN(new_n770));
  INV_X1    g345(.A(G2084), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n713), .A2(G26), .ZN(new_n774));
  OR3_X1    g349(.A1(KEYINPUT96), .A2(G104), .A3(G2105), .ZN(new_n775));
  INV_X1    g350(.A(G116), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n776), .A2(G2105), .ZN(new_n777));
  OAI21_X1  g352(.A(KEYINPUT96), .B1(G104), .B2(G2105), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n775), .A2(G2104), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT97), .ZN(new_n780));
  OAI21_X1  g355(.A(G128), .B1(new_n498), .B2(new_n500), .ZN(new_n781));
  OAI21_X1  g356(.A(G140), .B1(new_n504), .B2(new_n506), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n774), .B1(new_n784), .B2(new_n713), .ZN(new_n785));
  MUX2_X1   g360(.A(new_n774), .B(new_n785), .S(KEYINPUT28), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(G2067), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n764), .A2(new_n772), .A3(new_n773), .A4(new_n787), .ZN(new_n788));
  OAI22_X1  g363(.A1(new_n711), .A2(G2072), .B1(G2078), .B2(new_n752), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n749), .A2(new_n750), .A3(new_n753), .A4(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n721), .B1(new_n591), .B2(new_n593), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n721), .A2(G23), .ZN(new_n793));
  OR3_X1    g368(.A1(new_n792), .A2(KEYINPUT91), .A3(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(KEYINPUT91), .B1(new_n792), .B2(new_n793), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT33), .B(G1976), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT92), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n796), .B(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(G16), .A2(G22), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G166), .B2(G16), .ZN(new_n801));
  INV_X1    g376(.A(G1971), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n721), .A2(G6), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n600), .B2(new_n721), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT32), .B(G1981), .Z(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n799), .A2(new_n803), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(KEYINPUT34), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT34), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n799), .A2(new_n810), .A3(new_n803), .A4(new_n807), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(KEYINPUT93), .A2(KEYINPUT36), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n713), .A2(G25), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n632), .A2(G119), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n634), .A2(G131), .ZN(new_n816));
  OR2_X1    g391(.A1(G95), .A2(G2105), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n817), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n815), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n814), .B1(new_n820), .B2(new_n713), .ZN(new_n821));
  MUX2_X1   g396(.A(new_n814), .B(new_n821), .S(KEYINPUT87), .Z(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT35), .B(G1991), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n822), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n721), .A2(G24), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT88), .Z(new_n827));
  XOR2_X1   g402(.A(new_n607), .B(KEYINPUT89), .Z(new_n828));
  OAI21_X1  g403(.A(new_n827), .B1(new_n828), .B2(new_n721), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT90), .B(G1986), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n812), .A2(new_n813), .A3(new_n825), .A4(new_n831), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n809), .A2(new_n811), .A3(new_n825), .A4(new_n831), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n833), .A2(KEYINPUT93), .A3(KEYINPUT36), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n791), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n786), .A2(G2067), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n727), .A2(G1961), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n721), .A2(G4), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(new_n619), .B2(new_n721), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT94), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(G1348), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n835), .A2(new_n836), .A3(new_n837), .A4(new_n841), .ZN(G150));
  INV_X1    g417(.A(G150), .ZN(G311));
  NAND2_X1  g418(.A1(G80), .A2(G543), .ZN(new_n844));
  INV_X1    g419(.A(G67), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n844), .B1(new_n528), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(G651), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(KEYINPUT101), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n582), .A2(G93), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n551), .A2(G55), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT101), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n846), .A2(new_n851), .A3(G651), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n848), .A2(new_n849), .A3(new_n850), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(G860), .ZN(new_n854));
  XOR2_X1   g429(.A(KEYINPUT103), .B(KEYINPUT37), .Z(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT104), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n854), .B(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n618), .A2(new_n626), .ZN(new_n858));
  XNOR2_X1  g433(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT39), .Z(new_n861));
  OR2_X1    g436(.A1(new_n853), .A2(new_n571), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n853), .A2(new_n571), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n861), .B(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n857), .B1(new_n865), .B2(G860), .ZN(G145));
  AOI22_X1  g441(.A1(G130), .A2(new_n632), .B1(new_n634), .B2(G142), .ZN(new_n867));
  NOR2_X1   g442(.A1(G106), .A2(G2105), .ZN(new_n868));
  OAI21_X1  g443(.A(G2104), .B1(new_n464), .B2(G118), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n642), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n521), .A2(KEYINPUT106), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT106), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n516), .A2(new_n873), .A3(new_n520), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n735), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n734), .B1(new_n872), .B2(new_n874), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n784), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NOR3_X1   g454(.A1(new_n876), .A2(new_n877), .A3(new_n784), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n709), .A2(KEYINPUT107), .ZN(new_n881));
  NOR3_X1   g456(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n709), .A2(KEYINPUT107), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n881), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n876), .A2(new_n877), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n783), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n884), .B1(new_n886), .B2(new_n878), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n871), .B1(new_n882), .B2(new_n887), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n881), .B(new_n883), .C1(new_n879), .C2(new_n880), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n886), .A2(KEYINPUT107), .A3(new_n709), .A4(new_n878), .ZN(new_n890));
  INV_X1    g465(.A(new_n871), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n508), .A2(KEYINPUT105), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n508), .A2(KEYINPUT105), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n894), .A2(new_n638), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n638), .B1(new_n894), .B2(new_n895), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n769), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n894), .A2(new_n895), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n746), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n901), .A2(new_n896), .A3(G160), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n899), .A2(new_n819), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n819), .B1(new_n899), .B2(new_n902), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n893), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(G37), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n888), .B(new_n892), .C1(new_n904), .C2(new_n903), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(KEYINPUT108), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT108), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n906), .A2(new_n908), .A3(new_n911), .A4(new_n907), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT40), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n910), .A2(KEYINPUT40), .A3(new_n912), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(G395));
  XNOR2_X1  g492(.A(G166), .B(G290), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(new_n600), .ZN(new_n919));
  INV_X1    g494(.A(G288), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n918), .A2(G305), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n918), .A2(G305), .ZN(new_n923));
  OAI21_X1  g498(.A(G288), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g500(.A(new_n925), .B(KEYINPUT42), .Z(new_n926));
  XNOR2_X1  g501(.A(new_n628), .B(new_n864), .ZN(new_n927));
  NAND2_X1  g502(.A1(G299), .A2(KEYINPUT109), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT109), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n623), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n928), .A2(new_n618), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n619), .A2(new_n929), .A3(new_n623), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n927), .A2(new_n933), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n931), .A2(KEYINPUT41), .A3(new_n932), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT41), .B1(new_n931), .B2(new_n932), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n934), .B1(new_n937), .B2(new_n927), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n926), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n926), .A2(new_n938), .ZN(new_n940));
  OAI21_X1  g515(.A(G868), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(G868), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n853), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(G295));
  NAND2_X1  g519(.A1(new_n941), .A2(new_n943), .ZN(G331));
  NAND3_X1  g520(.A1(new_n862), .A2(G301), .A3(new_n863), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(G301), .B1(new_n862), .B2(new_n863), .ZN(new_n948));
  OAI21_X1  g523(.A(G286), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n948), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n950), .A2(G168), .A3(new_n946), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n952), .B1(new_n935), .B2(new_n936), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n933), .A2(new_n949), .A3(new_n951), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n925), .A2(new_n953), .A3(KEYINPUT110), .A4(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n953), .A2(KEYINPUT110), .A3(new_n954), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n956), .A2(new_n921), .A3(new_n924), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n955), .A2(new_n957), .A3(new_n907), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n955), .A2(new_n957), .A3(new_n960), .A4(new_n907), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT44), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n959), .A2(KEYINPUT44), .A3(new_n961), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(G397));
  INV_X1    g541(.A(G1981), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n600), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT49), .ZN(new_n969));
  OAI21_X1  g544(.A(G1981), .B1(new_n596), .B2(new_n599), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n969), .B1(new_n968), .B2(new_n970), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  XOR2_X1   g549(.A(KEYINPUT117), .B(G8), .Z(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G1384), .ZN(new_n977));
  INV_X1    g552(.A(new_n511), .ZN(new_n978));
  INV_X1    g553(.A(G126), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n979), .B1(new_n468), .B2(new_n469), .ZN(new_n980));
  INV_X1    g555(.A(new_n513), .ZN(new_n981));
  OAI21_X1  g556(.A(G2105), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n978), .B1(new_n982), .B2(KEYINPUT4), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n977), .B1(new_n983), .B2(new_n519), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT115), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n521), .A2(KEYINPUT115), .A3(new_n977), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G40), .ZN(new_n989));
  AOI211_X1 g564(.A(new_n989), .B(new_n476), .C1(new_n490), .C2(new_n487), .ZN(new_n990));
  AOI211_X1 g565(.A(KEYINPUT118), .B(new_n976), .C1(new_n988), .C2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT118), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT115), .B1(new_n521), .B2(new_n977), .ZN(new_n993));
  AOI211_X1 g568(.A(new_n985), .B(G1384), .C1(new_n516), .C2(new_n520), .ZN(new_n994));
  OAI211_X1 g569(.A(G40), .B(G160), .C1(new_n993), .C2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n992), .B1(new_n995), .B2(new_n975), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n974), .B1(new_n991), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT119), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n473), .A2(new_n475), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n486), .B1(new_n485), .B2(G2105), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n489), .A2(KEYINPUT69), .A3(new_n464), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n999), .B(G40), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1002), .B1(new_n986), .B2(new_n987), .ZN(new_n1003));
  OAI21_X1  g578(.A(KEYINPUT118), .B1(new_n1003), .B2(new_n976), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n995), .A2(new_n992), .A3(new_n975), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT119), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1006), .A2(new_n1007), .A3(new_n974), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n998), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n874), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n873), .B1(new_n516), .B2(new_n520), .ZN(new_n1011));
  OAI211_X1 g586(.A(KEYINPUT45), .B(new_n977), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT45), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n984), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1012), .A2(new_n990), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n802), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1017), .B1(new_n521), .B2(new_n977), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1002), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1017), .B1(new_n993), .B2(new_n994), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1016), .B1(G2090), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(G8), .ZN(new_n1023));
  NAND2_X1  g598(.A1(G303), .A2(G8), .ZN(new_n1024));
  XNOR2_X1  g599(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n1024), .B(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n920), .A2(G1976), .ZN(new_n1028));
  INV_X1    g603(.A(G1976), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT52), .B1(G288), .B2(new_n1029), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1028), .B(new_n1030), .C1(new_n991), .C2(new_n996), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1028), .B1(new_n991), .B2(new_n996), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT52), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1009), .A2(new_n1027), .A3(new_n1031), .A4(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n968), .ZN(new_n1035));
  NOR2_X1   g610(.A1(G288), .A2(G1976), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1035), .B1(new_n1009), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1006), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1034), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  XOR2_X1   g614(.A(new_n1024), .B(new_n1025), .Z(new_n1040));
  NAND3_X1  g615(.A1(new_n1040), .A2(G8), .A3(new_n1022), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1009), .A2(new_n1041), .A3(new_n1031), .A4(new_n1033), .ZN(new_n1042));
  XOR2_X1   g617(.A(KEYINPUT121), .B(G2084), .Z(new_n1043));
  AND3_X1   g618(.A1(new_n1019), .A2(new_n1020), .A3(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n984), .A2(new_n1013), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1002), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n986), .A2(new_n1013), .A3(new_n987), .ZN(new_n1047));
  AOI21_X1  g622(.A(G1966), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G8), .ZN(new_n1049));
  NOR2_X1   g624(.A1(G168), .A2(new_n976), .ZN(new_n1050));
  OAI22_X1  g625(.A1(new_n1044), .A2(new_n1048), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n993), .A2(new_n994), .A3(KEYINPUT45), .ZN(new_n1052));
  OAI211_X1 g627(.A(G160), .B(G40), .C1(new_n1013), .C2(new_n984), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n739), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1019), .A2(new_n1020), .A3(new_n1043), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1054), .B(new_n1055), .C1(G168), .C2(new_n976), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1051), .A2(new_n1056), .A3(KEYINPUT51), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n975), .B1(new_n1044), .B2(new_n1048), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1050), .A2(KEYINPUT51), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1057), .A2(new_n1060), .A3(KEYINPUT62), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n986), .A2(KEYINPUT50), .A3(new_n987), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n990), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n984), .A2(KEYINPUT50), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1062), .A2(KEYINPUT120), .A3(new_n990), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1065), .A2(new_n717), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n1016), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1040), .B1(new_n1070), .B2(new_n975), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1042), .A2(new_n1061), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G2078), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1012), .A2(new_n990), .A3(new_n1073), .A4(new_n1014), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G1961), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1021), .A2(new_n1077), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1075), .A2(G2078), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1046), .A2(new_n1080), .A3(new_n1047), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(G171), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT62), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1083), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1039), .B1(new_n1072), .B2(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g662(.A(new_n623), .B(KEYINPUT57), .ZN(new_n1088));
  XOR2_X1   g663(.A(KEYINPUT56), .B(G2072), .Z(new_n1089));
  NOR2_X1   g664(.A1(new_n1015), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1062), .A2(KEYINPUT120), .A3(new_n990), .ZN(new_n1092));
  AOI21_X1  g667(.A(KEYINPUT120), .B1(new_n1062), .B2(new_n990), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1092), .A2(new_n1093), .A3(new_n1066), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1088), .B(new_n1091), .C1(new_n1094), .C2(G1956), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1065), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1096));
  INV_X1    g671(.A(G1956), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1090), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1098), .A2(new_n1088), .ZN(new_n1099));
  INV_X1    g674(.A(G1348), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1021), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(G2067), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1003), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n618), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1095), .B1(new_n1099), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1095), .A2(KEYINPUT61), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT61), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1098), .A2(new_n1107), .A3(new_n1088), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n1101), .A2(new_n618), .A3(new_n1103), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT60), .B1(new_n1110), .B2(new_n1104), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT58), .B(G1341), .ZN(new_n1112));
  OAI22_X1  g687(.A1(new_n1015), .A2(G1996), .B1(new_n1003), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n571), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1113), .A2(KEYINPUT59), .A3(new_n571), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT60), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1101), .A2(new_n1118), .A3(new_n619), .A4(new_n1103), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1111), .A2(new_n1116), .A3(new_n1117), .A4(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1105), .B1(new_n1109), .B2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1042), .A2(new_n1071), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n1082), .B2(G171), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n977), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n476), .B1(new_n1126), .B2(new_n1013), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n1128));
  OAI21_X1  g703(.A(G2105), .B1(new_n485), .B2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n489), .A2(KEYINPUT122), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1131), .A2(new_n989), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1127), .A2(new_n1012), .A3(new_n1080), .A4(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1079), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1125), .B1(new_n1134), .B2(G171), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1079), .A2(KEYINPUT123), .A3(G301), .A4(new_n1081), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1124), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1079), .A2(G301), .A3(new_n1133), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1083), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1084), .B1(new_n1139), .B2(new_n1125), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1121), .A2(new_n1122), .A3(new_n1137), .A4(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1007), .B1(new_n1006), .B2(new_n974), .ZN(new_n1142));
  AOI211_X1 g717(.A(KEYINPUT119), .B(new_n973), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1031), .B(new_n1033), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1058), .A2(G286), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT63), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1147), .B1(new_n1023), .B2(new_n1026), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1145), .A2(new_n1041), .A3(new_n1146), .A4(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1146), .ZN(new_n1150));
  NOR4_X1   g725(.A1(new_n1144), .A2(new_n1071), .A3(new_n1027), .A4(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1149), .B1(new_n1151), .B2(KEYINPUT63), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1087), .A2(new_n1141), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(G1384), .B1(new_n872), .B2(new_n874), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1154), .A2(new_n1002), .A3(KEYINPUT45), .ZN(new_n1155));
  INV_X1    g730(.A(G1986), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n607), .A2(new_n1156), .ZN(new_n1157));
  XOR2_X1   g732(.A(new_n1157), .B(KEYINPUT111), .Z(new_n1158));
  NOR2_X1   g733(.A1(new_n607), .A2(new_n1156), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1155), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT113), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n783), .A2(G2067), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n780), .A2(new_n781), .A3(new_n782), .A4(new_n1102), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1155), .A2(new_n1161), .A3(new_n1164), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n990), .A2(new_n1126), .A3(new_n1164), .A4(new_n1013), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(KEYINPUT113), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  NOR4_X1   g743(.A1(new_n735), .A2(new_n1154), .A3(new_n1002), .A4(KEYINPUT45), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(G1996), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(G1996), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1155), .A2(KEYINPUT112), .A3(new_n1172), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n990), .A2(new_n1126), .A3(new_n1013), .A4(new_n1172), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT112), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n734), .B1(new_n1173), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(KEYINPUT114), .B1(new_n1171), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(KEYINPUT112), .B1(new_n1155), .B2(new_n1172), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n735), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT114), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1181), .A2(new_n1182), .A3(new_n1170), .A4(new_n1168), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n820), .A2(new_n824), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n819), .A2(new_n823), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1155), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  AND4_X1   g761(.A1(new_n1160), .A2(new_n1178), .A3(new_n1183), .A4(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1153), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1178), .A2(new_n1183), .A3(new_n1185), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1189), .A2(new_n1163), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1190), .A2(new_n1155), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1158), .A2(new_n1155), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n1192), .B(KEYINPUT125), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n1193), .B(KEYINPUT48), .ZN(new_n1194));
  NAND4_X1  g769(.A1(new_n1194), .A2(new_n1178), .A3(new_n1183), .A4(new_n1186), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT46), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1196), .A2(KEYINPUT124), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1197), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1166), .B1(KEYINPUT124), .B2(new_n1196), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1199), .A2(new_n1169), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1173), .A2(new_n1176), .A3(KEYINPUT124), .A4(new_n1196), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1198), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1202), .B(KEYINPUT47), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1191), .A2(new_n1195), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1204), .A2(KEYINPUT126), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT126), .ZN(new_n1206));
  NAND4_X1  g781(.A1(new_n1191), .A2(new_n1195), .A3(new_n1203), .A4(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1188), .A2(new_n1208), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g784(.A1(G227), .A2(new_n462), .ZN(new_n1211));
  NAND3_X1  g785(.A1(new_n702), .A2(new_n1211), .A3(new_n664), .ZN(new_n1212));
  OR2_X1    g786(.A1(new_n1212), .A2(KEYINPUT127), .ZN(new_n1213));
  NAND2_X1  g787(.A1(new_n1212), .A2(KEYINPUT127), .ZN(new_n1214));
  NAND4_X1  g788(.A1(new_n1213), .A2(new_n962), .A3(new_n909), .A4(new_n1214), .ZN(G225));
  INV_X1    g789(.A(G225), .ZN(G308));
endmodule


