

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U555 ( .A1(G2104), .A2(n548), .ZN(n897) );
  XOR2_X1 U556 ( .A(KEYINPUT69), .B(n611), .Z(n521) );
  INV_X1 U557 ( .A(KEYINPUT96), .ZN(n656) );
  BUF_X1 U558 ( .A(n650), .Z(n668) );
  INV_X1 U559 ( .A(KEYINPUT99), .ZN(n666) );
  XNOR2_X1 U560 ( .A(n667), .B(n666), .ZN(n673) );
  AND2_X1 U561 ( .A1(n590), .A2(G40), .ZN(n591) );
  NAND2_X1 U562 ( .A1(n694), .A2(n696), .ZN(n650) );
  NOR2_X1 U563 ( .A1(G2105), .A2(G2104), .ZN(n544) );
  XNOR2_X1 U564 ( .A(n522), .B(KEYINPUT65), .ZN(n538) );
  NOR2_X2 U565 ( .A1(G651), .A2(n538), .ZN(n817) );
  NOR2_X2 U566 ( .A1(n538), .A2(n529), .ZN(n813) );
  AND2_X2 U567 ( .A1(n548), .A2(G2104), .ZN(n900) );
  XOR2_X1 U568 ( .A(KEYINPUT15), .B(n633), .Z(n935) );
  XOR2_X1 U569 ( .A(KEYINPUT1), .B(n524), .Z(n820) );
  NOR2_X1 U570 ( .A1(n588), .A2(n587), .ZN(n782) );
  XNOR2_X1 U571 ( .A(G543), .B(KEYINPUT0), .ZN(n522) );
  NAND2_X1 U572 ( .A1(n817), .A2(G51), .ZN(n523) );
  XNOR2_X1 U573 ( .A(n523), .B(KEYINPUT74), .ZN(n526) );
  INV_X1 U574 ( .A(G651), .ZN(n529) );
  NOR2_X1 U575 ( .A1(G543), .A2(n529), .ZN(n524) );
  NAND2_X1 U576 ( .A1(G63), .A2(n820), .ZN(n525) );
  NAND2_X1 U577 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U578 ( .A(KEYINPUT6), .B(n527), .ZN(n535) );
  NOR2_X1 U579 ( .A1(G651), .A2(G543), .ZN(n811) );
  NAND2_X1 U580 ( .A1(n811), .A2(G89), .ZN(n528) );
  XNOR2_X1 U581 ( .A(n528), .B(KEYINPUT4), .ZN(n531) );
  NAND2_X1 U582 ( .A1(G76), .A2(n813), .ZN(n530) );
  NAND2_X1 U583 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U584 ( .A(KEYINPUT5), .B(n532), .ZN(n533) );
  XNOR2_X1 U585 ( .A(KEYINPUT73), .B(n533), .ZN(n534) );
  NOR2_X1 U586 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U587 ( .A(KEYINPUT7), .B(n536), .Z(G168) );
  XNOR2_X1 U588 ( .A(G168), .B(KEYINPUT8), .ZN(n537) );
  XNOR2_X1 U589 ( .A(n537), .B(KEYINPUT75), .ZN(G286) );
  NAND2_X1 U590 ( .A1(G49), .A2(n817), .ZN(n540) );
  NAND2_X1 U591 ( .A1(G87), .A2(n538), .ZN(n539) );
  NAND2_X1 U592 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U593 ( .A1(n820), .A2(n541), .ZN(n543) );
  NAND2_X1 U594 ( .A1(G651), .A2(G74), .ZN(n542) );
  NAND2_X1 U595 ( .A1(n543), .A2(n542), .ZN(G288) );
  INV_X1 U596 ( .A(G2105), .ZN(n548) );
  NAND2_X1 U597 ( .A1(G102), .A2(n900), .ZN(n547) );
  XOR2_X1 U598 ( .A(KEYINPUT17), .B(n544), .Z(n545) );
  XNOR2_X1 U599 ( .A(n545), .B(KEYINPUT64), .ZN(n697) );
  NAND2_X1 U600 ( .A1(G138), .A2(n697), .ZN(n546) );
  NAND2_X1 U601 ( .A1(n547), .A2(n546), .ZN(n552) );
  AND2_X1 U602 ( .A1(G2105), .A2(G2104), .ZN(n896) );
  NAND2_X1 U603 ( .A1(G114), .A2(n896), .ZN(n550) );
  NAND2_X1 U604 ( .A1(G126), .A2(n897), .ZN(n549) );
  NAND2_X1 U605 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U606 ( .A1(n552), .A2(n551), .ZN(G164) );
  NAND2_X1 U607 ( .A1(G52), .A2(n817), .ZN(n554) );
  NAND2_X1 U608 ( .A1(G64), .A2(n820), .ZN(n553) );
  NAND2_X1 U609 ( .A1(n554), .A2(n553), .ZN(n559) );
  NAND2_X1 U610 ( .A1(G90), .A2(n811), .ZN(n556) );
  NAND2_X1 U611 ( .A1(G77), .A2(n813), .ZN(n555) );
  NAND2_X1 U612 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U613 ( .A(KEYINPUT9), .B(n557), .Z(n558) );
  NOR2_X1 U614 ( .A1(n559), .A2(n558), .ZN(G171) );
  NAND2_X1 U615 ( .A1(n820), .A2(G62), .ZN(n561) );
  NAND2_X1 U616 ( .A1(n817), .A2(G50), .ZN(n560) );
  NAND2_X1 U617 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U618 ( .A(KEYINPUT84), .B(n562), .ZN(n566) );
  NAND2_X1 U619 ( .A1(G88), .A2(n811), .ZN(n564) );
  NAND2_X1 U620 ( .A1(G75), .A2(n813), .ZN(n563) );
  NAND2_X1 U621 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U622 ( .A1(n566), .A2(n565), .ZN(G166) );
  INV_X1 U623 ( .A(G166), .ZN(G303) );
  NAND2_X1 U624 ( .A1(G48), .A2(n817), .ZN(n568) );
  NAND2_X1 U625 ( .A1(G86), .A2(n811), .ZN(n567) );
  NAND2_X1 U626 ( .A1(n568), .A2(n567), .ZN(n571) );
  NAND2_X1 U627 ( .A1(n813), .A2(G73), .ZN(n569) );
  XOR2_X1 U628 ( .A(KEYINPUT2), .B(n569), .Z(n570) );
  NOR2_X1 U629 ( .A1(n571), .A2(n570), .ZN(n573) );
  NAND2_X1 U630 ( .A1(n820), .A2(G61), .ZN(n572) );
  NAND2_X1 U631 ( .A1(n573), .A2(n572), .ZN(G305) );
  NAND2_X1 U632 ( .A1(G85), .A2(n811), .ZN(n575) );
  NAND2_X1 U633 ( .A1(G72), .A2(n813), .ZN(n574) );
  NAND2_X1 U634 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U635 ( .A(KEYINPUT66), .B(n576), .ZN(n579) );
  NAND2_X1 U636 ( .A1(G47), .A2(n817), .ZN(n577) );
  XNOR2_X1 U637 ( .A(KEYINPUT67), .B(n577), .ZN(n578) );
  NOR2_X1 U638 ( .A1(n579), .A2(n578), .ZN(n581) );
  NAND2_X1 U639 ( .A1(n820), .A2(G60), .ZN(n580) );
  NAND2_X1 U640 ( .A1(n581), .A2(n580), .ZN(G290) );
  NOR2_X1 U641 ( .A1(G1976), .A2(G288), .ZN(n942) );
  NAND2_X1 U642 ( .A1(n896), .A2(G113), .ZN(n584) );
  NAND2_X1 U643 ( .A1(G101), .A2(n900), .ZN(n582) );
  XOR2_X1 U644 ( .A(KEYINPUT23), .B(n582), .Z(n583) );
  NAND2_X1 U645 ( .A1(n584), .A2(n583), .ZN(n588) );
  NAND2_X1 U646 ( .A1(n697), .A2(G137), .ZN(n586) );
  NAND2_X1 U647 ( .A1(n897), .A2(G125), .ZN(n585) );
  NAND2_X1 U648 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U649 ( .A1(n782), .A2(G40), .ZN(n589) );
  NAND2_X1 U650 ( .A1(n589), .A2(KEYINPUT87), .ZN(n593) );
  INV_X1 U651 ( .A(KEYINPUT87), .ZN(n590) );
  NAND2_X1 U652 ( .A1(n782), .A2(n591), .ZN(n592) );
  NAND2_X1 U653 ( .A1(n593), .A2(n592), .ZN(n694) );
  NOR2_X1 U654 ( .A1(G164), .A2(G1384), .ZN(n696) );
  NAND2_X1 U655 ( .A1(n668), .A2(G1961), .ZN(n595) );
  INV_X1 U656 ( .A(n668), .ZN(n634) );
  XOR2_X1 U657 ( .A(G2078), .B(KEYINPUT25), .Z(n1019) );
  NAND2_X1 U658 ( .A1(n634), .A2(n1019), .ZN(n594) );
  NAND2_X1 U659 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U660 ( .A(n596), .B(KEYINPUT92), .Z(n658) );
  NAND2_X1 U661 ( .A1(n658), .A2(G171), .ZN(n649) );
  NAND2_X1 U662 ( .A1(G53), .A2(n817), .ZN(n598) );
  NAND2_X1 U663 ( .A1(G65), .A2(n820), .ZN(n597) );
  NAND2_X1 U664 ( .A1(n598), .A2(n597), .ZN(n602) );
  NAND2_X1 U665 ( .A1(G91), .A2(n811), .ZN(n600) );
  NAND2_X1 U666 ( .A1(G78), .A2(n813), .ZN(n599) );
  NAND2_X1 U667 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U668 ( .A1(n602), .A2(n601), .ZN(n939) );
  NAND2_X1 U669 ( .A1(n634), .A2(G2072), .ZN(n603) );
  XNOR2_X1 U670 ( .A(n603), .B(KEYINPUT27), .ZN(n605) );
  AND2_X1 U671 ( .A1(G1956), .A2(n668), .ZN(n604) );
  NOR2_X1 U672 ( .A1(n605), .A2(n604), .ZN(n608) );
  NOR2_X1 U673 ( .A1(n939), .A2(n608), .ZN(n607) );
  XNOR2_X1 U674 ( .A(KEYINPUT28), .B(KEYINPUT93), .ZN(n606) );
  XNOR2_X1 U675 ( .A(n607), .B(n606), .ZN(n646) );
  NAND2_X1 U676 ( .A1(n939), .A2(n608), .ZN(n644) );
  NAND2_X1 U677 ( .A1(G81), .A2(n811), .ZN(n609) );
  XNOR2_X1 U678 ( .A(n609), .B(KEYINPUT68), .ZN(n610) );
  XNOR2_X1 U679 ( .A(KEYINPUT12), .B(n610), .ZN(n612) );
  NAND2_X1 U680 ( .A1(n813), .A2(G68), .ZN(n611) );
  NAND2_X1 U681 ( .A1(n612), .A2(n521), .ZN(n613) );
  XNOR2_X1 U682 ( .A(n613), .B(KEYINPUT13), .ZN(n615) );
  NAND2_X1 U683 ( .A1(G43), .A2(n817), .ZN(n614) );
  NAND2_X1 U684 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U685 ( .A1(n820), .A2(G56), .ZN(n616) );
  XOR2_X1 U686 ( .A(KEYINPUT14), .B(n616), .Z(n617) );
  NOR2_X1 U687 ( .A1(n618), .A2(n617), .ZN(n619) );
  XOR2_X2 U688 ( .A(KEYINPUT70), .B(n619), .Z(n951) );
  INV_X1 U689 ( .A(G1996), .ZN(n879) );
  NOR2_X1 U690 ( .A1(n650), .A2(n879), .ZN(n621) );
  XOR2_X1 U691 ( .A(KEYINPUT26), .B(KEYINPUT94), .Z(n620) );
  XNOR2_X1 U692 ( .A(n621), .B(n620), .ZN(n623) );
  NAND2_X1 U693 ( .A1(n668), .A2(G1341), .ZN(n622) );
  NAND2_X1 U694 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U695 ( .A(n624), .B(KEYINPUT95), .ZN(n638) );
  NAND2_X1 U696 ( .A1(n820), .A2(G66), .ZN(n632) );
  NAND2_X1 U697 ( .A1(G54), .A2(n817), .ZN(n626) );
  NAND2_X1 U698 ( .A1(G79), .A2(n813), .ZN(n625) );
  NAND2_X1 U699 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U700 ( .A(KEYINPUT72), .B(n627), .ZN(n630) );
  NAND2_X1 U701 ( .A1(G92), .A2(n811), .ZN(n628) );
  XNOR2_X1 U702 ( .A(KEYINPUT71), .B(n628), .ZN(n629) );
  NOR2_X1 U703 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U704 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U705 ( .A1(G1348), .A2(n668), .ZN(n636) );
  NAND2_X1 U706 ( .A1(n634), .A2(G2067), .ZN(n635) );
  NAND2_X1 U707 ( .A1(n636), .A2(n635), .ZN(n640) );
  NAND2_X1 U708 ( .A1(n935), .A2(n640), .ZN(n637) );
  NAND2_X1 U709 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U710 ( .A1(n951), .A2(n639), .ZN(n642) );
  NOR2_X1 U711 ( .A1(n640), .A2(n935), .ZN(n641) );
  NOR2_X1 U712 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U713 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U714 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U715 ( .A(KEYINPUT29), .B(n647), .Z(n648) );
  NAND2_X1 U716 ( .A1(n649), .A2(n648), .ZN(n665) );
  NAND2_X1 U717 ( .A1(G8), .A2(n650), .ZN(n746) );
  NOR2_X1 U718 ( .A1(G1966), .A2(n746), .ZN(n681) );
  NOR2_X1 U719 ( .A1(G2084), .A2(n650), .ZN(n651) );
  INV_X1 U720 ( .A(n651), .ZN(n677) );
  NAND2_X1 U721 ( .A1(G8), .A2(n677), .ZN(n652) );
  NOR2_X1 U722 ( .A1(n681), .A2(n652), .ZN(n654) );
  INV_X1 U723 ( .A(KEYINPUT30), .ZN(n653) );
  XNOR2_X1 U724 ( .A(n654), .B(n653), .ZN(n655) );
  NOR2_X1 U725 ( .A1(G168), .A2(n655), .ZN(n657) );
  XNOR2_X1 U726 ( .A(n657), .B(n656), .ZN(n660) );
  OR2_X1 U727 ( .A1(G171), .A2(n658), .ZN(n659) );
  NAND2_X1 U728 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U729 ( .A(n661), .B(KEYINPUT31), .ZN(n663) );
  INV_X1 U730 ( .A(KEYINPUT97), .ZN(n662) );
  XNOR2_X1 U731 ( .A(n663), .B(n662), .ZN(n664) );
  NAND2_X1 U732 ( .A1(n665), .A2(n664), .ZN(n676) );
  NAND2_X1 U733 ( .A1(n676), .A2(G286), .ZN(n667) );
  NOR2_X1 U734 ( .A1(G1971), .A2(n746), .ZN(n670) );
  NOR2_X1 U735 ( .A1(G2090), .A2(n668), .ZN(n669) );
  NOR2_X1 U736 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U737 ( .A1(G303), .A2(n671), .ZN(n672) );
  NAND2_X1 U738 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U739 ( .A1(n674), .A2(G8), .ZN(n675) );
  XOR2_X1 U740 ( .A(n675), .B(KEYINPUT32), .Z(n683) );
  XNOR2_X1 U741 ( .A(n676), .B(KEYINPUT98), .ZN(n679) );
  NAND2_X1 U742 ( .A1(n651), .A2(G8), .ZN(n678) );
  NAND2_X1 U743 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U744 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U745 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U746 ( .A(KEYINPUT100), .B(n684), .ZN(n739) );
  NOR2_X1 U747 ( .A1(n942), .A2(n739), .ZN(n687) );
  NOR2_X1 U748 ( .A1(G1971), .A2(G303), .ZN(n685) );
  XNOR2_X1 U749 ( .A(n685), .B(KEYINPUT101), .ZN(n686) );
  NAND2_X1 U750 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U751 ( .A1(G1976), .A2(G288), .ZN(n943) );
  NAND2_X1 U752 ( .A1(n688), .A2(n943), .ZN(n689) );
  XNOR2_X1 U753 ( .A(n689), .B(KEYINPUT102), .ZN(n731) );
  NAND2_X1 U754 ( .A1(n942), .A2(KEYINPUT33), .ZN(n690) );
  NOR2_X1 U755 ( .A1(n690), .A2(n746), .ZN(n693) );
  XNOR2_X1 U756 ( .A(G1981), .B(KEYINPUT103), .ZN(n691) );
  XNOR2_X1 U757 ( .A(n691), .B(G305), .ZN(n932) );
  INV_X1 U758 ( .A(n932), .ZN(n692) );
  NOR2_X1 U759 ( .A1(n693), .A2(n692), .ZN(n710) );
  INV_X1 U760 ( .A(n694), .ZN(n695) );
  NOR2_X1 U761 ( .A1(n696), .A2(n695), .ZN(n765) );
  XNOR2_X1 U762 ( .A(G2067), .B(KEYINPUT37), .ZN(n762) );
  INV_X1 U763 ( .A(n697), .ZN(n698) );
  INV_X1 U764 ( .A(n698), .ZN(n902) );
  NAND2_X1 U765 ( .A1(G140), .A2(n902), .ZN(n699) );
  XNOR2_X1 U766 ( .A(n699), .B(KEYINPUT88), .ZN(n701) );
  NAND2_X1 U767 ( .A1(G104), .A2(n900), .ZN(n700) );
  NAND2_X1 U768 ( .A1(n701), .A2(n700), .ZN(n703) );
  XOR2_X1 U769 ( .A(KEYINPUT89), .B(KEYINPUT34), .Z(n702) );
  XNOR2_X1 U770 ( .A(n703), .B(n702), .ZN(n708) );
  NAND2_X1 U771 ( .A1(G116), .A2(n896), .ZN(n705) );
  NAND2_X1 U772 ( .A1(G128), .A2(n897), .ZN(n704) );
  NAND2_X1 U773 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U774 ( .A(KEYINPUT35), .B(n706), .Z(n707) );
  NOR2_X1 U775 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U776 ( .A(KEYINPUT36), .B(n709), .ZN(n921) );
  NOR2_X1 U777 ( .A1(n762), .A2(n921), .ZN(n1009) );
  NAND2_X1 U778 ( .A1(n765), .A2(n1009), .ZN(n760) );
  AND2_X1 U779 ( .A1(n710), .A2(n760), .ZN(n729) );
  XOR2_X1 U780 ( .A(G1986), .B(G290), .Z(n945) );
  NAND2_X1 U781 ( .A1(G95), .A2(n900), .ZN(n712) );
  NAND2_X1 U782 ( .A1(G131), .A2(n902), .ZN(n711) );
  NAND2_X1 U783 ( .A1(n712), .A2(n711), .ZN(n716) );
  NAND2_X1 U784 ( .A1(G107), .A2(n896), .ZN(n714) );
  NAND2_X1 U785 ( .A1(G119), .A2(n897), .ZN(n713) );
  NAND2_X1 U786 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U787 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U788 ( .A(n717), .B(KEYINPUT90), .Z(n916) );
  AND2_X1 U789 ( .A1(G1991), .A2(n916), .ZN(n727) );
  NAND2_X1 U790 ( .A1(G105), .A2(n900), .ZN(n718) );
  XNOR2_X1 U791 ( .A(n718), .B(KEYINPUT38), .ZN(n721) );
  NAND2_X1 U792 ( .A1(G117), .A2(n896), .ZN(n719) );
  XOR2_X1 U793 ( .A(KEYINPUT91), .B(n719), .Z(n720) );
  NAND2_X1 U794 ( .A1(n721), .A2(n720), .ZN(n725) );
  NAND2_X1 U795 ( .A1(n897), .A2(G129), .ZN(n723) );
  NAND2_X1 U796 ( .A1(G141), .A2(n902), .ZN(n722) );
  NAND2_X1 U797 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U798 ( .A1(n725), .A2(n724), .ZN(n909) );
  NOR2_X1 U799 ( .A1(n909), .A2(n879), .ZN(n726) );
  NOR2_X1 U800 ( .A1(n727), .A2(n726), .ZN(n999) );
  NAND2_X1 U801 ( .A1(n945), .A2(n999), .ZN(n728) );
  NAND2_X1 U802 ( .A1(n728), .A2(n765), .ZN(n736) );
  NAND2_X1 U803 ( .A1(n729), .A2(n736), .ZN(n732) );
  OR2_X1 U804 ( .A1(n746), .A2(n732), .ZN(n730) );
  NOR2_X1 U805 ( .A1(n731), .A2(n730), .ZN(n735) );
  INV_X1 U806 ( .A(n732), .ZN(n733) );
  AND2_X1 U807 ( .A1(n733), .A2(KEYINPUT33), .ZN(n734) );
  NOR2_X1 U808 ( .A1(n735), .A2(n734), .ZN(n770) );
  INV_X1 U809 ( .A(n736), .ZN(n751) );
  NOR2_X1 U810 ( .A1(G2090), .A2(G303), .ZN(n737) );
  XNOR2_X1 U811 ( .A(KEYINPUT104), .B(n737), .ZN(n738) );
  NAND2_X1 U812 ( .A1(n738), .A2(G8), .ZN(n741) );
  INV_X1 U813 ( .A(n739), .ZN(n740) );
  NAND2_X1 U814 ( .A1(n741), .A2(n740), .ZN(n743) );
  AND2_X1 U815 ( .A1(n746), .A2(n760), .ZN(n742) );
  AND2_X1 U816 ( .A1(n743), .A2(n742), .ZN(n749) );
  NOR2_X1 U817 ( .A1(G1981), .A2(G305), .ZN(n744) );
  XOR2_X1 U818 ( .A(n744), .B(KEYINPUT24), .Z(n745) );
  NOR2_X1 U819 ( .A1(n746), .A2(n745), .ZN(n747) );
  AND2_X1 U820 ( .A1(n760), .A2(n747), .ZN(n748) );
  NOR2_X1 U821 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U822 ( .A1(n751), .A2(n750), .ZN(n768) );
  AND2_X1 U823 ( .A1(n879), .A2(n909), .ZN(n989) );
  INV_X1 U824 ( .A(n999), .ZN(n756) );
  NOR2_X1 U825 ( .A1(G1986), .A2(G290), .ZN(n753) );
  NOR2_X1 U826 ( .A1(G1991), .A2(n916), .ZN(n752) );
  XOR2_X1 U827 ( .A(KEYINPUT105), .B(n752), .Z(n992) );
  NOR2_X1 U828 ( .A1(n753), .A2(n992), .ZN(n754) );
  XNOR2_X1 U829 ( .A(n754), .B(KEYINPUT106), .ZN(n755) );
  NOR2_X1 U830 ( .A1(n756), .A2(n755), .ZN(n757) );
  NOR2_X1 U831 ( .A1(n989), .A2(n757), .ZN(n758) );
  XOR2_X1 U832 ( .A(KEYINPUT39), .B(n758), .Z(n759) );
  XNOR2_X1 U833 ( .A(n759), .B(KEYINPUT107), .ZN(n761) );
  NAND2_X1 U834 ( .A1(n761), .A2(n760), .ZN(n763) );
  NAND2_X1 U835 ( .A1(n762), .A2(n921), .ZN(n1006) );
  NAND2_X1 U836 ( .A1(n763), .A2(n1006), .ZN(n764) );
  XNOR2_X1 U837 ( .A(KEYINPUT108), .B(n764), .ZN(n766) );
  AND2_X1 U838 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U839 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U840 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U841 ( .A(n771), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U842 ( .A(G2446), .B(G2451), .Z(n773) );
  XNOR2_X1 U843 ( .A(G2454), .B(KEYINPUT109), .ZN(n772) );
  XNOR2_X1 U844 ( .A(n773), .B(n772), .ZN(n780) );
  XOR2_X1 U845 ( .A(G2438), .B(G2430), .Z(n775) );
  XNOR2_X1 U846 ( .A(G2435), .B(G2443), .ZN(n774) );
  XNOR2_X1 U847 ( .A(n775), .B(n774), .ZN(n776) );
  XOR2_X1 U848 ( .A(n776), .B(G2427), .Z(n778) );
  XNOR2_X1 U849 ( .A(G1348), .B(G1341), .ZN(n777) );
  XNOR2_X1 U850 ( .A(n778), .B(n777), .ZN(n779) );
  XNOR2_X1 U851 ( .A(n780), .B(n779), .ZN(n781) );
  AND2_X1 U852 ( .A1(n781), .A2(G14), .ZN(G401) );
  AND2_X1 U853 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U854 ( .A(G860), .ZN(n790) );
  OR2_X1 U855 ( .A1(n790), .A2(n951), .ZN(G153) );
  INV_X1 U856 ( .A(G132), .ZN(G219) );
  INV_X1 U857 ( .A(G82), .ZN(G220) );
  INV_X1 U858 ( .A(G57), .ZN(G237) );
  INV_X1 U859 ( .A(G108), .ZN(G238) );
  INV_X1 U860 ( .A(G120), .ZN(G236) );
  BUF_X1 U861 ( .A(n782), .Z(G160) );
  INV_X1 U862 ( .A(G171), .ZN(G301) );
  NAND2_X1 U863 ( .A1(G7), .A2(G661), .ZN(n783) );
  XNOR2_X1 U864 ( .A(n783), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U865 ( .A(G223), .ZN(n850) );
  NAND2_X1 U866 ( .A1(n850), .A2(G567), .ZN(n784) );
  XOR2_X1 U867 ( .A(KEYINPUT11), .B(n784), .Z(G234) );
  NAND2_X1 U868 ( .A1(G868), .A2(G301), .ZN(n786) );
  INV_X1 U869 ( .A(G868), .ZN(n832) );
  NAND2_X1 U870 ( .A1(n935), .A2(n832), .ZN(n785) );
  NAND2_X1 U871 ( .A1(n786), .A2(n785), .ZN(G284) );
  INV_X1 U872 ( .A(n939), .ZN(G299) );
  NOR2_X1 U873 ( .A1(G868), .A2(G299), .ZN(n787) );
  XNOR2_X1 U874 ( .A(n787), .B(KEYINPUT76), .ZN(n789) );
  NOR2_X1 U875 ( .A1(n832), .A2(G286), .ZN(n788) );
  NOR2_X1 U876 ( .A1(n789), .A2(n788), .ZN(G297) );
  NAND2_X1 U877 ( .A1(n790), .A2(G559), .ZN(n791) );
  INV_X1 U878 ( .A(n935), .ZN(n809) );
  NAND2_X1 U879 ( .A1(n791), .A2(n809), .ZN(n792) );
  XNOR2_X1 U880 ( .A(n792), .B(KEYINPUT77), .ZN(n793) );
  XOR2_X1 U881 ( .A(KEYINPUT16), .B(n793), .Z(G148) );
  NOR2_X1 U882 ( .A1(n935), .A2(n832), .ZN(n794) );
  XOR2_X1 U883 ( .A(KEYINPUT78), .B(n794), .Z(n795) );
  NOR2_X1 U884 ( .A1(G559), .A2(n795), .ZN(n796) );
  XOR2_X1 U885 ( .A(KEYINPUT79), .B(n796), .Z(n798) );
  NOR2_X1 U886 ( .A1(n951), .A2(G868), .ZN(n797) );
  NOR2_X1 U887 ( .A1(n798), .A2(n797), .ZN(G282) );
  NAND2_X1 U888 ( .A1(G123), .A2(n897), .ZN(n799) );
  XNOR2_X1 U889 ( .A(n799), .B(KEYINPUT18), .ZN(n802) );
  NAND2_X1 U890 ( .A1(G111), .A2(n896), .ZN(n800) );
  XNOR2_X1 U891 ( .A(n800), .B(KEYINPUT80), .ZN(n801) );
  NAND2_X1 U892 ( .A1(n802), .A2(n801), .ZN(n806) );
  NAND2_X1 U893 ( .A1(G99), .A2(n900), .ZN(n804) );
  NAND2_X1 U894 ( .A1(G135), .A2(n902), .ZN(n803) );
  NAND2_X1 U895 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U896 ( .A1(n806), .A2(n805), .ZN(n991) );
  XNOR2_X1 U897 ( .A(n991), .B(G2096), .ZN(n808) );
  INV_X1 U898 ( .A(G2100), .ZN(n807) );
  NAND2_X1 U899 ( .A1(n808), .A2(n807), .ZN(G156) );
  NAND2_X1 U900 ( .A1(G559), .A2(n809), .ZN(n810) );
  XNOR2_X1 U901 ( .A(n810), .B(n951), .ZN(n830) );
  NOR2_X1 U902 ( .A1(G860), .A2(n830), .ZN(n824) );
  NAND2_X1 U903 ( .A1(G93), .A2(n811), .ZN(n812) );
  XNOR2_X1 U904 ( .A(n812), .B(KEYINPUT81), .ZN(n816) );
  NAND2_X1 U905 ( .A1(G80), .A2(n813), .ZN(n814) );
  XOR2_X1 U906 ( .A(KEYINPUT82), .B(n814), .Z(n815) );
  NOR2_X1 U907 ( .A1(n816), .A2(n815), .ZN(n819) );
  NAND2_X1 U908 ( .A1(n817), .A2(G55), .ZN(n818) );
  NAND2_X1 U909 ( .A1(n819), .A2(n818), .ZN(n823) );
  NAND2_X1 U910 ( .A1(G67), .A2(n820), .ZN(n821) );
  XNOR2_X1 U911 ( .A(KEYINPUT83), .B(n821), .ZN(n822) );
  OR2_X1 U912 ( .A1(n823), .A2(n822), .ZN(n833) );
  XOR2_X1 U913 ( .A(n824), .B(n833), .Z(G145) );
  XNOR2_X1 U914 ( .A(KEYINPUT19), .B(n833), .ZN(n825) );
  XNOR2_X1 U915 ( .A(G288), .B(n825), .ZN(n826) );
  XNOR2_X1 U916 ( .A(G305), .B(n826), .ZN(n828) );
  XNOR2_X1 U917 ( .A(G166), .B(n939), .ZN(n827) );
  XNOR2_X1 U918 ( .A(n828), .B(n827), .ZN(n829) );
  XNOR2_X1 U919 ( .A(n829), .B(G290), .ZN(n858) );
  XOR2_X1 U920 ( .A(n858), .B(n830), .Z(n831) );
  NOR2_X1 U921 ( .A1(n832), .A2(n831), .ZN(n835) );
  NOR2_X1 U922 ( .A1(G868), .A2(n833), .ZN(n834) );
  NOR2_X1 U923 ( .A1(n835), .A2(n834), .ZN(G295) );
  NAND2_X1 U924 ( .A1(G2084), .A2(G2078), .ZN(n836) );
  XOR2_X1 U925 ( .A(KEYINPUT20), .B(n836), .Z(n837) );
  NAND2_X1 U926 ( .A1(G2090), .A2(n837), .ZN(n838) );
  XNOR2_X1 U927 ( .A(KEYINPUT21), .B(n838), .ZN(n839) );
  NAND2_X1 U928 ( .A1(n839), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U929 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U930 ( .A1(G236), .A2(G238), .ZN(n840) );
  NAND2_X1 U931 ( .A1(G69), .A2(n840), .ZN(n841) );
  NOR2_X1 U932 ( .A1(n841), .A2(G237), .ZN(n842) );
  XNOR2_X1 U933 ( .A(n842), .B(KEYINPUT85), .ZN(n855) );
  NAND2_X1 U934 ( .A1(n855), .A2(G567), .ZN(n847) );
  NOR2_X1 U935 ( .A1(G220), .A2(G219), .ZN(n843) );
  XOR2_X1 U936 ( .A(KEYINPUT22), .B(n843), .Z(n844) );
  NOR2_X1 U937 ( .A1(G218), .A2(n844), .ZN(n845) );
  NAND2_X1 U938 ( .A1(G96), .A2(n845), .ZN(n854) );
  NAND2_X1 U939 ( .A1(n854), .A2(G2106), .ZN(n846) );
  NAND2_X1 U940 ( .A1(n847), .A2(n846), .ZN(n931) );
  NAND2_X1 U941 ( .A1(G661), .A2(G483), .ZN(n848) );
  XNOR2_X1 U942 ( .A(KEYINPUT86), .B(n848), .ZN(n849) );
  NOR2_X1 U943 ( .A1(n931), .A2(n849), .ZN(n853) );
  NAND2_X1 U944 ( .A1(n853), .A2(G36), .ZN(G176) );
  NAND2_X1 U945 ( .A1(G2106), .A2(n850), .ZN(G217) );
  AND2_X1 U946 ( .A1(G15), .A2(G2), .ZN(n851) );
  NAND2_X1 U947 ( .A1(G661), .A2(n851), .ZN(G259) );
  NAND2_X1 U948 ( .A1(G3), .A2(G1), .ZN(n852) );
  NAND2_X1 U949 ( .A1(n853), .A2(n852), .ZN(G188) );
  INV_X1 U951 ( .A(G96), .ZN(G221) );
  NOR2_X1 U952 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U953 ( .A(n856), .B(KEYINPUT110), .ZN(G325) );
  INV_X1 U954 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U955 ( .A(G286), .B(G301), .ZN(n857) );
  XNOR2_X1 U956 ( .A(n857), .B(n935), .ZN(n860) );
  XNOR2_X1 U957 ( .A(n951), .B(n858), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n860), .B(n859), .ZN(n861) );
  NOR2_X1 U959 ( .A1(G37), .A2(n861), .ZN(G397) );
  XOR2_X1 U960 ( .A(G2100), .B(G2096), .Z(n863) );
  XNOR2_X1 U961 ( .A(KEYINPUT42), .B(G2678), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n863), .B(n862), .ZN(n867) );
  XOR2_X1 U963 ( .A(KEYINPUT43), .B(G2072), .Z(n865) );
  XNOR2_X1 U964 ( .A(G2090), .B(G2067), .ZN(n864) );
  XNOR2_X1 U965 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U966 ( .A(n867), .B(n866), .Z(n869) );
  XNOR2_X1 U967 ( .A(G2084), .B(G2078), .ZN(n868) );
  XNOR2_X1 U968 ( .A(n869), .B(n868), .ZN(G227) );
  XOR2_X1 U969 ( .A(G1991), .B(G1986), .Z(n871) );
  XNOR2_X1 U970 ( .A(G1961), .B(G1971), .ZN(n870) );
  XNOR2_X1 U971 ( .A(n871), .B(n870), .ZN(n875) );
  XOR2_X1 U972 ( .A(G1976), .B(G1981), .Z(n873) );
  XNOR2_X1 U973 ( .A(G1966), .B(G1956), .ZN(n872) );
  XNOR2_X1 U974 ( .A(n873), .B(n872), .ZN(n874) );
  XOR2_X1 U975 ( .A(n875), .B(n874), .Z(n877) );
  XNOR2_X1 U976 ( .A(KEYINPUT111), .B(G2474), .ZN(n876) );
  XNOR2_X1 U977 ( .A(n877), .B(n876), .ZN(n878) );
  XNOR2_X1 U978 ( .A(KEYINPUT41), .B(n878), .ZN(n880) );
  XNOR2_X1 U979 ( .A(n880), .B(n879), .ZN(G229) );
  NAND2_X1 U980 ( .A1(G124), .A2(n897), .ZN(n881) );
  XNOR2_X1 U981 ( .A(n881), .B(KEYINPUT44), .ZN(n883) );
  NAND2_X1 U982 ( .A1(n896), .A2(G112), .ZN(n882) );
  NAND2_X1 U983 ( .A1(n883), .A2(n882), .ZN(n887) );
  NAND2_X1 U984 ( .A1(G100), .A2(n900), .ZN(n885) );
  NAND2_X1 U985 ( .A1(G136), .A2(n902), .ZN(n884) );
  NAND2_X1 U986 ( .A1(n885), .A2(n884), .ZN(n886) );
  NOR2_X1 U987 ( .A1(n887), .A2(n886), .ZN(G162) );
  NAND2_X1 U988 ( .A1(G103), .A2(n900), .ZN(n889) );
  NAND2_X1 U989 ( .A1(G139), .A2(n902), .ZN(n888) );
  NAND2_X1 U990 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U991 ( .A(KEYINPUT113), .B(n890), .Z(n895) );
  NAND2_X1 U992 ( .A1(G115), .A2(n896), .ZN(n892) );
  NAND2_X1 U993 ( .A1(G127), .A2(n897), .ZN(n891) );
  NAND2_X1 U994 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U995 ( .A(KEYINPUT47), .B(n893), .Z(n894) );
  NOR2_X1 U996 ( .A1(n895), .A2(n894), .ZN(n1000) );
  NAND2_X1 U997 ( .A1(G118), .A2(n896), .ZN(n899) );
  NAND2_X1 U998 ( .A1(G130), .A2(n897), .ZN(n898) );
  NAND2_X1 U999 ( .A1(n899), .A2(n898), .ZN(n907) );
  NAND2_X1 U1000 ( .A1(n900), .A2(G106), .ZN(n901) );
  XNOR2_X1 U1001 ( .A(n901), .B(KEYINPUT112), .ZN(n904) );
  NAND2_X1 U1002 ( .A1(G142), .A2(n902), .ZN(n903) );
  NAND2_X1 U1003 ( .A1(n904), .A2(n903), .ZN(n905) );
  XOR2_X1 U1004 ( .A(KEYINPUT45), .B(n905), .Z(n906) );
  NOR2_X1 U1005 ( .A1(n907), .A2(n906), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n1000), .B(n908), .ZN(n920) );
  XOR2_X1 U1007 ( .A(G162), .B(n991), .Z(n911) );
  XNOR2_X1 U1008 ( .A(G160), .B(n909), .ZN(n910) );
  XNOR2_X1 U1009 ( .A(n911), .B(n910), .ZN(n915) );
  XOR2_X1 U1010 ( .A(KEYINPUT115), .B(KEYINPUT46), .Z(n913) );
  XNOR2_X1 U1011 ( .A(KEYINPUT114), .B(KEYINPUT48), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(n913), .B(n912), .ZN(n914) );
  XOR2_X1 U1013 ( .A(n915), .B(n914), .Z(n918) );
  XNOR2_X1 U1014 ( .A(G164), .B(n916), .ZN(n917) );
  XNOR2_X1 U1015 ( .A(n918), .B(n917), .ZN(n919) );
  XNOR2_X1 U1016 ( .A(n920), .B(n919), .ZN(n922) );
  XOR2_X1 U1017 ( .A(n922), .B(n921), .Z(n923) );
  NOR2_X1 U1018 ( .A1(G37), .A2(n923), .ZN(G395) );
  NOR2_X1 U1019 ( .A1(G227), .A2(G229), .ZN(n924) );
  XOR2_X1 U1020 ( .A(KEYINPUT117), .B(n924), .Z(n925) );
  XNOR2_X1 U1021 ( .A(n925), .B(KEYINPUT49), .ZN(n926) );
  NOR2_X1 U1022 ( .A1(G397), .A2(n926), .ZN(n930) );
  NOR2_X1 U1023 ( .A1(n931), .A2(G401), .ZN(n927) );
  XOR2_X1 U1024 ( .A(KEYINPUT116), .B(n927), .Z(n928) );
  NOR2_X1 U1025 ( .A1(G395), .A2(n928), .ZN(n929) );
  NAND2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(G225) );
  INV_X1 U1027 ( .A(G225), .ZN(G308) );
  INV_X1 U1028 ( .A(n931), .ZN(G319) );
  INV_X1 U1029 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1030 ( .A(G16), .B(KEYINPUT56), .ZN(n958) );
  XNOR2_X1 U1031 ( .A(G1966), .B(G168), .ZN(n933) );
  NAND2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1033 ( .A(n934), .B(KEYINPUT57), .ZN(n956) );
  XNOR2_X1 U1034 ( .A(G301), .B(G1961), .ZN(n937) );
  XNOR2_X1 U1035 ( .A(n935), .B(G1348), .ZN(n936) );
  NOR2_X1 U1036 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1037 ( .A(KEYINPUT120), .B(n938), .ZN(n950) );
  XNOR2_X1 U1038 ( .A(n939), .B(G1956), .ZN(n940) );
  XNOR2_X1 U1039 ( .A(n940), .B(KEYINPUT121), .ZN(n941) );
  NOR2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n944) );
  NAND2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n948) );
  XNOR2_X1 U1042 ( .A(G166), .B(G1971), .ZN(n946) );
  NAND2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n954) );
  XNOR2_X1 U1046 ( .A(G1341), .B(n951), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(KEYINPUT122), .B(n952), .ZN(n953) );
  NOR2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1050 ( .A1(n958), .A2(n957), .ZN(n986) );
  INV_X1 U1051 ( .A(G16), .ZN(n984) );
  XNOR2_X1 U1052 ( .A(G1348), .B(KEYINPUT59), .ZN(n959) );
  XNOR2_X1 U1053 ( .A(n959), .B(G4), .ZN(n963) );
  XNOR2_X1 U1054 ( .A(G1956), .B(G20), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(G6), .B(G1981), .ZN(n960) );
  NOR2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n966) );
  XOR2_X1 U1058 ( .A(KEYINPUT123), .B(G1341), .Z(n964) );
  XNOR2_X1 U1059 ( .A(G19), .B(n964), .ZN(n965) );
  NOR2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1061 ( .A(n967), .B(KEYINPUT60), .ZN(n970) );
  XOR2_X1 U1062 ( .A(G1966), .B(G21), .Z(n968) );
  XNOR2_X1 U1063 ( .A(KEYINPUT124), .B(n968), .ZN(n969) );
  NAND2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(KEYINPUT125), .B(n971), .ZN(n973) );
  XOR2_X1 U1066 ( .A(G1961), .B(G5), .Z(n972) );
  NAND2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n980) );
  XNOR2_X1 U1068 ( .A(G1971), .B(G22), .ZN(n975) );
  XNOR2_X1 U1069 ( .A(G23), .B(G1976), .ZN(n974) );
  NOR2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n977) );
  XOR2_X1 U1071 ( .A(G1986), .B(G24), .Z(n976) );
  NAND2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1073 ( .A(KEYINPUT58), .B(n978), .ZN(n979) );
  NOR2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1075 ( .A(n981), .B(KEYINPUT126), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(n982), .B(KEYINPUT61), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1079 ( .A(n987), .B(KEYINPUT127), .ZN(n1015) );
  XOR2_X1 U1080 ( .A(G2090), .B(G162), .Z(n988) );
  NOR2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n990) );
  XOR2_X1 U1082 ( .A(KEYINPUT51), .B(n990), .Z(n995) );
  NOR2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(n993), .B(KEYINPUT118), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n997) );
  XOR2_X1 U1086 ( .A(G160), .B(G2084), .Z(n996) );
  NOR2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1005) );
  XOR2_X1 U1089 ( .A(G2072), .B(n1000), .Z(n1002) );
  XOR2_X1 U1090 ( .A(G164), .B(G2078), .Z(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1092 ( .A(KEYINPUT50), .B(n1003), .Z(n1004) );
  NOR2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  NAND2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1096 ( .A(KEYINPUT52), .B(n1010), .ZN(n1012) );
  INV_X1 U1097 ( .A(KEYINPUT55), .ZN(n1011) );
  NAND2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1099 ( .A1(n1013), .A2(G29), .ZN(n1014) );
  NAND2_X1 U1100 ( .A1(n1015), .A2(n1014), .ZN(n1038) );
  XNOR2_X1 U1101 ( .A(G1996), .B(G32), .ZN(n1017) );
  XNOR2_X1 U1102 ( .A(G33), .B(G2072), .ZN(n1016) );
  NOR2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1025) );
  XOR2_X1 U1104 ( .A(G2067), .B(G26), .Z(n1018) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(G28), .ZN(n1023) );
  XOR2_X1 U1106 ( .A(n1019), .B(G27), .Z(n1021) );
  XOR2_X1 U1107 ( .A(G1991), .B(G25), .Z(n1020) );
  NAND2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1111 ( .A(n1026), .B(KEYINPUT53), .ZN(n1029) );
  XOR2_X1 U1112 ( .A(G2084), .B(G34), .Z(n1027) );
  XNOR2_X1 U1113 ( .A(KEYINPUT54), .B(n1027), .ZN(n1028) );
  NAND2_X1 U1114 ( .A1(n1029), .A2(n1028), .ZN(n1031) );
  XNOR2_X1 U1115 ( .A(G35), .B(G2090), .ZN(n1030) );
  NOR2_X1 U1116 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1117 ( .A(KEYINPUT55), .B(n1032), .ZN(n1034) );
  INV_X1 U1118 ( .A(G29), .ZN(n1033) );
  NAND2_X1 U1119 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1120 ( .A1(n1035), .A2(G11), .ZN(n1036) );
  XOR2_X1 U1121 ( .A(KEYINPUT119), .B(n1036), .Z(n1037) );
  NOR2_X1 U1122 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  XNOR2_X1 U1123 ( .A(KEYINPUT62), .B(n1039), .ZN(G311) );
  INV_X1 U1124 ( .A(G311), .ZN(G150) );
endmodule

