//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 1 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 1 0 1 0 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n209, new_n210, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1263,
    new_n1264, new_n1265;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NOR3_X1   g0007(.A1(new_n207), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0008(.A1(G97), .A2(G107), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G87), .ZN(G355));
  INV_X1    g0011(.A(G1), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G13), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT0), .Z(new_n219));
  INV_X1    g0019(.A(KEYINPUT1), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT66), .Z(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  AND3_X1   g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n214), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n219), .B1(new_n220), .B2(new_n227), .ZN(new_n228));
  OR2_X1    g0028(.A1(new_n207), .A2(KEYINPUT65), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n207), .A2(KEYINPUT65), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n229), .A2(G50), .A3(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n233), .A2(new_n213), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n228), .B(new_n235), .C1(new_n220), .C2(new_n227), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n236), .B(KEYINPUT67), .Z(G361));
  XOR2_X1   g0037(.A(G238), .B(G244), .Z(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT68), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G250), .B(G257), .Z(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n242), .B(new_n247), .Z(G358));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G50), .B(G68), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G58), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n251), .B(new_n254), .Z(G351));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G264), .A3(G1698), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n260), .A2(G257), .A3(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G303), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n261), .A2(new_n263), .A3(new_n267), .ZN(new_n268));
  AND2_X1   g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(new_n233), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G179), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n212), .A2(G13), .A3(G20), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G116), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n212), .A2(G33), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n273), .A2(new_n277), .A3(new_n233), .A4(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n276), .B1(new_n279), .B2(new_n275), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G283), .ZN(new_n281));
  INV_X1    g0081(.A(G97), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n281), .B(new_n213), .C1(G33), .C2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n278), .A2(new_n233), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n275), .A2(G20), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT20), .ZN(new_n287));
  OR2_X1    g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n287), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n280), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n272), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT82), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT5), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n292), .B1(new_n293), .B2(G41), .ZN(new_n294));
  INV_X1    g0094(.A(G41), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n295), .A2(KEYINPUT82), .A3(KEYINPUT5), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n293), .A2(G41), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT81), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n298), .A2(new_n299), .A3(new_n212), .A4(G45), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(KEYINPUT71), .B1(new_n269), .B2(new_n233), .ZN(new_n302));
  NAND2_X1  g0102(.A1(G33), .A2(G41), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT71), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n303), .A2(new_n304), .A3(G1), .A4(G13), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n295), .A2(KEYINPUT5), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n212), .A2(G45), .ZN(new_n308));
  OAI21_X1  g0108(.A(KEYINPUT81), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n301), .A2(G274), .A3(new_n306), .A4(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n297), .A2(new_n300), .A3(new_n309), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT84), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n311), .A2(new_n306), .A3(new_n312), .A4(G270), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n311), .A2(new_n306), .A3(G270), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT84), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n291), .A2(KEYINPUT85), .A3(new_n314), .A4(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT85), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n316), .A2(new_n310), .A3(new_n313), .ZN(new_n319));
  INV_X1    g0119(.A(G179), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n320), .B1(new_n268), .B2(new_n270), .ZN(new_n321));
  XNOR2_X1  g0121(.A(new_n286), .B(KEYINPUT20), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n321), .B1(new_n322), .B2(new_n280), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n318), .B1(new_n319), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n317), .A2(new_n324), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n314), .A2(G190), .A3(new_n316), .A4(new_n271), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n316), .A2(new_n310), .A3(new_n313), .A4(new_n271), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G200), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n326), .A2(new_n328), .A3(new_n290), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT21), .ZN(new_n330));
  INV_X1    g0130(.A(G169), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n290), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n330), .B1(new_n327), .B2(new_n332), .ZN(new_n333));
  AND3_X1   g0133(.A1(new_n327), .A2(new_n330), .A3(new_n332), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n325), .B(new_n329), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(G1698), .B1(new_n258), .B2(new_n259), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G222), .ZN(new_n338));
  INV_X1    g0138(.A(G77), .ZN(new_n339));
  INV_X1    g0139(.A(G223), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n260), .A2(G1698), .ZN(new_n341));
  OAI221_X1 g0141(.A(new_n338), .B1(new_n339), .B2(new_n260), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n270), .ZN(new_n343));
  INV_X1    g0143(.A(G45), .ZN(new_n344));
  AOI21_X1  g0144(.A(G1), .B1(new_n295), .B2(new_n344), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n302), .A2(G274), .A3(new_n305), .A4(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n345), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n348), .A2(new_n302), .A3(new_n305), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT72), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n348), .A2(new_n302), .A3(KEYINPUT72), .A4(new_n305), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n347), .B1(G226), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G190), .ZN(new_n355));
  INV_X1    g0155(.A(G50), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n213), .B1(new_n206), .B2(new_n356), .ZN(new_n357));
  XNOR2_X1  g0157(.A(KEYINPUT8), .B(G58), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n213), .A2(G33), .ZN(new_n359));
  INV_X1    g0159(.A(G150), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n213), .A2(new_n257), .ZN(new_n361));
  OAI22_X1  g0161(.A1(new_n358), .A2(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n284), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n212), .A2(G20), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(G50), .ZN(new_n365));
  XOR2_X1   g0165(.A(new_n365), .B(KEYINPUT73), .Z(new_n366));
  NOR2_X1   g0166(.A1(new_n274), .A2(new_n284), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  OAI221_X1 g0168(.A(new_n363), .B1(G50), .B2(new_n273), .C1(new_n366), .C2(new_n368), .ZN(new_n369));
  XNOR2_X1  g0169(.A(new_n369), .B(KEYINPUT9), .ZN(new_n370));
  INV_X1    g0170(.A(G200), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n355), .B(new_n370), .C1(new_n371), .C2(new_n354), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n372), .B(KEYINPUT10), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT16), .ZN(new_n374));
  INV_X1    g0174(.A(G159), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n361), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G58), .A2(G68), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n204), .A2(new_n205), .A3(new_n377), .ZN(new_n378));
  AOI211_X1 g0178(.A(new_n374), .B(new_n376), .C1(new_n378), .C2(G20), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT7), .ZN(new_n380));
  NOR4_X1   g0180(.A1(new_n264), .A2(new_n265), .A3(new_n380), .A4(G20), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT77), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(new_n264), .B2(new_n265), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n258), .A2(KEYINPUT77), .A3(new_n259), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(new_n384), .A3(new_n213), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n381), .B1(new_n385), .B2(new_n380), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n379), .B1(new_n386), .B2(new_n203), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n258), .A2(new_n213), .A3(new_n259), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n380), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n266), .A2(KEYINPUT7), .A3(new_n213), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n203), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n378), .A2(G20), .ZN(new_n392));
  INV_X1    g0192(.A(new_n376), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n374), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n387), .A2(new_n284), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n358), .B1(new_n212), .B2(G20), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n397), .A2(new_n367), .B1(new_n274), .B2(new_n358), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G232), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n346), .B1(new_n349), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n270), .ZN(new_n402));
  MUX2_X1   g0202(.A(G223), .B(G226), .S(G1698), .Z(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n260), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G87), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n402), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n331), .B1(new_n401), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n404), .A2(new_n405), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT78), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(new_n409), .A3(new_n270), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n403), .A2(new_n260), .B1(G33), .B2(G87), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT78), .B1(new_n411), .B2(new_n402), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n346), .B(new_n320), .C1(new_n349), .C2(new_n400), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n407), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n399), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT18), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n371), .B1(new_n401), .B2(new_n406), .ZN(new_n419));
  INV_X1    g0219(.A(G190), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n346), .B(new_n420), .C1(new_n349), .C2(new_n400), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n419), .B1(new_n413), .B2(new_n421), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n422), .A2(new_n396), .A3(new_n398), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT17), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n415), .B1(new_n396), .B2(new_n398), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT18), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n422), .A2(new_n396), .A3(new_n398), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT17), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n418), .A2(new_n424), .A3(new_n427), .A4(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n354), .A2(new_n320), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n433), .B(new_n369), .C1(G169), .C2(new_n354), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n260), .A2(G232), .A3(new_n262), .ZN(new_n435));
  INV_X1    g0235(.A(G107), .ZN(new_n436));
  INV_X1    g0236(.A(G238), .ZN(new_n437));
  OAI221_X1 g0237(.A(new_n435), .B1(new_n436), .B2(new_n260), .C1(new_n341), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n270), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n346), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n353), .A2(G244), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n320), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n367), .A2(G77), .A3(new_n364), .ZN(new_n444));
  XNOR2_X1  g0244(.A(KEYINPUT15), .B(G87), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(new_n359), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(KEYINPUT74), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT74), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n445), .A2(new_n448), .A3(new_n359), .ZN(new_n449));
  OAI22_X1  g0249(.A1(new_n358), .A2(new_n361), .B1(new_n213), .B2(new_n339), .ZN(new_n450));
  NOR3_X1   g0250(.A1(new_n447), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n284), .ZN(new_n452));
  OAI221_X1 g0252(.A(new_n444), .B1(G77), .B2(new_n273), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n331), .B1(new_n440), .B2(new_n441), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n443), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(G200), .B1(new_n440), .B2(new_n441), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n453), .B1(new_n442), .B2(G190), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n373), .A2(new_n432), .A3(new_n434), .A4(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT76), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n461), .B1(new_n273), .B2(G68), .ZN(new_n462));
  XNOR2_X1  g0262(.A(new_n462), .B(KEYINPUT12), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT11), .ZN(new_n464));
  OAI22_X1  g0264(.A1(new_n359), .A2(new_n339), .B1(new_n213), .B2(G68), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n361), .A2(new_n356), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n284), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n463), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  OR2_X1    g0268(.A1(new_n467), .A2(new_n464), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n367), .A2(G68), .A3(new_n364), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  OAI211_X1 g0272(.A(G232), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G97), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT75), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n337), .A2(new_n476), .A3(G226), .ZN(new_n477));
  OAI211_X1 g0277(.A(G226), .B(new_n262), .C1(new_n264), .C2(new_n265), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT75), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n475), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  OR2_X1    g0280(.A1(new_n480), .A2(new_n402), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT13), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n353), .A2(G238), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n481), .A2(new_n482), .A3(new_n483), .A4(new_n346), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n346), .B1(new_n480), .B2(new_n402), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n437), .B1(new_n351), .B2(new_n352), .ZN(new_n486));
  OAI21_X1  g0286(.A(KEYINPUT13), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT14), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n488), .A2(new_n489), .A3(G169), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n484), .A2(G179), .A3(new_n487), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n489), .B1(new_n488), .B2(G169), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n472), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n471), .B1(new_n488), .B2(new_n420), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n371), .B1(new_n484), .B2(new_n487), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n460), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n337), .A2(KEYINPUT4), .A3(G244), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n260), .A2(G250), .A3(G1698), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n501), .A2(new_n281), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(KEYINPUT4), .B1(new_n337), .B2(G244), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n270), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n311), .A2(new_n306), .A3(G257), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n505), .A2(new_n420), .A3(new_n310), .A4(new_n506), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n505), .A2(new_n310), .A3(new_n506), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n507), .B1(new_n508), .B2(G200), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n274), .A2(KEYINPUT80), .A3(new_n282), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT80), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n273), .B2(G97), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n510), .B(new_n512), .C1(new_n282), .C2(new_n279), .ZN(new_n513));
  AOI21_X1  g0313(.A(KEYINPUT7), .B1(new_n266), .B2(new_n213), .ZN(new_n514));
  OAI21_X1  g0314(.A(G107), .B1(new_n514), .B2(new_n381), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT6), .ZN(new_n516));
  AND2_X1   g0316(.A1(G97), .A2(G107), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n516), .B1(new_n517), .B2(new_n209), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n436), .A2(KEYINPUT6), .A3(G97), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n361), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n520), .A2(G20), .B1(G77), .B2(new_n521), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n515), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(KEYINPUT79), .B1(new_n523), .B2(new_n452), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n452), .B1(new_n515), .B2(new_n522), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT79), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n513), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n509), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n508), .A2(new_n320), .ZN(new_n530));
  INV_X1    g0330(.A(new_n513), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n525), .A2(new_n526), .ZN(new_n532));
  AOI211_X1 g0332(.A(KEYINPUT79), .B(new_n452), .C1(new_n515), .C2(new_n522), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n505), .A2(new_n310), .A3(new_n506), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n331), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n530), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G33), .A2(G116), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n538), .A2(G20), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n213), .A2(G107), .ZN(new_n540));
  OR2_X1    g0340(.A1(new_n540), .A2(KEYINPUT23), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(KEYINPUT23), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n539), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n260), .A2(new_n213), .A3(G87), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT22), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n545), .A2(KEYINPUT86), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n544), .A2(new_n546), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n543), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n549), .A2(KEYINPUT24), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT24), .ZN(new_n551));
  XNOR2_X1  g0351(.A(new_n544), .B(new_n546), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n551), .B1(new_n552), .B2(new_n543), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n284), .B1(new_n550), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n215), .A2(G1), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n540), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n556), .A2(KEYINPUT87), .A3(KEYINPUT25), .ZN(new_n557));
  OR2_X1    g0357(.A1(KEYINPUT87), .A2(KEYINPUT25), .ZN(new_n558));
  NAND2_X1  g0358(.A1(KEYINPUT87), .A2(KEYINPUT25), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n555), .A2(new_n540), .A3(new_n558), .A4(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n557), .B(new_n560), .C1(new_n436), .C2(new_n279), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n337), .A2(G250), .B1(G33), .B2(G294), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n260), .A2(G257), .A3(G1698), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n270), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n311), .A2(new_n306), .A3(G264), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n566), .A2(new_n310), .A3(G190), .A4(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n310), .A3(new_n567), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(G200), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n554), .A2(new_n562), .A3(new_n568), .A4(new_n570), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n529), .A2(new_n537), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n337), .A2(G238), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n260), .A2(G244), .A3(G1698), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(new_n538), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n270), .ZN(new_n576));
  MUX2_X1   g0376(.A(G274), .B(G250), .S(new_n308), .Z(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n306), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n331), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n260), .A2(new_n213), .A3(G68), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT19), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n213), .B1(new_n474), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(G87), .B2(new_n210), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n213), .A2(G33), .A3(G97), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n585), .A2(KEYINPUT83), .A3(new_n582), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT83), .B1(new_n585), .B2(new_n582), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n581), .B(new_n584), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n588), .A2(new_n284), .B1(new_n274), .B2(new_n445), .ZN(new_n589));
  INV_X1    g0389(.A(new_n279), .ZN(new_n590));
  INV_X1    g0390(.A(new_n445), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n575), .A2(new_n270), .B1(new_n577), .B2(new_n306), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n320), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n580), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n579), .A2(new_n420), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n590), .A2(G87), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n589), .B(new_n598), .C1(new_n594), .C2(new_n371), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n596), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  OR2_X1    g0400(.A1(new_n569), .A2(G179), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n569), .A2(new_n331), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n554), .A2(new_n562), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n600), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AND4_X1   g0405(.A1(new_n336), .A2(new_n500), .A3(new_n572), .A4(new_n605), .ZN(G372));
  NAND3_X1  g0406(.A1(new_n498), .A2(new_n430), .A3(new_n424), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n607), .B1(new_n494), .B2(new_n455), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n418), .A2(new_n427), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n373), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n610), .A2(new_n434), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n549), .A2(KEYINPUT24), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n552), .A2(new_n551), .A3(new_n543), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n452), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n601), .B(new_n602), .C1(new_n614), .C2(new_n561), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n615), .B(new_n325), .C1(new_n333), .C2(new_n334), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n596), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT88), .ZN(new_n619));
  OR2_X1    g0419(.A1(new_n599), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n597), .B1(new_n599), .B2(new_n619), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n618), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n622), .A2(new_n537), .A3(new_n529), .A4(new_n571), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n596), .B1(new_n617), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n537), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT26), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n622), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n537), .A2(new_n600), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n627), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n500), .B1(new_n624), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n611), .A2(new_n630), .ZN(G369));
  NAND2_X1  g0431(.A1(new_n555), .A2(new_n213), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(G213), .A3(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(G343), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n638), .A2(new_n290), .ZN(new_n639));
  XNOR2_X1  g0439(.A(new_n639), .B(KEYINPUT89), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n336), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n334), .A2(new_n333), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n324), .B2(new_n317), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n641), .B1(new_n643), .B2(new_n640), .ZN(new_n644));
  XOR2_X1   g0444(.A(new_n644), .B(KEYINPUT90), .Z(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(G330), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n604), .A2(new_n637), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n648), .A2(new_n571), .B1(new_n603), .B2(new_n604), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n615), .A2(new_n637), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n643), .A2(new_n637), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n650), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n652), .A2(new_n654), .ZN(G399));
  NOR2_X1   g0455(.A1(new_n216), .A2(G41), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n210), .A2(G87), .A3(G116), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(G1), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n231), .B2(new_n657), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(KEYINPUT28), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n620), .A2(new_n621), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n596), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT26), .B1(new_n663), .B2(new_n537), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n628), .A2(new_n626), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  OAI211_X1 g0466(.A(KEYINPUT29), .B(new_n638), .C1(new_n624), .C2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(KEYINPUT91), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n667), .A2(KEYINPUT91), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n638), .B1(new_n624), .B2(new_n629), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT29), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n668), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n336), .A2(new_n572), .A3(new_n605), .A4(new_n638), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n594), .A2(G179), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n327), .A2(new_n535), .A3(new_n675), .A4(new_n569), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n594), .A2(new_n321), .A3(new_n566), .A4(new_n567), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n677), .A2(new_n535), .A3(new_n319), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n676), .B1(new_n678), .B2(KEYINPUT30), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n677), .A2(new_n535), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT30), .ZN(new_n681));
  NOR3_X1   g0481(.A1(new_n680), .A2(new_n681), .A3(new_n319), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n637), .B1(new_n679), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT31), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI211_X1 g0485(.A(KEYINPUT31), .B(new_n637), .C1(new_n679), .C2(new_n682), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n674), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(G330), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n673), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n661), .B1(new_n690), .B2(G1), .ZN(G364));
  NOR2_X1   g0491(.A1(new_n215), .A2(G20), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n212), .B1(new_n692), .B2(G45), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n656), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n647), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(G330), .B2(new_n645), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n217), .A2(G355), .A3(new_n260), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(G116), .B2(new_n217), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n232), .A2(new_n344), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n383), .A2(new_n384), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(new_n216), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n703), .B1(G45), .B2(new_n254), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n699), .B1(new_n700), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(G20), .B1(KEYINPUT92), .B2(G169), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(KEYINPUT92), .A2(G169), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n233), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(G13), .A2(G33), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(G20), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n695), .B1(new_n705), .B2(new_n714), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n420), .A2(G179), .A3(G200), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(new_n213), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n213), .A2(new_n320), .ZN(new_n718));
  NOR2_X1   g0518(.A1(G190), .A2(G200), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OAI22_X1  g0520(.A1(new_n717), .A2(new_n282), .B1(new_n720), .B2(new_n339), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n718), .A2(G190), .A3(new_n371), .ZN(new_n722));
  XOR2_X1   g0522(.A(new_n722), .B(KEYINPUT93), .Z(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n721), .B1(new_n724), .B2(G58), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n213), .A2(G179), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n726), .A2(new_n420), .A3(G200), .ZN(new_n727));
  INV_X1    g0527(.A(G87), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n726), .A2(G190), .A3(G200), .ZN(new_n729));
  OAI221_X1 g0529(.A(new_n260), .B1(new_n727), .B2(new_n436), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT94), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n718), .A2(G200), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n420), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(G190), .ZN(new_n734));
  AOI22_X1  g0534(.A1(G50), .A2(new_n733), .B1(new_n734), .B2(G68), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n726), .A2(new_n719), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n375), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT32), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n725), .A2(new_n731), .A3(new_n735), .A4(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n722), .ZN(new_n740));
  INV_X1    g0540(.A(new_n736), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n740), .A2(G322), .B1(new_n741), .B2(G329), .ZN(new_n742));
  INV_X1    g0542(.A(G283), .ZN(new_n743));
  INV_X1    g0543(.A(new_n734), .ZN(new_n744));
  XOR2_X1   g0544(.A(KEYINPUT33), .B(G317), .Z(new_n745));
  OAI221_X1 g0545(.A(new_n742), .B1(new_n743), .B2(new_n727), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(G303), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n266), .B1(new_n729), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n746), .B1(KEYINPUT96), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n749), .B1(KEYINPUT96), .B2(new_n748), .ZN(new_n750));
  INV_X1    g0550(.A(G294), .ZN(new_n751));
  INV_X1    g0551(.A(G311), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n717), .A2(new_n751), .B1(new_n720), .B2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n753), .B1(G326), .B2(new_n733), .ZN(new_n754));
  XOR2_X1   g0554(.A(new_n754), .B(KEYINPUT95), .Z(new_n755));
  OAI21_X1  g0555(.A(new_n739), .B1(new_n750), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n715), .B1(new_n756), .B2(new_n709), .ZN(new_n757));
  XOR2_X1   g0557(.A(new_n712), .B(KEYINPUT97), .Z(new_n758));
  OAI21_X1  g0558(.A(new_n757), .B1(new_n644), .B2(new_n758), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n697), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(G396));
  NOR2_X1   g0561(.A1(new_n455), .A2(new_n637), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n458), .A2(new_n457), .B1(new_n453), .B2(new_n637), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n763), .B1(new_n456), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n670), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n765), .ZN(new_n767));
  OAI211_X1 g0567(.A(new_n767), .B(new_n638), .C1(new_n624), .C2(new_n629), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n695), .B1(new_n769), .B2(new_n688), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n770), .B1(new_n688), .B2(new_n769), .ZN(new_n771));
  INV_X1    g0571(.A(new_n695), .ZN(new_n772));
  INV_X1    g0572(.A(new_n709), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(new_n711), .ZN(new_n774));
  XOR2_X1   g0574(.A(new_n774), .B(KEYINPUT98), .Z(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n772), .B1(new_n776), .B2(new_n339), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n260), .B1(new_n741), .B2(G311), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n778), .B1(new_n275), .B2(new_n720), .C1(new_n751), .C2(new_n722), .ZN(new_n779));
  INV_X1    g0579(.A(new_n727), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n733), .A2(G303), .B1(new_n780), .B2(G87), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(new_n436), .B2(new_n729), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n744), .A2(new_n743), .B1(new_n282), .B2(new_n717), .ZN(new_n783));
  NOR3_X1   g0583(.A1(new_n779), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n720), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n733), .A2(G137), .B1(new_n785), .B2(G159), .ZN(new_n786));
  INV_X1    g0586(.A(G143), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n786), .B1(new_n360), .B2(new_n744), .C1(new_n723), .C2(new_n787), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n788), .B(KEYINPUT34), .Z(new_n789));
  NOR2_X1   g0589(.A1(new_n727), .A2(new_n203), .ZN(new_n790));
  INV_X1    g0590(.A(new_n729), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n790), .B1(G50), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT99), .ZN(new_n793));
  INV_X1    g0593(.A(new_n717), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G58), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n741), .A2(G132), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n793), .A2(new_n701), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n789), .B1(KEYINPUT100), .B2(new_n797), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n797), .A2(KEYINPUT100), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n784), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n777), .B1(new_n800), .B2(new_n773), .C1(new_n767), .C2(new_n711), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n771), .A2(new_n801), .ZN(G384));
  NAND3_X1  g0602(.A1(new_n232), .A2(G77), .A3(new_n377), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n356), .A2(G68), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n212), .B(G13), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n520), .A2(KEYINPUT35), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n520), .A2(KEYINPUT35), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n806), .A2(G116), .A3(new_n234), .A4(new_n807), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(KEYINPUT36), .Z(new_n809));
  NOR2_X1   g0609(.A1(new_n805), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT40), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n385), .A2(new_n380), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n390), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G68), .ZN(new_n814));
  INV_X1    g0614(.A(new_n394), .ZN(new_n815));
  AOI21_X1  g0615(.A(KEYINPUT16), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n387), .A2(new_n284), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n398), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(KEYINPUT101), .ZN(new_n819));
  INV_X1    g0619(.A(new_n635), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT101), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n821), .B(new_n398), .C1(new_n816), .C2(new_n817), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n819), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n432), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n819), .A2(new_n416), .A3(new_n822), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n823), .A2(new_n825), .A3(new_n428), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT102), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n826), .A2(new_n827), .A3(KEYINPUT37), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n423), .A2(new_n425), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT37), .ZN(new_n830));
  AOI211_X1 g0630(.A(KEYINPUT103), .B(new_n635), .C1(new_n396), .C2(new_n398), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT103), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(new_n399), .B2(new_n820), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n829), .B(new_n830), .C1(new_n831), .C2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n828), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n827), .B1(new_n826), .B2(KEYINPUT37), .ZN(new_n836));
  OAI211_X1 g0636(.A(KEYINPUT38), .B(new_n824), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n826), .A2(KEYINPUT37), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(KEYINPUT102), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n840), .A2(new_n834), .A3(new_n828), .ZN(new_n841));
  AOI21_X1  g0641(.A(KEYINPUT38), .B1(new_n841), .B2(new_n824), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n472), .A2(new_n637), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n494), .A2(new_n498), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n488), .A2(G169), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(KEYINPUT14), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n847), .A2(new_n491), .A3(new_n490), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n472), .B(new_n637), .C1(new_n848), .C2(new_n497), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n765), .B1(new_n845), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(KEYINPUT106), .B1(new_n850), .B2(new_n687), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n850), .A2(KEYINPUT106), .A3(new_n687), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n811), .B1(new_n843), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n833), .A2(new_n831), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n417), .A2(new_n428), .ZN(new_n857));
  OAI21_X1  g0657(.A(KEYINPUT37), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n834), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n431), .A2(new_n856), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT38), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n861), .A2(KEYINPUT104), .A3(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT104), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n858), .A2(new_n834), .B1(new_n431), .B2(new_n856), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n864), .B1(new_n865), .B2(KEYINPUT38), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n837), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n845), .A2(new_n849), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n869), .A2(new_n687), .A3(new_n767), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n870), .A2(new_n811), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n855), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n500), .A2(new_n687), .ZN(new_n874));
  OAI21_X1  g0674(.A(G330), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(new_n873), .B2(new_n874), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n848), .A2(new_n472), .A3(new_n638), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT39), .B1(new_n838), .B2(new_n842), .ZN(new_n878));
  XOR2_X1   g0678(.A(KEYINPUT105), .B(KEYINPUT39), .Z(new_n879));
  NAND3_X1  g0679(.A1(new_n867), .A2(new_n837), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n877), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n609), .A2(new_n635), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n768), .A2(new_n763), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n869), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n882), .B1(new_n843), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n500), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n611), .B1(new_n673), .B2(new_n887), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n886), .B(new_n888), .ZN(new_n889));
  OAI22_X1  g0689(.A1(new_n876), .A2(new_n889), .B1(new_n212), .B2(new_n692), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n876), .A2(new_n889), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n810), .B1(new_n890), .B2(new_n891), .ZN(G367));
  XOR2_X1   g0692(.A(new_n656), .B(KEYINPUT41), .Z(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n529), .B(new_n537), .C1(new_n528), .C2(new_n638), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n625), .A2(new_n637), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n654), .A2(new_n897), .ZN(new_n898));
  XOR2_X1   g0698(.A(new_n898), .B(KEYINPUT45), .Z(new_n899));
  NOR2_X1   g0699(.A1(new_n654), .A2(new_n897), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT44), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n652), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n646), .A2(new_n650), .A3(new_n649), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n899), .A2(new_n901), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n651), .B(new_n653), .Z(new_n907));
  XNOR2_X1  g0707(.A(new_n646), .B(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n690), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n894), .B1(new_n910), .B2(new_n689), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n693), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n903), .A2(new_n897), .ZN(new_n913));
  OR2_X1    g0713(.A1(new_n895), .A2(new_n615), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n637), .B1(new_n914), .B2(new_n537), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n651), .A2(new_n653), .A3(new_n897), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n915), .B1(new_n916), .B2(KEYINPUT42), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n916), .A2(KEYINPUT42), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n589), .A2(new_n598), .ZN(new_n919));
  OR3_X1    g0719(.A1(new_n596), .A2(new_n919), .A3(new_n638), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n919), .A2(new_n638), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n920), .B1(new_n663), .B2(new_n921), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n917), .A2(new_n918), .B1(KEYINPUT43), .B2(new_n922), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n922), .A2(KEYINPUT43), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n923), .B(new_n924), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n913), .B(new_n925), .Z(new_n926));
  NAND2_X1  g0726(.A1(new_n912), .A2(new_n926), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n247), .A2(new_n702), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n713), .B1(new_n217), .B2(new_n445), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n695), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n780), .A2(G77), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n260), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n932), .B(KEYINPUT107), .Z(new_n933));
  AOI22_X1  g0733(.A1(G50), .A2(new_n785), .B1(new_n741), .B2(G137), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n360), .B2(new_n722), .ZN(new_n935));
  INV_X1    g0735(.A(new_n733), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n787), .A2(new_n936), .B1(new_n744), .B2(new_n375), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n717), .A2(new_n203), .B1(new_n729), .B2(new_n202), .ZN(new_n938));
  NOR4_X1   g0738(.A1(new_n933), .A2(new_n935), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT108), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n724), .A2(G303), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n744), .A2(new_n751), .B1(new_n436), .B2(new_n717), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n780), .A2(G97), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n936), .B2(new_n752), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(G317), .ZN(new_n946));
  OAI22_X1  g0746(.A1(new_n720), .A2(new_n743), .B1(new_n736), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n947), .A2(new_n701), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n791), .A2(G116), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT46), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n941), .A2(new_n945), .A3(new_n948), .A4(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n940), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT47), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n930), .B1(new_n953), .B2(new_n709), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n758), .B2(new_n922), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n927), .A2(new_n955), .ZN(G387));
  AOI21_X1  g0756(.A(new_n657), .B1(new_n908), .B2(new_n690), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n690), .B2(new_n908), .ZN(new_n958));
  INV_X1    g0758(.A(new_n658), .ZN(new_n959));
  AOI211_X1 g0759(.A(G45), .B(new_n959), .C1(G68), .C2(G77), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT110), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OR3_X1    g0762(.A1(new_n358), .A2(KEYINPUT50), .A3(G50), .ZN(new_n963));
  OAI21_X1  g0763(.A(KEYINPUT50), .B1(new_n358), .B2(G50), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n960), .A2(new_n961), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n702), .B1(new_n344), .B2(new_n242), .C1(new_n965), .C2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n959), .A2(new_n217), .A3(new_n260), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(G107), .B2(new_n217), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT109), .Z(new_n970));
  AND2_X1   g0770(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n695), .B1(new_n714), .B2(new_n971), .C1(new_n651), .C2(new_n758), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n717), .A2(new_n445), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n791), .A2(G77), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n744), .B2(new_n358), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n973), .B(new_n975), .C1(G159), .C2(new_n733), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n722), .A2(new_n356), .B1(new_n720), .B2(new_n203), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(G150), .B2(new_n741), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n976), .A2(new_n701), .A3(new_n943), .A4(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT111), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n724), .A2(G317), .B1(G303), .B2(new_n785), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n981), .A2(KEYINPUT113), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(KEYINPUT113), .ZN(new_n983));
  AOI22_X1  g0783(.A1(G311), .A2(new_n734), .B1(new_n733), .B2(G322), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT48), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n717), .A2(new_n743), .B1(new_n729), .B2(new_n751), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT112), .Z(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(new_n985), .B2(new_n986), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n987), .A2(KEYINPUT49), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n701), .B1(G326), .B2(new_n741), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n991), .B(new_n992), .C1(new_n275), .C2(new_n727), .ZN(new_n993));
  AOI21_X1  g0793(.A(KEYINPUT49), .B1(new_n987), .B2(new_n990), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n980), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT114), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n972), .B1(new_n996), .B2(new_n709), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(new_n908), .B2(new_n694), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n958), .A2(new_n998), .ZN(G393));
  INV_X1    g0799(.A(KEYINPUT115), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n902), .A2(new_n1000), .A3(new_n905), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n903), .A2(new_n904), .A3(KEYINPUT115), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n693), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n895), .A2(new_n896), .A3(new_n712), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n936), .A2(new_n946), .B1(new_n752), .B2(new_n722), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT52), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n266), .B1(new_n720), .B2(new_n751), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(G322), .B2(new_n741), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n791), .A2(G283), .B1(new_n780), .B2(G107), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(G116), .A2(new_n794), .B1(new_n734), .B2(G303), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1006), .A2(new_n1008), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n936), .A2(new_n360), .B1(new_n375), .B2(new_n722), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT51), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n358), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n1014), .A2(new_n785), .B1(new_n741), .B2(G143), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n717), .A2(new_n339), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n203), .A2(new_n729), .B1(new_n727), .B2(new_n728), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n1016), .B(new_n1017), .C1(G50), .C2(new_n734), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1013), .A2(new_n701), .A3(new_n1015), .A4(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n773), .B1(new_n1011), .B2(new_n1019), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n703), .A2(new_n251), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n714), .B1(G97), .B2(new_n216), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n772), .B(new_n1020), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1003), .B1(new_n1004), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1001), .A2(new_n909), .A3(new_n1002), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1025), .B(new_n656), .C1(new_n909), .C2(new_n906), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1024), .A2(new_n1026), .ZN(G390));
  INV_X1    g0827(.A(G330), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n686), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n681), .B1(new_n680), .B2(new_n319), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n678), .A2(KEYINPUT30), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1030), .A2(new_n1031), .A3(new_n676), .ZN(new_n1032));
  AOI21_X1  g0832(.A(KEYINPUT31), .B1(new_n1032), .B2(new_n637), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1029), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1028), .B1(new_n1034), .B2(new_n674), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n500), .A2(new_n1035), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n611), .B(new_n1036), .C1(new_n673), .C2(new_n887), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n687), .A2(G330), .A3(new_n767), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n869), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT117), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1038), .A2(KEYINPUT117), .A3(new_n1039), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT116), .ZN(new_n1044));
  AND3_X1   g0844(.A1(new_n1035), .A2(new_n1044), .A3(new_n850), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1044), .B1(new_n1035), .B2(new_n850), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1042), .B(new_n1043), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n883), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n626), .B1(new_n622), .B2(new_n625), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n626), .B2(new_n628), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n529), .A2(new_n537), .A3(new_n571), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1051), .A2(new_n663), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n618), .B1(new_n1052), .B2(new_n616), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n637), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n764), .A2(new_n456), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n762), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1035), .A2(new_n850), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1057), .A2(new_n1058), .A3(new_n1040), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1037), .B1(new_n1048), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n884), .A2(new_n877), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n878), .A2(new_n1061), .A3(new_n880), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n868), .B(new_n877), .C1(new_n1039), .C2(new_n1057), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1062), .A2(new_n1063), .A3(new_n1058), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1060), .B(new_n1064), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT118), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1060), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1059), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n1047), .B2(new_n883), .ZN(new_n1071));
  OAI21_X1  g0871(.A(KEYINPUT118), .B1(new_n1071), .B2(new_n1037), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1073));
  AND3_X1   g0873(.A1(new_n1062), .A2(new_n1063), .A3(new_n1058), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1066), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n656), .B(new_n1067), .C1(new_n1073), .C2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n878), .A2(new_n880), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1078), .A2(new_n711), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G97), .A2(new_n785), .B1(new_n741), .B2(G294), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1080), .B(new_n266), .C1(new_n275), .C2(new_n722), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n790), .B(new_n1081), .C1(G87), .C2(new_n791), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n744), .A2(new_n436), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1016), .B(new_n1083), .C1(G283), .C2(new_n733), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(KEYINPUT54), .B(G143), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n785), .A2(new_n1086), .B1(new_n741), .B2(G125), .ZN(new_n1087));
  INV_X1    g0887(.A(G132), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1087), .B(new_n260), .C1(new_n1088), .C2(new_n722), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n734), .A2(G137), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n356), .B2(new_n727), .ZN(new_n1091));
  INV_X1    g0891(.A(G128), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n936), .A2(new_n1092), .B1(new_n375), .B2(new_n717), .ZN(new_n1093));
  NOR3_X1   g0893(.A1(new_n1089), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n729), .A2(new_n360), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT53), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n1082), .A2(new_n1084), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n695), .B1(new_n1014), .B2(new_n775), .C1(new_n1097), .C2(new_n773), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1079), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(new_n1076), .B2(new_n694), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1077), .A2(new_n1100), .ZN(G378));
  INV_X1    g0901(.A(KEYINPUT123), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1028), .B1(new_n868), .B2(new_n871), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n373), .A2(new_n434), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n369), .A2(new_n820), .ZN(new_n1105));
  XOR2_X1   g0905(.A(new_n1105), .B(KEYINPUT121), .Z(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  XOR2_X1   g0907(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1108));
  INV_X1    g0908(.A(new_n1106), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n373), .A2(new_n434), .A3(new_n1109), .ZN(new_n1110));
  AND3_X1   g0910(.A1(new_n1107), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1108), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n855), .A2(new_n1103), .A3(new_n1114), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n850), .A2(KEYINPUT106), .A3(new_n687), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1116), .A2(new_n851), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n824), .B1(new_n835), .B2(new_n836), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n862), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n837), .ZN(new_n1120));
  AOI21_X1  g0920(.A(KEYINPUT40), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n872), .A2(G330), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1113), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  AND3_X1   g0923(.A1(new_n886), .A2(new_n1115), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n877), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1078), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n884), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1127), .A2(new_n1120), .B1(new_n609), .B2(new_n635), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n1115), .A2(new_n1123), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1102), .B1(new_n1124), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1037), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1067), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1114), .B1(new_n855), .B2(new_n1103), .ZN(new_n1134));
  NOR3_X1   g0934(.A1(new_n1121), .A2(new_n1122), .A3(new_n1113), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1133), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n886), .A2(new_n1115), .A3(new_n1123), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1136), .A2(KEYINPUT123), .A3(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1130), .A2(new_n1132), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT57), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1037), .B1(new_n1076), .B2(new_n1060), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1136), .A2(KEYINPUT57), .A3(new_n1137), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n656), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1141), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1130), .A2(new_n694), .A3(new_n1138), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n936), .A2(new_n275), .B1(new_n203), .B2(new_n717), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT119), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n701), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n295), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n974), .B1(new_n202), .B2(new_n727), .C1(new_n744), .C2(new_n282), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n591), .A2(new_n785), .B1(new_n741), .B2(G283), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(new_n436), .B2(new_n722), .ZN(new_n1154));
  NOR4_X1   g0954(.A1(new_n1149), .A2(new_n1151), .A3(new_n1152), .A4(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1155), .B(new_n1156), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1151), .B(new_n356), .C1(G33), .C2(G41), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n733), .A2(G125), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n744), .B2(new_n1088), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n740), .A2(G128), .B1(new_n785), .B2(G137), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n729), .B2(new_n1085), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1160), .B(new_n1162), .C1(G150), .C2(new_n794), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1164), .A2(KEYINPUT59), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(KEYINPUT59), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n780), .A2(G159), .ZN(new_n1167));
  AOI211_X1 g0967(.A(G33), .B(G41), .C1(new_n741), .C2(G124), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1157), .B(new_n1158), .C1(new_n1165), .C2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n709), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1171), .B(new_n695), .C1(G50), .C2(new_n775), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n1114), .B2(new_n710), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT122), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1147), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1146), .A2(new_n1176), .ZN(G375));
  OAI22_X1  g0977(.A1(new_n275), .A2(new_n744), .B1(new_n936), .B2(new_n751), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G97), .B2(new_n791), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n973), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n722), .A2(new_n743), .B1(new_n720), .B2(new_n436), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n260), .B(new_n1181), .C1(G303), .C2(new_n741), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1179), .A2(new_n931), .A3(new_n1180), .A4(new_n1182), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n936), .A2(new_n1088), .B1(new_n729), .B2(new_n375), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(G50), .B2(new_n794), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n724), .A2(G137), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n720), .A2(new_n360), .B1(new_n736), .B2(new_n1092), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1150), .A2(new_n1187), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n734), .A2(new_n1086), .B1(new_n780), .B2(G58), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1185), .A2(new_n1186), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n773), .B1(new_n1183), .B2(new_n1190), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n772), .B(new_n1191), .C1(new_n203), .C2(new_n776), .ZN(new_n1192));
  XOR2_X1   g0992(.A(new_n1192), .B(KEYINPUT124), .Z(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n711), .B2(new_n869), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n1071), .B2(new_n693), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1071), .A2(new_n1037), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n894), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1196), .B1(new_n1073), .B2(new_n1198), .ZN(G381));
  INV_X1    g0999(.A(G387), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n958), .A2(new_n760), .A3(new_n998), .ZN(new_n1201));
  NOR3_X1   g1001(.A1(G390), .A2(new_n1201), .A3(G384), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  OR4_X1    g1003(.A1(G378), .A2(new_n1203), .A3(G375), .A4(G381), .ZN(G407));
  AOI21_X1  g1004(.A(new_n1175), .B1(new_n1141), .B2(new_n1145), .ZN(new_n1205));
  INV_X1    g1005(.A(G378), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n636), .A2(G213), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT125), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1205), .A2(new_n1206), .A3(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(G407), .A2(G213), .A3(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT126), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(G407), .A2(KEYINPUT126), .A3(G213), .A4(new_n1209), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(G409));
  NAND2_X1  g1014(.A1(new_n1200), .A2(G390), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1201), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n760), .B1(new_n958), .B2(new_n998), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(G387), .A2(new_n1026), .A3(new_n1024), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1215), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1218), .B1(new_n1215), .B2(new_n1219), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1208), .ZN(new_n1224));
  OAI21_X1  g1024(.A(KEYINPUT60), .B1(new_n1071), .B2(new_n1037), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n1197), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1071), .A2(KEYINPUT60), .A3(new_n1037), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1226), .A2(new_n656), .A3(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n1196), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1229), .A2(new_n771), .A3(new_n801), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1228), .A2(G384), .A3(new_n1196), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1144), .B1(new_n1140), .B2(new_n1139), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(new_n1234), .A2(new_n1206), .A3(new_n1175), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1130), .A2(new_n1132), .A3(new_n894), .A4(new_n1138), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1136), .A2(new_n694), .A3(new_n1137), .ZN(new_n1237));
  AND2_X1   g1037(.A1(new_n1237), .A2(new_n1174), .ZN(new_n1238));
  AOI21_X1  g1038(.A(G378), .B1(new_n1236), .B2(new_n1238), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1224), .B(new_n1233), .C1(new_n1235), .C2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT127), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1146), .A2(G378), .A3(new_n1176), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1239), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1208), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1245), .A2(KEYINPUT127), .A3(new_n1233), .ZN(new_n1246));
  AOI21_X1  g1046(.A(KEYINPUT62), .B1(new_n1242), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1208), .A2(G2897), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n1232), .B(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1239), .B1(new_n1205), .B2(G378), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1249), .B1(new_n1250), .B2(new_n1208), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT61), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n1208), .B(new_n1232), .C1(new_n1243), .C2(new_n1244), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT62), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1251), .B(new_n1252), .C1(new_n1253), .C2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1223), .B1(new_n1247), .B2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT63), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1242), .A2(new_n1246), .A3(new_n1257), .ZN(new_n1258));
  AND2_X1   g1058(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1253), .A2(KEYINPUT63), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1258), .A2(new_n1259), .A3(new_n1222), .A4(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1256), .A2(new_n1261), .ZN(G405));
  NAND2_X1  g1062(.A1(G375), .A2(new_n1206), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1243), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1264), .B(new_n1232), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1265), .B(new_n1222), .ZN(G402));
endmodule


