//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 1 0 1 0 0 1 0 0 0 0 1 0 0 1 1 0 0 0 0 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 1 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n564, new_n565, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XOR2_X1   g014(.A(KEYINPUT67), .B(G120), .Z(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT68), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n448));
  AND2_X1   g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  NAND2_X1  g025(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(KEYINPUT70), .B(KEYINPUT2), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n453), .B(new_n454), .Z(new_n455));
  OR4_X1    g030(.A1(G237), .A2(G236), .A3(G235), .A4(G238), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n455), .A2(new_n456), .ZN(G325));
  XNOR2_X1  g032(.A(G325), .B(KEYINPUT71), .ZN(G261));
  NAND2_X1  g033(.A1(new_n455), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT72), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT72), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(new_n467), .A3(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n469));
  AND4_X1   g044(.A1(new_n463), .A2(new_n465), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G137), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n467), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(new_n469), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n464), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G101), .ZN(new_n479));
  AND3_X1   g054(.A1(new_n471), .A2(new_n477), .A3(new_n479), .ZN(G160));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n482));
  OR2_X1    g057(.A1(new_n470), .A2(KEYINPUT73), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n470), .A2(KEYINPUT73), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(G136), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n482), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NOR3_X1   g063(.A1(new_n464), .A2(KEYINPUT72), .A3(KEYINPUT3), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n467), .A2(G2104), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n491), .A2(G2105), .A3(new_n465), .ZN(new_n492));
  XNOR2_X1  g067(.A(new_n492), .B(KEYINPUT74), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n488), .B1(G124), .B2(new_n493), .ZN(G162));
  AND2_X1   g069(.A1(KEYINPUT4), .A2(G138), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n473), .A2(new_n469), .A3(G138), .A4(new_n463), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n470), .A2(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(G114), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  AND2_X1   g078(.A1(G126), .A2(G2105), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n465), .A2(new_n468), .A3(new_n469), .A4(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT75), .ZN(new_n506));
  AND2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n505), .A2(new_n506), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n503), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT76), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n491), .A2(KEYINPUT75), .A3(new_n465), .A4(new_n504), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n505), .A2(new_n506), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n502), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT76), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n499), .B1(new_n511), .B2(new_n515), .ZN(G164));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G50), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT5), .ZN(new_n521));
  OAI21_X1  g096(.A(KEYINPUT77), .B1(new_n521), .B2(G543), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT77), .ZN(new_n523));
  INV_X1    g098(.A(G543), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(new_n524), .A3(KEYINPUT5), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n521), .A2(G543), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(new_n517), .ZN(new_n529));
  INV_X1    g104(.A(G88), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n520), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n528), .A2(G62), .ZN(new_n533));
  NAND2_X1  g108(.A1(G75), .A2(G543), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT78), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n532), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n531), .A2(new_n536), .ZN(G303));
  INV_X1    g112(.A(G303), .ZN(G166));
  AND2_X1   g113(.A1(new_n528), .A2(new_n517), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G89), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n528), .A2(G63), .A3(G651), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n519), .A2(G51), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n541), .A2(KEYINPUT79), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT7), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n540), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g121(.A(KEYINPUT79), .B1(new_n541), .B2(new_n542), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n546), .A2(new_n547), .ZN(G168));
  XNOR2_X1  g123(.A(KEYINPUT80), .B(G52), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n539), .A2(G90), .B1(new_n519), .B2(new_n549), .ZN(new_n550));
  XOR2_X1   g125(.A(new_n550), .B(KEYINPUT81), .Z(new_n551));
  AOI22_X1  g126(.A1(new_n528), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(new_n532), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n551), .A2(new_n553), .ZN(G301));
  INV_X1    g129(.A(G301), .ZN(G171));
  AOI22_X1  g130(.A1(new_n528), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n556), .A2(new_n532), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n519), .A2(G43), .ZN(new_n558));
  INV_X1    g133(.A(G81), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n529), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND4_X1  g140(.A1(G319), .A2(G483), .A3(G661), .A4(new_n565), .ZN(G188));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n526), .A2(new_n527), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OR2_X1    g145(.A1(new_n570), .A2(KEYINPUT82), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(KEYINPUT82), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n571), .A2(G651), .A3(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(G53), .ZN(new_n574));
  OR3_X1    g149(.A1(new_n518), .A2(KEYINPUT9), .A3(new_n574), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT9), .B1(new_n518), .B2(new_n574), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n539), .A2(G91), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n573), .A2(new_n577), .ZN(G299));
  INV_X1    g153(.A(G168), .ZN(G286));
  OAI21_X1  g154(.A(G651), .B1(new_n528), .B2(G74), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT83), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n539), .A2(G87), .B1(G49), .B2(new_n519), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G288));
  AOI22_X1  g158(.A1(new_n528), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n532), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n519), .A2(G48), .ZN(new_n586));
  INV_X1    g161(.A(G86), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n529), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G305));
  AOI22_X1  g165(.A1(new_n539), .A2(G85), .B1(G47), .B2(new_n519), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n528), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n532), .B2(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(new_n539), .A2(G92), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n594), .B(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  XNOR2_X1  g172(.A(KEYINPUT84), .B(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n568), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n599), .A2(G651), .B1(G54), .B2(new_n519), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G171), .B2(new_n602), .ZN(G284));
  OAI21_X1  g179(.A(new_n603), .B1(G171), .B2(new_n602), .ZN(G321));
  NAND2_X1  g180(.A1(G299), .A2(new_n602), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(new_n602), .B2(G168), .ZN(G297));
  OAI21_X1  g182(.A(new_n606), .B1(new_n602), .B2(G168), .ZN(G280));
  AND2_X1   g183(.A1(new_n596), .A2(new_n600), .ZN(new_n609));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G860), .ZN(G148));
  NAND2_X1  g186(.A1(new_n609), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n613), .A2(KEYINPUT85), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(KEYINPUT85), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n614), .B(new_n615), .C1(G868), .C2(new_n561), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n485), .A2(G135), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n493), .A2(G123), .ZN(new_n619));
  NOR3_X1   g194(.A1(new_n463), .A2(KEYINPUT87), .A3(G111), .ZN(new_n620));
  OAI21_X1  g195(.A(KEYINPUT87), .B1(new_n463), .B2(G111), .ZN(new_n621));
  OR2_X1    g196(.A1(G99), .A2(G2105), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n621), .A2(G2104), .A3(new_n622), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n618), .B(new_n619), .C1(new_n620), .C2(new_n623), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n624), .A2(G2096), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(G2096), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT86), .B(G2100), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT12), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n628), .B(new_n630), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n625), .A2(new_n626), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT88), .ZN(G156));
  XNOR2_X1  g208(.A(G2427), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n637), .A2(new_n638), .A3(KEYINPUT14), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n639), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2451), .B(G2454), .Z(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT89), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n643), .A2(new_n646), .ZN(new_n648));
  AND3_X1   g223(.A1(new_n647), .A2(G14), .A3(new_n648), .ZN(G401));
  XOR2_X1   g224(.A(G2072), .B(G2078), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT90), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT17), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2084), .B(G2090), .ZN(new_n654));
  NOR3_X1   g229(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n654), .B1(new_n651), .B2(new_n653), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n656), .B1(new_n652), .B2(new_n653), .ZN(new_n657));
  INV_X1    g232(.A(new_n653), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n658), .A2(new_n654), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n651), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT18), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n655), .A2(new_n657), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2096), .B(G2100), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(G227));
  XNOR2_X1  g239(.A(G1971), .B(G1976), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1956), .B(G2474), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1961), .B(G1966), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n669), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n667), .A2(KEYINPUT92), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n673), .B(new_n674), .Z(new_n675));
  NOR3_X1   g250(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT20), .Z(new_n677));
  NAND2_X1  g252(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT93), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n680), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G1981), .B(G1986), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G229));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G23), .ZN(new_n687));
  INV_X1    g262(.A(G288), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n687), .B1(new_n688), .B2(new_n686), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT98), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT33), .B(G1976), .Z(new_n691));
  AND2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n686), .A2(G6), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(new_n589), .B2(new_n686), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT32), .B(G1981), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT97), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n695), .B(new_n697), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n686), .A2(KEYINPUT96), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n686), .A2(KEYINPUT96), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n701), .A2(G22), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(G166), .B2(new_n701), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G1971), .ZN(new_n704));
  OR4_X1    g279(.A1(new_n692), .A2(new_n693), .A3(new_n698), .A4(new_n704), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n705), .A2(KEYINPUT34), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(KEYINPUT34), .ZN(new_n707));
  INV_X1    g282(.A(G25), .ZN(new_n708));
  OR3_X1    g283(.A1(new_n708), .A2(KEYINPUT94), .A3(G29), .ZN(new_n709));
  OAI21_X1  g284(.A(KEYINPUT94), .B1(new_n708), .B2(G29), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n485), .A2(G131), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT95), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  OAI21_X1  g288(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n714));
  INV_X1    g289(.A(G107), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(G2105), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n493), .B2(G119), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n709), .B(new_n710), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT35), .B(G1991), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  MUX2_X1   g298(.A(G24), .B(G290), .S(new_n701), .Z(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(G1986), .Z(new_n725));
  NAND4_X1  g300(.A1(new_n706), .A2(new_n707), .A3(new_n723), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT36), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n686), .A2(G4), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n609), .B2(new_n686), .ZN(new_n729));
  INV_X1    g304(.A(G1348), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n686), .A2(G21), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G168), .B2(new_n686), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n731), .B1(G1966), .B2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G34), .ZN(new_n735));
  AOI21_X1  g310(.A(G29), .B1(new_n735), .B2(KEYINPUT24), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(KEYINPUT24), .B2(new_n735), .ZN(new_n737));
  INV_X1    g312(.A(G160), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(new_n720), .ZN(new_n739));
  INV_X1    g314(.A(G2084), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT30), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n742), .A2(G28), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n720), .B1(new_n742), .B2(G28), .ZN(new_n744));
  AND2_X1   g319(.A1(KEYINPUT31), .A2(G11), .ZN(new_n745));
  NOR2_X1   g320(.A1(KEYINPUT31), .A2(G11), .ZN(new_n746));
  OAI22_X1  g321(.A1(new_n743), .A2(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AND3_X1   g322(.A1(new_n699), .A2(G19), .A3(new_n700), .ZN(new_n748));
  INV_X1    g323(.A(new_n561), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(new_n701), .ZN(new_n750));
  INV_X1    g325(.A(G1341), .ZN(new_n751));
  AOI211_X1 g326(.A(new_n741), .B(new_n747), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  OAI221_X1 g327(.A(new_n752), .B1(new_n720), .B2(new_n624), .C1(new_n751), .C2(new_n750), .ZN(new_n753));
  NAND3_X1  g328(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT26), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n478), .A2(G105), .ZN(new_n756));
  AOI211_X1 g331(.A(new_n755), .B(new_n756), .C1(new_n493), .C2(G129), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n485), .A2(G141), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n759), .A2(new_n720), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n720), .B2(G32), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT27), .B(G1996), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n720), .A2(G27), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G164), .B2(new_n720), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G2078), .ZN(new_n766));
  NOR4_X1   g341(.A1(new_n734), .A2(new_n753), .A3(new_n763), .A4(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n699), .A2(G20), .A3(new_n700), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT23), .Z(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G299), .B2(G16), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G1956), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n733), .A2(G1966), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT101), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n686), .A2(G5), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G171), .B2(new_n686), .ZN(new_n775));
  INV_X1    g350(.A(G1961), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n767), .A2(new_n771), .A3(new_n773), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(G115), .A2(G2104), .ZN(new_n779));
  INV_X1    g354(.A(G127), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n474), .B2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT25), .ZN(new_n782));
  NAND2_X1  g357(.A1(G103), .A2(G2104), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(G2105), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n463), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n785));
  AOI22_X1  g360(.A1(new_n781), .A2(G2105), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(G139), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n486), .B2(new_n787), .ZN(new_n788));
  MUX2_X1   g363(.A(G33), .B(new_n788), .S(G29), .Z(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(G2072), .Z(new_n790));
  NAND2_X1  g365(.A1(new_n761), .A2(new_n762), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n790), .B(new_n791), .C1(new_n740), .C2(new_n739), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT100), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n720), .A2(G26), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT28), .Z(new_n795));
  OAI21_X1  g370(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n796));
  INV_X1    g371(.A(G116), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(G2105), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n485), .B2(G140), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT99), .ZN(new_n800));
  AND3_X1   g375(.A1(new_n493), .A2(new_n800), .A3(G128), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n800), .B1(new_n493), .B2(G128), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n799), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n795), .B1(new_n803), .B2(G29), .ZN(new_n804));
  INV_X1    g379(.A(G2067), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n720), .A2(G35), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G162), .B2(new_n720), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT29), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G2090), .ZN(new_n810));
  NOR4_X1   g385(.A1(new_n778), .A2(new_n793), .A3(new_n806), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n727), .A2(new_n811), .ZN(G150));
  INV_X1    g387(.A(G150), .ZN(G311));
  NAND2_X1  g388(.A1(new_n609), .A2(G559), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT38), .ZN(new_n815));
  NAND2_X1  g390(.A1(G80), .A2(G543), .ZN(new_n816));
  INV_X1    g391(.A(G67), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n568), .B2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT102), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n532), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(new_n819), .B2(new_n818), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n539), .A2(G93), .B1(G55), .B2(new_n519), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(new_n561), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n821), .A2(new_n822), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n749), .A2(new_n825), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n815), .B(new_n827), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n828), .A2(KEYINPUT39), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n828), .A2(KEYINPUT39), .ZN(new_n830));
  NOR3_X1   g405(.A1(new_n829), .A2(new_n830), .A3(G860), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n825), .A2(G860), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT37), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n831), .A2(new_n833), .ZN(G145));
  INV_X1    g409(.A(new_n630), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n713), .A2(new_n835), .A3(new_n717), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n835), .B1(new_n713), .B2(new_n717), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n493), .A2(G130), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT103), .ZN(new_n840));
  OR2_X1    g415(.A1(G106), .A2(G2105), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n841), .B(G2104), .C1(G118), .C2(new_n463), .ZN(new_n842));
  INV_X1    g417(.A(G142), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n842), .B1(new_n486), .B2(new_n843), .ZN(new_n844));
  OAI22_X1  g419(.A1(new_n837), .A2(new_n838), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n838), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n840), .A2(new_n844), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n846), .A2(new_n847), .A3(new_n836), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n759), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n803), .A2(new_n788), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n514), .A2(new_n498), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n803), .A2(new_n788), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n853), .B1(new_n852), .B2(new_n854), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n851), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n857), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n859), .A2(new_n759), .A3(new_n855), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n850), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT105), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n850), .A2(new_n858), .A3(KEYINPUT105), .A4(new_n860), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n624), .B(new_n738), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(G162), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n858), .A2(new_n860), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n867), .B1(new_n868), .B2(new_n849), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n863), .A2(new_n864), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(KEYINPUT106), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT106), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n863), .A2(new_n872), .A3(new_n869), .A4(new_n864), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT104), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n861), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n876), .A2(new_n866), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n868), .A2(new_n849), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n878), .A2(new_n861), .A3(new_n875), .ZN(new_n879));
  AOI21_X1  g454(.A(G37), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n874), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g457(.A(new_n609), .B1(KEYINPUT107), .B2(G299), .ZN(new_n883));
  INV_X1    g458(.A(G299), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT107), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n601), .B1(new_n885), .B2(new_n884), .ZN(new_n888));
  INV_X1    g463(.A(new_n886), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n824), .A2(new_n826), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n612), .B(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT108), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n891), .A2(KEYINPUT108), .A3(new_n893), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT41), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n898), .B1(new_n887), .B2(new_n890), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n883), .A2(new_n886), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n888), .A2(new_n889), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n900), .A2(new_n901), .A3(KEYINPUT41), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  OAI211_X1 g478(.A(new_n896), .B(new_n897), .C1(new_n893), .C2(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XOR2_X1   g483(.A(G290), .B(G303), .Z(new_n909));
  XNOR2_X1  g484(.A(G288), .B(new_n589), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n909), .B(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n911), .B1(KEYINPUT109), .B2(KEYINPUT42), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n908), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n906), .A2(new_n912), .A3(new_n907), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(G868), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT110), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n823), .A2(G868), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n917), .A2(new_n918), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n602), .B1(new_n914), .B2(new_n915), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT110), .B1(new_n922), .B2(new_n919), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(G295));
  NAND2_X1  g499(.A1(new_n917), .A2(new_n920), .ZN(G331));
  INV_X1    g500(.A(KEYINPUT111), .ZN(new_n926));
  NAND2_X1  g501(.A1(G171), .A2(new_n892), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n827), .A2(G301), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(G286), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n927), .A2(new_n928), .A3(G168), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n930), .A2(new_n899), .A3(new_n902), .A4(new_n931), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n927), .A2(new_n928), .A3(G168), .ZN(new_n933));
  AOI21_X1  g508(.A(G168), .B1(new_n927), .B2(new_n928), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n891), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n911), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n926), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n932), .A2(new_n935), .A3(KEYINPUT111), .A4(new_n911), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(G37), .B1(new_n936), .B2(new_n937), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n940), .A2(new_n944), .A3(new_n941), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  XOR2_X1   g521(.A(new_n946), .B(KEYINPUT44), .Z(G397));
  NAND2_X1  g522(.A1(G160), .A2(G40), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G1384), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n853), .A2(new_n950), .ZN(new_n951));
  XOR2_X1   g526(.A(KEYINPUT112), .B(KEYINPUT45), .Z(new_n952));
  AND3_X1   g527(.A1(new_n949), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  XOR2_X1   g528(.A(new_n718), .B(new_n722), .Z(new_n954));
  XNOR2_X1  g529(.A(new_n759), .B(G1996), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n803), .B(new_n805), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(G290), .B(G1986), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n953), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT125), .ZN(new_n962));
  INV_X1    g537(.A(G8), .ZN(new_n963));
  NOR2_X1   g538(.A1(G168), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT116), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n966), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT115), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n951), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT50), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n853), .A2(KEYINPUT115), .A3(new_n950), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n967), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n512), .A2(new_n513), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT76), .B1(new_n974), .B2(new_n503), .ZN(new_n975));
  AOI211_X1 g550(.A(new_n510), .B(new_n502), .C1(new_n512), .C2(new_n513), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n498), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n950), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n966), .B1(new_n978), .B2(KEYINPUT50), .ZN(new_n979));
  XOR2_X1   g554(.A(KEYINPUT121), .B(G2084), .Z(new_n980));
  NAND2_X1  g555(.A1(new_n949), .A2(new_n980), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n973), .A2(new_n979), .A3(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT115), .B1(new_n853), .B2(new_n950), .ZN(new_n984));
  AOI211_X1 g559(.A(new_n968), .B(G1384), .C1(new_n514), .C2(new_n498), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n952), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n977), .A2(new_n950), .A3(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n986), .A2(new_n988), .A3(new_n949), .ZN(new_n989));
  INV_X1    g564(.A(G1966), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT123), .B1(new_n982), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n511), .A2(new_n515), .ZN(new_n993));
  AOI21_X1  g568(.A(G1384), .B1(new_n993), .B2(new_n498), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT116), .B1(new_n994), .B2(new_n970), .ZN(new_n995));
  INV_X1    g570(.A(new_n981), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n995), .A2(new_n972), .A3(new_n967), .A4(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n989), .A2(new_n990), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT123), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n965), .B1(new_n992), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n963), .B1(new_n992), .B2(new_n1000), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT124), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n965), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AND3_X1   g579(.A1(new_n997), .A2(new_n999), .A3(new_n998), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n999), .B1(new_n997), .B2(new_n998), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1003), .B(G8), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT51), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(G8), .B1(new_n982), .B2(new_n991), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(new_n1011), .A3(new_n965), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1001), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1013));
  OR3_X1    g588(.A1(new_n585), .A2(new_n588), .A3(G1981), .ZN(new_n1014));
  OAI21_X1  g589(.A(G1981), .B1(new_n585), .B2(new_n588), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1014), .A2(KEYINPUT49), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT49), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n984), .A2(new_n985), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n963), .B1(new_n1019), .B2(new_n949), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT119), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT119), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1018), .A2(new_n1023), .A3(new_n1020), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1976), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1020), .B1(new_n1026), .B2(G288), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT52), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n688), .A2(G1976), .ZN(new_n1029));
  OR3_X1    g604(.A1(new_n1027), .A2(KEYINPUT52), .A3(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1025), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(G303), .A2(G8), .ZN(new_n1032));
  XOR2_X1   g607(.A(new_n1032), .B(KEYINPUT55), .Z(new_n1033));
  AOI21_X1  g608(.A(new_n948), .B1(new_n994), .B2(new_n970), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n970), .B2(new_n1019), .ZN(new_n1035));
  XOR2_X1   g610(.A(KEYINPUT117), .B(G2090), .Z(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n949), .B1(new_n951), .B2(new_n983), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1038), .B1(new_n952), .B2(new_n978), .ZN(new_n1039));
  XOR2_X1   g614(.A(KEYINPUT113), .B(G1971), .Z(new_n1040));
  OAI22_X1  g615(.A1(new_n1035), .A2(new_n1037), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1033), .B1(new_n1041), .B2(G8), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1031), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1044), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1040), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n994), .A2(new_n987), .ZN(new_n1047));
  OAI211_X1 g622(.A(KEYINPUT114), .B(new_n1046), .C1(new_n1047), .C2(new_n1038), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1049));
  NOR4_X1   g624(.A1(new_n973), .A2(new_n979), .A3(new_n948), .A4(new_n1037), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT118), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n973), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1052), .A2(new_n949), .A3(new_n995), .A4(new_n1036), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(new_n1045), .A4(new_n1048), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1051), .A2(new_n1055), .A3(G8), .A4(new_n1033), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1043), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G2078), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT53), .B1(new_n1039), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1052), .A2(new_n949), .A3(new_n995), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1059), .B1(new_n1060), .B2(new_n776), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1058), .A2(KEYINPUT53), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1061), .B1(new_n989), .B2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g638(.A(G301), .B(KEYINPUT54), .ZN(new_n1064));
  AOI211_X1 g639(.A(new_n1062), .B(new_n1038), .C1(new_n951), .C2(new_n952), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1063), .A2(new_n1064), .B1(new_n1061), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1057), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n962), .B1(new_n1013), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1001), .ZN(new_n1070));
  OAI21_X1  g645(.A(G8), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n964), .B1(new_n1071), .B2(KEYINPUT124), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1011), .B1(new_n1072), .B2(new_n1007), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1012), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1070), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1075), .A2(KEYINPUT125), .A3(new_n1057), .A4(new_n1067), .ZN(new_n1076));
  INV_X1    g651(.A(G1956), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT56), .B(G2072), .ZN(new_n1078));
  AOI22_X1  g653(.A1(new_n1035), .A2(new_n1077), .B1(new_n1039), .B2(new_n1078), .ZN(new_n1079));
  XOR2_X1   g654(.A(G299), .B(KEYINPUT57), .Z(new_n1080));
  NOR2_X1   g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1082), .A2(new_n601), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1060), .A2(new_n730), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1019), .A2(new_n949), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1084), .B1(G2067), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1081), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT60), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n601), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT61), .ZN(new_n1091));
  OR3_X1    g666(.A1(new_n1082), .A2(new_n1081), .A3(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1091), .B1(new_n1082), .B2(new_n1081), .ZN(new_n1093));
  INV_X1    g668(.A(G1996), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1039), .A2(new_n1094), .ZN(new_n1095));
  XOR2_X1   g670(.A(KEYINPUT58), .B(G1341), .Z(new_n1096));
  NAND2_X1  g671(.A1(new_n1085), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n749), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  XOR2_X1   g673(.A(new_n1098), .B(KEYINPUT59), .Z(new_n1099));
  NAND4_X1  g674(.A1(new_n1090), .A2(new_n1092), .A3(new_n1093), .A4(new_n1099), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1101), .A2(new_n1089), .A3(new_n601), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1087), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1069), .A2(new_n1076), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1071), .A2(KEYINPUT124), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1105), .A2(new_n1007), .A3(new_n965), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1074), .B1(new_n1106), .B2(KEYINPUT51), .ZN(new_n1107));
  OAI21_X1  g682(.A(KEYINPUT62), .B1(new_n1107), .B2(new_n1001), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1057), .A2(G171), .A3(new_n1063), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT62), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1110), .B(new_n1070), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1108), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  AOI211_X1 g687(.A(G1976), .B(G288), .C1(new_n1022), .C2(new_n1024), .ZN(new_n1113));
  XOR2_X1   g688(.A(new_n1014), .B(KEYINPUT120), .Z(new_n1114));
  OAI21_X1  g689(.A(new_n1020), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n1056), .B2(new_n1031), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1010), .A2(G286), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1056), .A2(KEYINPUT63), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1033), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1051), .A2(G8), .A3(new_n1055), .ZN(new_n1120));
  AOI211_X1 g695(.A(KEYINPUT122), .B(new_n1031), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1119), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1031), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1122), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1118), .B1(new_n1121), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT63), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1043), .A2(new_n1056), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1117), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1127), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1116), .B1(new_n1126), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1112), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n961), .B1(new_n1104), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n956), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n953), .B1(new_n1134), .B2(new_n851), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n953), .A2(new_n1094), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1136), .B(KEYINPUT46), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  XOR2_X1   g713(.A(new_n1138), .B(KEYINPUT47), .Z(new_n1139));
  NAND2_X1  g714(.A1(new_n719), .A2(new_n722), .ZN(new_n1140));
  OAI22_X1  g715(.A1(new_n957), .A2(new_n1140), .B1(G2067), .B2(new_n803), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n953), .ZN(new_n1142));
  XOR2_X1   g717(.A(new_n1142), .B(KEYINPUT126), .Z(new_n1143));
  NAND2_X1  g718(.A1(new_n959), .A2(new_n953), .ZN(new_n1144));
  NOR2_X1   g719(.A1(G290), .A2(G1986), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n953), .A2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(KEYINPUT48), .ZN(new_n1147));
  AOI211_X1 g722(.A(new_n1139), .B(new_n1143), .C1(new_n1144), .C2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1133), .A2(new_n1148), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g724(.A1(G227), .A2(new_n461), .ZN(new_n1151));
  OR3_X1    g725(.A1(G229), .A2(G401), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g726(.A(new_n1152), .B1(new_n874), .B2(new_n880), .ZN(new_n1153));
  INV_X1    g727(.A(KEYINPUT127), .ZN(new_n1154));
  AND3_X1   g728(.A1(new_n946), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g729(.A(new_n1154), .B1(new_n946), .B2(new_n1153), .ZN(new_n1156));
  NOR2_X1   g730(.A1(new_n1155), .A2(new_n1156), .ZN(G308));
  NAND2_X1  g731(.A1(new_n946), .A2(new_n1153), .ZN(G225));
endmodule


