//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 1 0 1 1 0 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n851, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT70), .ZN(new_n203));
  INV_X1    g002(.A(G113gat), .ZN(new_n204));
  OAI21_X1  g003(.A(KEYINPUT68), .B1(new_n204), .B2(G120gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT68), .ZN(new_n206));
  INV_X1    g005(.A(G120gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(new_n207), .A3(G113gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n204), .A2(G120gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n205), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(G127gat), .A2(G134gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT69), .ZN(new_n213));
  NAND2_X1  g012(.A1(G127gat), .A2(G134gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n214), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT69), .B1(new_n216), .B2(new_n211), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT1), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n210), .A2(new_n215), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G134gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT67), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT67), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G134gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n223), .A3(G127gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(G113gat), .B(G120gat), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n224), .B(new_n212), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n219), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G190gat), .ZN(new_n228));
  AND2_X1   g027(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT27), .B(G183gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n235), .A2(new_n228), .A3(new_n232), .ZN(new_n236));
  NAND2_X1  g035(.A1(G183gat), .A2(G190gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n234), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n240));
  NAND2_X1  g039(.A1(G169gat), .A2(G176gat), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n240), .B1(new_n239), .B2(new_n241), .ZN(new_n243));
  NOR3_X1   g042(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n244));
  NOR3_X1   g043(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n238), .A2(new_n245), .ZN(new_n246));
  AND2_X1   g045(.A1(G169gat), .A2(G176gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(G169gat), .A2(G176gat), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n247), .B1(KEYINPUT23), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(G183gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(new_n228), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n251), .A2(KEYINPUT24), .A3(new_n237), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT23), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n253), .B1(G169gat), .B2(G176gat), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT24), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(G183gat), .A3(G190gat), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n249), .A2(new_n252), .A3(new_n254), .A4(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT25), .ZN(new_n258));
  INV_X1    g057(.A(G169gat), .ZN(new_n259));
  INV_X1    g058(.A(G176gat), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n259), .A2(new_n260), .A3(KEYINPUT23), .ZN(new_n261));
  AND4_X1   g060(.A1(KEYINPUT25), .A2(new_n261), .A3(new_n254), .A4(new_n241), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT64), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n237), .A2(new_n263), .A3(new_n255), .ZN(new_n264));
  OAI211_X1 g063(.A(G183gat), .B(G190gat), .C1(KEYINPUT64), .C2(KEYINPUT24), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(new_n251), .A3(new_n265), .ZN(new_n266));
  AOI22_X1  g065(.A1(new_n257), .A2(new_n258), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n227), .B1(new_n246), .B2(new_n267), .ZN(new_n268));
  AND2_X1   g067(.A1(new_n219), .A2(new_n226), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n256), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n261), .A2(new_n254), .A3(new_n241), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n258), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n262), .A2(new_n266), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n243), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n276));
  INV_X1    g075(.A(new_n244), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n231), .A2(new_n233), .B1(G183gat), .B2(G190gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n278), .A2(new_n236), .A3(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n269), .A2(new_n274), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n268), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(G227gat), .ZN(new_n283));
  INV_X1    g082(.A(G233gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n203), .B1(new_n282), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n285), .ZN(new_n287));
  AOI211_X1 g086(.A(KEYINPUT70), .B(new_n287), .C1(new_n268), .C2(new_n281), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT32), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT33), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n290), .B1(new_n286), .B2(new_n288), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT71), .B(G71gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n292), .B(G99gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(G15gat), .B(G43gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n289), .A2(new_n291), .A3(new_n296), .ZN(new_n297));
  OAI221_X1 g096(.A(KEYINPUT32), .B1(new_n290), .B2(new_n295), .C1(new_n286), .C2(new_n288), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n268), .A2(new_n281), .A3(new_n287), .ZN(new_n300));
  XOR2_X1   g099(.A(new_n300), .B(KEYINPUT34), .Z(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT72), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n297), .A2(new_n301), .A3(new_n298), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n301), .B1(new_n297), .B2(new_n298), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT72), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n202), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT36), .B1(new_n303), .B2(new_n305), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT78), .ZN(new_n311));
  INV_X1    g110(.A(G148gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n311), .A2(new_n312), .A3(G141gat), .ZN(new_n313));
  INV_X1    g112(.A(G141gat), .ZN(new_n314));
  AOI21_X1  g113(.A(KEYINPUT78), .B1(new_n314), .B2(G148gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(G148gat), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n313), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT79), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI211_X1 g118(.A(KEYINPUT79), .B(new_n313), .C1(new_n315), .C2(new_n316), .ZN(new_n320));
  NOR2_X1   g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT2), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G155gat), .A2(G162gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n319), .A2(new_n320), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT76), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n327), .B1(G155gat), .B2(G162gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n324), .A2(KEYINPUT76), .ZN(new_n329));
  NOR3_X1   g128(.A1(new_n328), .A2(new_n329), .A3(new_n321), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n324), .A2(KEYINPUT2), .ZN(new_n331));
  XNOR2_X1  g130(.A(G141gat), .B(G148gat), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT77), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n314), .A2(G148gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n312), .A2(G141gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n335), .A2(new_n336), .A3(new_n333), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n330), .B1(new_n334), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n326), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT3), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(new_n227), .A3(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT80), .B(KEYINPUT5), .ZN(new_n345));
  NAND2_X1  g144(.A1(G225gat), .A2(G233gat), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT4), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n317), .A2(new_n318), .B1(new_n324), .B2(new_n323), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n312), .A2(G141gat), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT77), .B1(new_n351), .B2(new_n316), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n352), .A2(new_n337), .A3(new_n331), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n350), .A2(new_n320), .B1(new_n353), .B2(new_n330), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n349), .B1(new_n354), .B2(new_n269), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT82), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n354), .A2(new_n349), .A3(new_n269), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n354), .A2(new_n269), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n359), .A2(new_n356), .A3(KEYINPUT4), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n344), .B(new_n348), .C1(new_n358), .C2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT4), .B1(new_n340), .B2(new_n227), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(new_n357), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n364), .A2(new_n346), .A3(new_n344), .ZN(new_n365));
  INV_X1    g164(.A(new_n345), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n340), .A2(new_n227), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n359), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n366), .B1(new_n368), .B2(new_n347), .ZN(new_n369));
  AND3_X1   g168(.A1(new_n365), .A2(new_n369), .A3(KEYINPUT81), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT81), .B1(new_n365), .B2(new_n369), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n362), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(G1gat), .B(G29gat), .ZN(new_n373));
  INV_X1    g172(.A(G85gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT0), .B(G57gat), .ZN(new_n376));
  XOR2_X1   g175(.A(new_n375), .B(new_n376), .Z(new_n377));
  NAND2_X1  g176(.A1(new_n372), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT6), .ZN(new_n379));
  INV_X1    g178(.A(new_n377), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n380), .B(new_n362), .C1(new_n370), .C2(new_n371), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n378), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G8gat), .B(G36gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n383), .B(G92gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(KEYINPUT74), .B(G64gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n384), .B(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n274), .A2(new_n280), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT29), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(G226gat), .A2(G233gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G211gat), .B(G218gat), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT73), .ZN(new_n393));
  OR2_X1    g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n393), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n396));
  INV_X1    g195(.A(G197gat), .ZN(new_n397));
  INV_X1    g196(.A(G204gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(G197gat), .A2(G204gat), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n396), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n394), .A2(new_n395), .A3(new_n401), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n399), .A2(new_n400), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n393), .B(new_n392), .C1(new_n403), .C2(new_n396), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n390), .B1(new_n274), .B2(new_n280), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n391), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  AOI22_X1  g208(.A1(new_n387), .A2(new_n388), .B1(G226gat), .B2(G233gat), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n405), .B1(new_n410), .B2(new_n407), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT37), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n409), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n412), .B1(new_n409), .B2(new_n411), .ZN(new_n415));
  OAI211_X1 g214(.A(KEYINPUT38), .B(new_n386), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n386), .ZN(new_n417));
  INV_X1    g216(.A(new_n415), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n417), .B1(new_n418), .B2(new_n413), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n409), .A2(new_n411), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n417), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT38), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n416), .B1(new_n419), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n372), .A2(KEYINPUT6), .A3(new_n377), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n382), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n368), .A2(new_n347), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT39), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n344), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n357), .A2(new_n356), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n363), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n430), .B1(new_n432), .B2(new_n360), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n429), .B1(new_n433), .B2(new_n346), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n344), .B1(new_n358), .B2(new_n361), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n435), .A2(new_n428), .A3(new_n347), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n434), .A2(new_n380), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT40), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT30), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n421), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT75), .B1(new_n420), .B2(new_n417), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT75), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n409), .A2(new_n411), .A3(new_n443), .A4(new_n386), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n420), .A2(KEYINPUT30), .A3(new_n417), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n441), .A2(new_n442), .A3(new_n444), .A4(new_n445), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n434), .A2(new_n436), .A3(KEYINPUT40), .A4(new_n380), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n439), .A2(new_n446), .A3(new_n378), .A4(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n405), .B1(new_n388), .B2(new_n343), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n402), .A2(new_n388), .A3(new_n404), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n354), .B1(new_n450), .B2(new_n342), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT83), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(G228gat), .A2(G233gat), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  OAI211_X1 g254(.A(KEYINPUT83), .B(new_n453), .C1(new_n449), .C2(new_n451), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(G78gat), .B(G106gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(KEYINPUT31), .B(G50gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n459), .B(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(G22gat), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT85), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n452), .A2(new_n454), .ZN(new_n466));
  XOR2_X1   g265(.A(KEYINPUT84), .B(G22gat), .Z(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n466), .A2(new_n456), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n468), .B1(new_n466), .B2(new_n456), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n465), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n465), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n463), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n448), .A2(new_n475), .ZN(new_n476));
  OAI22_X1  g275(.A1(new_n309), .A2(new_n310), .B1(new_n426), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n382), .A2(new_n425), .ZN(new_n478));
  INV_X1    g277(.A(new_n446), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n463), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n467), .B1(new_n455), .B2(new_n457), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n473), .B1(new_n482), .B2(new_n469), .ZN(new_n483));
  INV_X1    g282(.A(new_n474), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n480), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT35), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n485), .B1(new_n306), .B2(new_n308), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n446), .B1(new_n382), .B2(new_n425), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT86), .ZN(new_n492));
  INV_X1    g291(.A(new_n305), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n492), .B1(new_n493), .B2(new_n307), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n303), .A2(KEYINPUT86), .A3(new_n305), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(new_n495), .A3(new_n475), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n381), .A2(new_n379), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT81), .ZN(new_n498));
  NOR3_X1   g297(.A1(new_n340), .A2(KEYINPUT4), .A3(new_n227), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n499), .A2(new_n355), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n343), .A2(new_n227), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n342), .B1(new_n326), .B2(new_n339), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n346), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n340), .A2(new_n227), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n326), .A2(new_n339), .B1(new_n226), .B2(new_n219), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n347), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n345), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n498), .B1(new_n504), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n365), .A2(new_n369), .A3(KEYINPUT81), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n380), .B1(new_n511), .B2(new_n362), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n497), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n425), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n488), .B(new_n479), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n496), .A2(new_n515), .ZN(new_n516));
  OAI22_X1  g315(.A1(new_n477), .A2(new_n487), .B1(new_n491), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  XOR2_X1   g317(.A(G43gat), .B(G50gat), .Z(new_n519));
  OR2_X1    g318(.A1(new_n519), .A2(KEYINPUT88), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT15), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n521), .B1(new_n519), .B2(KEYINPUT88), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  OR3_X1    g322(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT90), .B(G36gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(G29gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n519), .A2(new_n521), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n523), .A2(new_n526), .A3(new_n528), .A4(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n526), .A2(KEYINPUT89), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(new_n528), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n526), .A2(KEYINPUT89), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n520), .B(new_n522), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(KEYINPUT91), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT16), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n537), .A2(G1gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(G15gat), .B(G22gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(KEYINPUT92), .ZN(new_n540));
  MUX2_X1   g339(.A(G1gat), .B(new_n538), .S(new_n540), .Z(new_n541));
  INV_X1    g340(.A(G8gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n536), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(KEYINPUT93), .ZN(new_n545));
  NAND2_X1  g344(.A1(G229gat), .A2(G233gat), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT17), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n536), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n543), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n535), .A2(KEYINPUT17), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n545), .A2(KEYINPUT18), .A3(new_n546), .A4(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n544), .A2(KEYINPUT93), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT93), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n554), .B1(new_n536), .B2(new_n543), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n546), .B(new_n551), .C1(new_n553), .C2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT18), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI22_X1  g357(.A1(new_n553), .A2(new_n555), .B1(new_n543), .B2(new_n536), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n546), .B(KEYINPUT13), .Z(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(G113gat), .B(G141gat), .Z(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT87), .B(G197gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(KEYINPUT11), .B(G169gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n566), .B(KEYINPUT12), .Z(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n552), .A2(new_n558), .A3(new_n561), .A4(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  AOI22_X1  g369(.A1(new_n557), .A2(new_n556), .B1(new_n559), .B2(new_n560), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n568), .B1(new_n571), .B2(new_n552), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n518), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT94), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(G162gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT97), .B(G134gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G85gat), .A2(G92gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT7), .ZN(new_n582));
  INV_X1    g381(.A(G99gat), .ZN(new_n583));
  INV_X1    g382(.A(G106gat), .ZN(new_n584));
  OAI21_X1  g383(.A(KEYINPUT8), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n582), .B(new_n585), .C1(G85gat), .C2(G92gat), .ZN(new_n586));
  XOR2_X1   g385(.A(G99gat), .B(G106gat), .Z(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n536), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT98), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n590), .A2(KEYINPUT98), .A3(new_n591), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(G190gat), .B(G218gat), .Z(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n548), .A2(new_n550), .A3(new_n588), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n596), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n598), .B1(new_n596), .B2(new_n599), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n580), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n602), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n604), .A2(new_n600), .A3(new_n579), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G57gat), .B(G64gat), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G71gat), .B(G78gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT21), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n543), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n611), .B(KEYINPUT21), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n614), .B1(new_n543), .B2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G183gat), .B(G211gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT96), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT19), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT20), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n616), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G231gat), .A2(G233gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT95), .ZN(new_n623));
  XNOR2_X1  g422(.A(G127gat), .B(G155gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n621), .B(new_n625), .Z(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(G230gat), .A2(G233gat), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n588), .A2(new_n611), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n588), .A2(new_n611), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT99), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT10), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n629), .A2(new_n633), .A3(new_n630), .ZN(new_n634));
  OR3_X1    g433(.A1(new_n588), .A2(new_n633), .A3(new_n611), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n628), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n632), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G120gat), .B(G148gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(G204gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT100), .B(G176gat), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n640), .B(new_n641), .Z(new_n642));
  OR2_X1    g441(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n632), .A2(new_n642), .A3(new_n637), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n606), .A2(new_n627), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n575), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n478), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(G1gat), .ZN(G1324gat));
  INV_X1    g452(.A(KEYINPUT42), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT101), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(new_n542), .ZN(new_n656));
  AND4_X1   g455(.A1(new_n654), .A2(new_n650), .A3(new_n446), .A4(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n650), .A2(new_n446), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n654), .B1(new_n658), .B2(G8gat), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n650), .A2(new_n446), .A3(new_n656), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n657), .B1(new_n659), .B2(new_n660), .ZN(G1325gat));
  NAND2_X1  g460(.A1(new_n494), .A2(new_n495), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n649), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n663), .A2(G15gat), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n309), .A2(new_n310), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(G15gat), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n649), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(KEYINPUT102), .B1(new_n664), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT102), .ZN(new_n669));
  OAI221_X1 g468(.A(new_n669), .B1(new_n649), .B2(new_n666), .C1(new_n663), .C2(G15gat), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n670), .ZN(G1326gat));
  NOR2_X1   g470(.A1(new_n649), .A2(new_n475), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT43), .B(G22gat), .Z(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(G1327gat));
  NAND2_X1  g473(.A1(new_n306), .A2(new_n308), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n675), .A2(new_n490), .A3(new_n475), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(KEYINPUT35), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n494), .A2(new_n495), .A3(new_n475), .ZN(new_n678));
  AOI211_X1 g477(.A(KEYINPUT35), .B(new_n446), .C1(new_n382), .C2(new_n425), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n424), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n448), .B(new_n475), .C1(new_n478), .C2(new_n682), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n486), .B(new_n683), .C1(new_n309), .C2(new_n310), .ZN(new_n684));
  AOI211_X1 g483(.A(KEYINPUT44), .B(new_n606), .C1(new_n681), .C2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686));
  INV_X1    g485(.A(new_n606), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n686), .B1(new_n517), .B2(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n627), .A2(new_n645), .ZN(new_n690));
  INV_X1    g489(.A(new_n573), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(G29gat), .B1(new_n694), .B2(new_n478), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT45), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n606), .A2(new_n627), .A3(new_n645), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n575), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n478), .A2(G29gat), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n696), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NOR4_X1   g500(.A1(new_n698), .A2(KEYINPUT45), .A3(G29gat), .A4(new_n478), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n695), .B1(new_n701), .B2(new_n702), .ZN(G1328gat));
  NOR2_X1   g502(.A1(new_n479), .A2(new_n527), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT103), .B(KEYINPUT46), .Z(new_n705));
  NAND3_X1  g504(.A1(new_n699), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n527), .B1(new_n694), .B2(new_n479), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n705), .B1(new_n699), .B2(new_n704), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n708), .A2(new_n709), .ZN(G1329gat));
  INV_X1    g509(.A(G43gat), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n711), .B1(new_n698), .B2(new_n662), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n693), .A2(G43gat), .A3(new_n665), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n712), .A2(KEYINPUT47), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(KEYINPUT47), .B1(new_n712), .B2(new_n713), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n714), .A2(new_n715), .ZN(G1330gat));
  INV_X1    g515(.A(new_n688), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n517), .A2(new_n686), .A3(new_n687), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n719), .A2(new_n691), .A3(new_n485), .A4(new_n690), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(G50gat), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n475), .A2(G50gat), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n574), .A2(KEYINPUT94), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n574), .A2(KEYINPUT94), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n697), .B(new_n722), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n721), .A2(new_n725), .A3(KEYINPUT48), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT104), .B(KEYINPUT48), .ZN(new_n727));
  INV_X1    g526(.A(G50gat), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n728), .B1(new_n693), .B2(new_n485), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n727), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n721), .A2(new_n725), .A3(KEYINPUT105), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n731), .A2(new_n732), .A3(KEYINPUT106), .ZN(new_n733));
  AOI21_X1  g532(.A(KEYINPUT106), .B1(new_n731), .B2(new_n732), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n726), .B1(new_n733), .B2(new_n734), .ZN(G1331gat));
  NAND4_X1  g534(.A1(new_n573), .A2(new_n606), .A3(new_n627), .A4(new_n645), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n518), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n651), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(G57gat), .ZN(G1332gat));
  XOR2_X1   g538(.A(new_n737), .B(KEYINPUT107), .Z(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n446), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n742));
  XOR2_X1   g541(.A(KEYINPUT49), .B(G64gat), .Z(new_n743));
  OAI21_X1  g542(.A(new_n742), .B1(new_n741), .B2(new_n743), .ZN(G1333gat));
  NAND2_X1  g543(.A1(new_n740), .A2(new_n665), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n662), .A2(G71gat), .ZN(new_n746));
  AOI22_X1  g545(.A1(new_n745), .A2(G71gat), .B1(new_n737), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g547(.A1(new_n740), .A2(new_n485), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT109), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n740), .A2(new_n751), .A3(new_n485), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(KEYINPUT108), .B(G78gat), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n750), .A2(new_n752), .A3(new_n754), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(G1335gat));
  NOR2_X1   g557(.A1(new_n691), .A2(new_n627), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n759), .A2(new_n517), .A3(new_n687), .ZN(new_n760));
  OR2_X1    g559(.A1(new_n760), .A2(KEYINPUT51), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(KEYINPUT51), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n761), .A2(new_n645), .A3(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(G85gat), .B1(new_n764), .B2(new_n651), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n552), .A2(new_n558), .A3(new_n561), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n567), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n626), .A2(new_n767), .A3(new_n569), .A4(new_n645), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT110), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(new_n685), .B2(new_n688), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT111), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI211_X1 g571(.A(KEYINPUT111), .B(new_n769), .C1(new_n685), .C2(new_n688), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n478), .A2(new_n374), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n765), .B1(new_n774), .B2(new_n775), .ZN(G1336gat));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n479), .A2(G92gat), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n719), .A2(new_n446), .A3(new_n769), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT113), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(G92gat), .B1(new_n779), .B2(new_n780), .ZN(new_n782));
  OAI221_X1 g581(.A(new_n777), .B1(new_n763), .B2(new_n778), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n760), .A2(KEYINPUT112), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n760), .A2(KEYINPUT112), .A3(KEYINPUT51), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n786), .A2(new_n645), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(new_n778), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n446), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n789), .B1(new_n790), .B2(G92gat), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n783), .B1(new_n777), .B2(new_n791), .ZN(G1337gat));
  INV_X1    g591(.A(new_n662), .ZN(new_n793));
  AOI21_X1  g592(.A(G99gat), .B1(new_n764), .B2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n665), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n795), .A2(new_n583), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n794), .B1(new_n774), .B2(new_n796), .ZN(G1338gat));
  NOR2_X1   g596(.A1(new_n475), .A2(G106gat), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT53), .B1(new_n764), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n719), .A2(new_n485), .A3(new_n769), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n800), .A2(KEYINPUT115), .ZN(new_n801));
  OAI21_X1  g600(.A(G106gat), .B1(new_n800), .B2(KEYINPUT115), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n799), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n786), .A2(new_n645), .A3(new_n787), .A4(new_n798), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n475), .B1(new_n772), .B2(new_n773), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n805), .B2(new_n584), .ZN(new_n806));
  AND3_X1   g605(.A1(new_n806), .A2(KEYINPUT114), .A3(KEYINPUT53), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT114), .B1(new_n806), .B2(KEYINPUT53), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n803), .B1(new_n807), .B2(new_n808), .ZN(G1339gat));
  NOR2_X1   g608(.A1(new_n478), .A2(new_n446), .ZN(new_n810));
  INV_X1    g609(.A(new_n628), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n634), .A2(new_n811), .A3(new_n635), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n637), .A2(KEYINPUT54), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n811), .B1(new_n634), .B2(new_n635), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n642), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT55), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n818));
  OR2_X1    g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n813), .A2(KEYINPUT55), .A3(new_n816), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n644), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n817), .A2(new_n818), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n819), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n824), .B1(new_n767), .B2(new_n569), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n559), .A2(new_n560), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n546), .B1(new_n545), .B2(new_n551), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n566), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n828), .A2(new_n569), .A3(new_n645), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT117), .B1(new_n825), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n824), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n832), .B1(new_n570), .B2(new_n572), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n833), .A2(new_n834), .A3(new_n829), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n831), .A2(new_n835), .A3(new_n606), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n828), .A2(new_n569), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n687), .A2(new_n837), .A3(new_n832), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n627), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n647), .A2(new_n691), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n678), .B(new_n810), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(G113gat), .B1(new_n841), .B2(new_n573), .ZN(new_n842));
  OR2_X1    g641(.A1(new_n839), .A2(new_n840), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(new_n489), .A3(new_n810), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n691), .A2(new_n204), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n842), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(KEYINPUT118), .ZN(G1340gat));
  OAI21_X1  g646(.A(G120gat), .B1(new_n841), .B2(new_n646), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n645), .A2(new_n207), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n848), .B1(new_n844), .B2(new_n849), .ZN(G1341gat));
  INV_X1    g649(.A(G127gat), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n841), .A2(new_n851), .A3(new_n626), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n844), .A2(new_n626), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(new_n853), .B2(new_n851), .ZN(G1342gat));
  NAND2_X1  g653(.A1(new_n221), .A2(new_n223), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n687), .A2(new_n855), .ZN(new_n856));
  OR3_X1    g655(.A1(new_n844), .A2(KEYINPUT56), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(G134gat), .B1(new_n841), .B2(new_n606), .ZN(new_n858));
  OAI21_X1  g657(.A(KEYINPUT56), .B1(new_n844), .B2(new_n856), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(G1343gat));
  INV_X1    g659(.A(new_n810), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n665), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n821), .A2(new_n817), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n864), .B1(new_n767), .B2(new_n569), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n606), .B1(new_n865), .B2(new_n830), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n627), .B1(new_n838), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n485), .B1(new_n867), .B2(new_n840), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n863), .B1(new_n868), .B2(KEYINPUT57), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n870), .B(new_n485), .C1(new_n839), .C2(new_n840), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(G141gat), .B1(new_n872), .B2(new_n573), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n485), .B1(new_n839), .B2(new_n840), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n875), .A2(new_n314), .A3(new_n691), .A4(new_n862), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT58), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT58), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n873), .A2(new_n879), .A3(new_n876), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(G1344gat));
  NAND2_X1  g680(.A1(new_n312), .A2(KEYINPUT59), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n875), .A2(new_n862), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n882), .B1(new_n884), .B2(new_n645), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n874), .A2(KEYINPUT57), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n868), .A2(KEYINPUT57), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n888));
  OAI21_X1  g687(.A(KEYINPUT59), .B1(new_n863), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n889), .B1(new_n888), .B2(new_n863), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n886), .A2(new_n645), .A3(new_n887), .A4(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n872), .A2(new_n646), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n891), .B1(new_n892), .B2(KEYINPUT59), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n885), .B1(new_n893), .B2(G148gat), .ZN(G1345gat));
  INV_X1    g693(.A(G155gat), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n872), .A2(new_n895), .A3(new_n626), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n875), .A2(new_n627), .A3(new_n862), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n898));
  OR2_X1    g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(G155gat), .B1(new_n897), .B2(new_n898), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n896), .B1(new_n899), .B2(new_n900), .ZN(G1346gat));
  OR3_X1    g700(.A1(new_n883), .A2(G162gat), .A3(new_n606), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n869), .A2(new_n871), .A3(new_n687), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT121), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(G162gat), .B1(new_n903), .B2(new_n904), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n902), .B1(new_n905), .B2(new_n906), .ZN(G1347gat));
  INV_X1    g706(.A(new_n489), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n478), .A2(new_n446), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n843), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n259), .A3(new_n691), .ZN(new_n912));
  XOR2_X1   g711(.A(new_n909), .B(KEYINPUT122), .Z(new_n913));
  AND2_X1   g712(.A1(new_n913), .A2(new_n678), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n843), .A2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n691), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n912), .B1(new_n918), .B2(new_n259), .ZN(G1348gat));
  AOI21_X1  g718(.A(G176gat), .B1(new_n911), .B2(new_n645), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n646), .A2(new_n260), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n916), .B2(new_n921), .ZN(G1349gat));
  INV_X1    g721(.A(KEYINPUT123), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n923), .A2(KEYINPUT60), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n843), .A2(new_n910), .A3(new_n235), .A4(new_n627), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n914), .B(new_n627), .C1(new_n839), .C2(new_n840), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(G183gat), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n924), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n923), .A2(KEYINPUT60), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n928), .B(new_n929), .ZN(G1350gat));
  NAND4_X1  g729(.A1(new_n843), .A2(new_n910), .A3(new_n228), .A4(new_n687), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT124), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n931), .B(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(G190gat), .B1(new_n915), .B2(new_n606), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n934), .A2(KEYINPUT61), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n934), .A2(KEYINPUT61), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(G1351gat));
  AND2_X1   g736(.A1(new_n913), .A2(new_n795), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n886), .A2(new_n887), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g738(.A(G197gat), .B1(new_n939), .B2(new_n573), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n665), .A2(new_n909), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n941), .B(new_n485), .C1(new_n839), .C2(new_n840), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n691), .A2(new_n397), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(G1352gat));
  NOR3_X1   g743(.A1(new_n942), .A2(G204gat), .A3(new_n646), .ZN(new_n945));
  XNOR2_X1  g744(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n945), .B(new_n946), .ZN(new_n947));
  AND4_X1   g746(.A1(new_n645), .A2(new_n886), .A3(new_n887), .A4(new_n938), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n947), .B1(new_n398), .B2(new_n948), .ZN(G1353gat));
  OR3_X1    g748(.A1(new_n942), .A2(G211gat), .A3(new_n626), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n886), .A2(new_n627), .A3(new_n887), .A4(new_n938), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n951), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n952));
  AOI21_X1  g751(.A(KEYINPUT63), .B1(new_n951), .B2(G211gat), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n950), .B1(new_n952), .B2(new_n953), .ZN(G1354gat));
  INV_X1    g753(.A(KEYINPUT127), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n886), .A2(new_n955), .A3(new_n887), .A4(new_n938), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n956), .A2(G218gat), .A3(new_n687), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n939), .A2(KEYINPUT127), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n942), .A2(new_n606), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT126), .ZN(new_n960));
  OR3_X1    g759(.A1(new_n959), .A2(new_n960), .A3(G218gat), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n960), .B1(new_n959), .B2(G218gat), .ZN(new_n962));
  AOI22_X1  g761(.A1(new_n957), .A2(new_n958), .B1(new_n961), .B2(new_n962), .ZN(G1355gat));
endmodule


