//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0 1 1 0 0 1 1 1 1 0 1 0 1 0 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 0 1 1 1 1 1 1 1 1 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1339, new_n1340;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G20), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT64), .Z(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n210), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n213), .B1(new_n216), .B2(new_n217), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT2), .B(G226), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n230), .B(new_n233), .Z(G358));
  XOR2_X1   g0034(.A(G87), .B(G97), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT65), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G58), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G351));
  INV_X1    g0042(.A(KEYINPUT66), .ZN(new_n243));
  AND2_X1   g0043(.A1(G33), .A2(G41), .ZN(new_n244));
  OAI21_X1  g0044(.A(new_n243), .B1(new_n244), .B2(new_n214), .ZN(new_n245));
  OAI21_X1  g0045(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(G33), .A2(G41), .ZN(new_n248));
  NAND4_X1  g0048(.A1(new_n248), .A2(KEYINPUT66), .A3(G1), .A4(G13), .ZN(new_n249));
  NAND4_X1  g0049(.A1(new_n245), .A2(new_n247), .A3(G274), .A4(new_n249), .ZN(new_n250));
  NAND4_X1  g0050(.A1(new_n245), .A2(G232), .A3(new_n246), .A4(new_n249), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G87), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G223), .A2(G1698), .ZN(new_n255));
  INV_X1    g0055(.A(G226), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n255), .B1(new_n256), .B2(G1698), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT3), .B(G33), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n254), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n215), .A2(new_n248), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n250), .B(new_n251), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(G179), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT80), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n260), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n256), .A2(G1698), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(G223), .B2(G1698), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT3), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n265), .B1(new_n272), .B2(new_n254), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n273), .A2(KEYINPUT80), .A3(new_n250), .A4(new_n251), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n264), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G169), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n262), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g0077(.A(G58), .B(G68), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G20), .A2(G33), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n278), .A2(G20), .B1(G159), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n208), .A2(KEYINPUT7), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n281), .B1(new_n269), .B2(new_n270), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n268), .A2(G33), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n208), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT7), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n282), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI211_X1 g0087(.A(KEYINPUT16), .B(new_n280), .C1(new_n287), .C2(new_n203), .ZN(new_n288));
  NAND3_X1  g0088(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n214), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT16), .ZN(new_n292));
  AOI21_X1  g0092(.A(G20), .B1(new_n269), .B2(new_n270), .ZN(new_n293));
  OAI21_X1  g0093(.A(KEYINPUT76), .B1(new_n293), .B2(KEYINPUT7), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT76), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n295), .B(new_n286), .C1(new_n258), .C2(G20), .ZN(new_n296));
  INV_X1    g0096(.A(new_n281), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT77), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n269), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n268), .A2(KEYINPUT77), .A3(G33), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n299), .A2(new_n270), .A3(new_n300), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n294), .A2(new_n296), .B1(new_n297), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n280), .B1(new_n302), .B2(new_n203), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n291), .B1(new_n292), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT79), .ZN(new_n305));
  XNOR2_X1  g0105(.A(KEYINPUT8), .B(G58), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT8), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G58), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n207), .A2(G20), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n307), .A2(new_n214), .A3(new_n289), .ZN(new_n316));
  OAI211_X1 g0116(.A(KEYINPUT78), .B(new_n309), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n289), .A2(new_n214), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n319), .A2(new_n313), .A3(new_n307), .A4(new_n314), .ZN(new_n320));
  AOI21_X1  g0120(.A(KEYINPUT78), .B1(new_n320), .B2(new_n309), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n305), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n309), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT78), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n325), .A2(KEYINPUT79), .A3(new_n317), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n277), .B(KEYINPUT18), .C1(new_n304), .C2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n280), .ZN(new_n330));
  OAI22_X1  g0130(.A1(new_n293), .A2(KEYINPUT7), .B1(new_n258), .B2(new_n281), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n330), .B1(new_n331), .B2(G68), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n319), .B1(new_n332), .B2(KEYINPUT16), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n301), .A2(new_n297), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n295), .B1(new_n285), .B2(new_n286), .ZN(new_n335));
  NOR3_X1   g0135(.A1(new_n293), .A2(KEYINPUT76), .A3(KEYINPUT7), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n330), .B1(new_n337), .B2(G68), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n333), .B1(new_n338), .B2(KEYINPUT16), .ZN(new_n339));
  INV_X1    g0139(.A(new_n327), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT18), .B1(new_n341), .B2(new_n277), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n329), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(G200), .B1(new_n264), .B2(new_n274), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n261), .A2(G190), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n339), .B(new_n340), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT17), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n303), .A2(new_n292), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n327), .B1(new_n349), .B2(new_n333), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n264), .A2(new_n274), .ZN(new_n351));
  OAI22_X1  g0151(.A1(new_n351), .A2(G200), .B1(G190), .B2(new_n261), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n350), .A2(new_n352), .A3(KEYINPUT17), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n343), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n245), .A2(new_n246), .A3(new_n249), .ZN(new_n356));
  OR2_X1    g0156(.A1(new_n356), .A2(new_n256), .ZN(new_n357));
  INV_X1    g0157(.A(G77), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n260), .B1(new_n358), .B2(new_n271), .ZN(new_n359));
  MUX2_X1   g0159(.A(G222), .B(G223), .S(G1698), .Z(new_n360));
  OAI21_X1  g0160(.A(new_n359), .B1(new_n271), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n357), .A2(new_n361), .A3(new_n250), .ZN(new_n362));
  XOR2_X1   g0162(.A(KEYINPUT68), .B(G200), .Z(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n208), .A2(G33), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n313), .A2(new_n366), .B1(G150), .B2(new_n279), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n204), .A2(G20), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n319), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n314), .A2(G50), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n316), .A2(new_n370), .B1(G50), .B2(new_n307), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT9), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n357), .A2(new_n361), .A3(G190), .A4(new_n250), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT9), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n369), .B2(new_n371), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n364), .A2(new_n373), .A3(new_n374), .A4(new_n376), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n377), .A2(KEYINPUT10), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n377), .A2(KEYINPUT10), .ZN(new_n379));
  OR2_X1    g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n258), .A2(G238), .A3(G1698), .ZN(new_n381));
  INV_X1    g0181(.A(G1698), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n258), .A2(G232), .A3(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(G107), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n381), .B(new_n383), .C1(new_n384), .C2(new_n258), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n265), .ZN(new_n386));
  INV_X1    g0186(.A(G244), .ZN(new_n387));
  OR2_X1    g0187(.A1(new_n356), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(new_n250), .A3(new_n388), .ZN(new_n389));
  OR2_X1    g0189(.A1(new_n389), .A2(G179), .ZN(new_n390));
  INV_X1    g0190(.A(new_n279), .ZN(new_n391));
  OAI22_X1  g0191(.A1(new_n306), .A2(new_n391), .B1(new_n208), .B2(new_n358), .ZN(new_n392));
  XNOR2_X1  g0192(.A(KEYINPUT15), .B(G87), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n393), .A2(new_n365), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n290), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  XNOR2_X1  g0195(.A(new_n395), .B(KEYINPUT67), .ZN(new_n396));
  INV_X1    g0196(.A(new_n316), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n358), .B1(new_n207), .B2(G20), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n397), .A2(new_n398), .B1(new_n358), .B2(new_n308), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n389), .A2(new_n276), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n390), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n389), .A2(new_n363), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n386), .A2(G190), .A3(new_n250), .A4(new_n388), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n403), .A2(new_n404), .A3(new_n396), .A4(new_n399), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT69), .ZN(new_n408));
  OR2_X1    g0208(.A1(new_n362), .A2(G179), .ZN(new_n409));
  INV_X1    g0209(.A(new_n372), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n362), .A2(new_n276), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n380), .A2(new_n407), .A3(new_n408), .A4(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n412), .B1(new_n378), .B2(new_n379), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT69), .B1(new_n414), .B2(new_n406), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n355), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n366), .A2(G77), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n279), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n319), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  XNOR2_X1  g0219(.A(new_n419), .B(KEYINPUT11), .ZN(new_n420));
  OR2_X1    g0220(.A1(new_n420), .A2(KEYINPUT74), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(KEYINPUT74), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT12), .B1(new_n307), .B2(G68), .ZN(new_n423));
  OR3_X1    g0223(.A1(new_n307), .A2(KEYINPUT12), .A3(G68), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n203), .B1(new_n207), .B2(G20), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n423), .A2(new_n424), .B1(new_n397), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n421), .A2(new_n422), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n256), .A2(G1698), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n429), .A2(new_n269), .A3(new_n270), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT70), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(G33), .A2(G97), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n269), .A2(new_n270), .A3(G232), .A4(G1698), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n429), .A2(new_n269), .A3(new_n270), .A4(KEYINPUT70), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n432), .A2(new_n433), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(KEYINPUT71), .B1(new_n436), .B2(new_n265), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n436), .A2(KEYINPUT71), .A3(new_n265), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT73), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT13), .ZN(new_n442));
  INV_X1    g0242(.A(G238), .ZN(new_n443));
  OR2_X1    g0243(.A1(new_n356), .A2(new_n443), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n444), .A2(new_n250), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n440), .A2(new_n441), .A3(new_n442), .A4(new_n445), .ZN(new_n446));
  AND3_X1   g0246(.A1(new_n436), .A2(KEYINPUT71), .A3(new_n265), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n445), .B(new_n442), .C1(new_n447), .C2(new_n437), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT73), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n445), .B1(new_n447), .B2(new_n437), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT13), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G190), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n428), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n452), .A2(KEYINPUT72), .A3(new_n448), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT72), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n451), .A2(new_n456), .A3(KEYINPUT13), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n454), .B1(G200), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n455), .A2(G169), .A3(new_n457), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT14), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT14), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n455), .A2(new_n462), .A3(G169), .A4(new_n457), .ZN(new_n463));
  INV_X1    g0263(.A(G179), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n464), .B1(new_n451), .B2(KEYINPUT13), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n465), .A2(new_n446), .A3(new_n449), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT75), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n465), .A2(new_n446), .A3(new_n449), .A4(KEYINPUT75), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n461), .A2(new_n463), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n459), .B1(new_n470), .B2(new_n427), .ZN(new_n471));
  AND3_X1   g0271(.A1(new_n416), .A2(KEYINPUT81), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(KEYINPUT81), .B1(new_n416), .B2(new_n471), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(G257), .A2(G1698), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n382), .A2(G264), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n258), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n477), .B(new_n265), .C1(G303), .C2(new_n258), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n207), .A2(G45), .ZN(new_n479));
  NOR2_X1   g0279(.A1(KEYINPUT5), .A2(G41), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(KEYINPUT5), .A2(G41), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n479), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n483), .A2(G274), .A3(new_n245), .A4(new_n249), .ZN(new_n484));
  INV_X1    g0284(.A(new_n482), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n207), .B(G45), .C1(new_n485), .C2(new_n480), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n486), .A2(new_n245), .A3(G270), .A4(new_n249), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n478), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G169), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT21), .ZN(new_n490));
  OAI22_X1  g0290(.A1(new_n489), .A2(new_n490), .B1(new_n464), .B2(new_n488), .ZN(new_n491));
  NAND2_X1  g0291(.A1(G33), .A2(G283), .ZN(new_n492));
  INV_X1    g0292(.A(G97), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n492), .B(new_n208), .C1(G33), .C2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(G116), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G20), .ZN(new_n496));
  AND3_X1   g0296(.A1(new_n290), .A2(KEYINPUT84), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(KEYINPUT84), .B1(new_n290), .B2(new_n496), .ZN(new_n498));
  OAI211_X1 g0298(.A(KEYINPUT20), .B(new_n494), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT85), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n290), .A2(new_n496), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT84), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n290), .A2(KEYINPUT84), .A3(new_n496), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT85), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT20), .A4(new_n494), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n494), .B1(new_n497), .B2(new_n498), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT20), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n500), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n307), .A2(new_n495), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n316), .B1(new_n207), .B2(G33), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n513), .B2(new_n495), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n491), .A2(new_n515), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n511), .A2(new_n514), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n488), .A2(G200), .ZN(new_n518));
  INV_X1    g0318(.A(G190), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n517), .B(new_n518), .C1(new_n519), .C2(new_n488), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT86), .ZN(new_n521));
  INV_X1    g0321(.A(new_n489), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n515), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n490), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n489), .B1(new_n511), .B2(new_n514), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n525), .A2(new_n521), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n516), .B(new_n520), .C1(new_n524), .C2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n443), .A2(new_n382), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n387), .A2(G1698), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n258), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G116), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n260), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(G45), .ZN(new_n533));
  OR3_X1    g0333(.A1(new_n533), .A2(G1), .A3(G274), .ZN(new_n534));
  INV_X1    g0334(.A(G250), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n479), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n245), .A2(new_n534), .A3(new_n249), .A4(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n363), .B1(new_n532), .B2(new_n538), .ZN(new_n539));
  AND2_X1   g0339(.A1(new_n528), .A2(new_n529), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n540), .A2(new_n258), .B1(G33), .B2(G116), .ZN(new_n541));
  OAI211_X1 g0341(.A(G190), .B(new_n537), .C1(new_n541), .C2(new_n260), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT19), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n208), .B1(new_n433), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n253), .A2(new_n493), .A3(new_n384), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n269), .A2(new_n270), .A3(new_n208), .A4(G68), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n543), .B1(new_n365), .B2(new_n493), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n549), .A2(new_n290), .B1(new_n308), .B2(new_n393), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n513), .A2(G87), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n539), .A2(new_n542), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n549), .A2(new_n290), .ZN(new_n553));
  INV_X1    g0353(.A(new_n393), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n397), .B(new_n554), .C1(G1), .C2(new_n252), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n393), .A2(new_n308), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n553), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n276), .B1(new_n532), .B2(new_n538), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n464), .B(new_n537), .C1(new_n541), .C2(new_n260), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n552), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT25), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(new_n307), .B2(G107), .ZN(new_n563));
  NOR3_X1   g0363(.A1(new_n307), .A2(new_n562), .A3(G107), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n513), .A2(G107), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n269), .A2(new_n270), .A3(new_n208), .A4(G87), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT22), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT22), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n258), .A2(new_n570), .A3(new_n208), .A4(G87), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT23), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n208), .B2(G107), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n384), .A2(KEYINPUT23), .A3(G20), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT87), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n531), .B2(G20), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n208), .A2(KEYINPUT87), .A3(G33), .A4(G116), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n576), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n572), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT24), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT24), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n572), .A2(new_n583), .A3(new_n580), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n567), .B1(new_n585), .B2(new_n290), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n486), .A2(new_n245), .A3(G264), .A4(new_n249), .ZN(new_n587));
  MUX2_X1   g0387(.A(G250), .B(G257), .S(G1698), .Z(new_n588));
  AOI22_X1  g0388(.A1(new_n588), .A2(new_n258), .B1(G33), .B2(G294), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n484), .B(new_n587), .C1(new_n589), .C2(new_n260), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n590), .A2(new_n519), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(G200), .B2(new_n590), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n561), .B1(new_n586), .B2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n486), .A2(new_n245), .A3(G257), .A4(new_n249), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n484), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n269), .A2(new_n270), .A3(G250), .A4(G1698), .ZN(new_n596));
  AND2_X1   g0396(.A1(new_n596), .A2(new_n492), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n387), .A2(G1698), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n258), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT4), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n598), .A2(new_n269), .A3(new_n270), .A4(KEYINPUT4), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT82), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT82), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n258), .A2(new_n604), .A3(KEYINPUT4), .A4(new_n598), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n597), .A2(new_n601), .A3(new_n603), .A4(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n595), .B1(new_n606), .B2(new_n265), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(G190), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n307), .A2(G97), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n609), .B1(new_n513), .B2(G97), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  XNOR2_X1  g0411(.A(G97), .B(G107), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT6), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n613), .A2(new_n493), .A3(G107), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n617), .A2(G20), .B1(G77), .B2(new_n279), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n618), .B1(new_n302), .B2(new_n384), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n611), .B1(new_n619), .B2(new_n290), .ZN(new_n620));
  OAI21_X1  g0420(.A(G200), .B1(new_n607), .B2(KEYINPUT83), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n606), .A2(new_n265), .ZN(new_n622));
  INV_X1    g0422(.A(new_n595), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n622), .A2(KEYINPUT83), .A3(new_n623), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n608), .B(new_n620), .C1(new_n621), .C2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n584), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n583), .B1(new_n572), .B2(new_n580), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n290), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n566), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n590), .A2(G179), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n630), .B1(new_n276), .B2(new_n590), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n615), .B1(new_n613), .B2(new_n612), .ZN(new_n633));
  OAI22_X1  g0433(.A1(new_n633), .A2(new_n208), .B1(new_n358), .B2(new_n391), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n634), .B1(new_n337), .B2(G107), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n610), .B1(new_n635), .B2(new_n319), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n622), .A2(new_n623), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n276), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n607), .A2(new_n464), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n593), .A2(new_n625), .A3(new_n632), .A4(new_n640), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n474), .A2(new_n527), .A3(new_n641), .ZN(G372));
  INV_X1    g0442(.A(new_n412), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT88), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n644), .B1(new_n329), .B2(new_n342), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n277), .B1(new_n304), .B2(new_n327), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT18), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n648), .A2(KEYINPUT88), .A3(new_n328), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n459), .ZN(new_n651));
  INV_X1    g0451(.A(new_n402), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n651), .A2(new_n652), .B1(new_n470), .B2(new_n427), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n650), .B1(new_n653), .B2(new_n354), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n643), .B1(new_n654), .B2(new_n380), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n629), .A2(new_n631), .B1(new_n491), .B2(new_n515), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n656), .B1(new_n524), .B2(new_n526), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n625), .A2(new_n640), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(new_n658), .A3(new_n593), .ZN(new_n659));
  INV_X1    g0459(.A(new_n560), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n640), .B2(new_n561), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n638), .A2(new_n639), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n552), .A2(new_n560), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n663), .A2(KEYINPUT26), .A3(new_n664), .A4(new_n636), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n660), .B1(new_n662), .B2(new_n665), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n659), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n655), .B1(new_n474), .B2(new_n667), .ZN(G369));
  INV_X1    g0468(.A(new_n526), .ZN(new_n669));
  AOI21_X1  g0469(.A(KEYINPUT21), .B1(new_n525), .B2(new_n521), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n669), .A2(new_n670), .B1(new_n491), .B2(new_n515), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n517), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n672), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n527), .B2(new_n680), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n682), .A2(G330), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n586), .A2(new_n592), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n586), .A2(new_n679), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n632), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n632), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n679), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n671), .A2(new_n678), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n691), .A2(new_n689), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n692), .B1(new_n687), .B2(new_n679), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n690), .A2(new_n693), .ZN(G399));
  INV_X1    g0494(.A(new_n211), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G41), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n545), .A2(G116), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G1), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n217), .B2(new_n697), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n678), .B1(new_n659), .B2(new_n666), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT29), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n593), .A2(new_n625), .A3(new_n640), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT89), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n705), .B1(new_n657), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n706), .B2(new_n657), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n678), .B1(new_n708), .B2(new_n666), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n704), .B1(new_n709), .B2(new_n703), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n527), .A2(new_n641), .A3(new_n678), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n488), .A2(new_n464), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n537), .B1(new_n541), .B2(new_n260), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n587), .B1(new_n589), .B2(new_n260), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n712), .A2(new_n607), .A3(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT30), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n712), .A2(new_n715), .A3(new_n607), .A4(KEYINPUT30), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n713), .A2(new_n464), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n637), .A2(new_n488), .A3(new_n720), .A4(new_n590), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n718), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n678), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT31), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n722), .A2(KEYINPUT31), .A3(new_n678), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n711), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(G330), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n710), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n701), .B1(new_n732), .B2(G1), .ZN(G364));
  NOR2_X1   g0533(.A1(new_n682), .A2(G330), .ZN(new_n734));
  INV_X1    g0534(.A(G13), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(G20), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n207), .B1(new_n736), .B2(G45), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n697), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n683), .A2(new_n734), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G13), .A2(G33), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G20), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n682), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n214), .B1(G20), .B2(new_n276), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n208), .A2(new_n464), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(G200), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n749), .A2(new_n750), .A3(G190), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(KEYINPUT91), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n752), .A2(KEYINPUT91), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  XNOR2_X1  g0557(.A(KEYINPUT33), .B(G317), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n363), .A2(G20), .A3(new_n464), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n519), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n757), .A2(new_n758), .B1(G303), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n759), .A2(G190), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G283), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G179), .A2(G200), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n208), .B1(new_n764), .B2(G190), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n765), .A2(KEYINPUT92), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(KEYINPUT92), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G294), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n749), .A2(G190), .A3(G200), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n258), .B1(new_n771), .B2(G311), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n764), .A2(G20), .A3(new_n519), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G329), .ZN(new_n775));
  INV_X1    g0575(.A(G322), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n748), .A2(G190), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(G200), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  OAI211_X1 g0579(.A(new_n772), .B(new_n775), .C1(new_n776), .C2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n777), .A2(new_n750), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT93), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n780), .B1(G326), .B2(new_n783), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n761), .A2(new_n763), .A3(new_n770), .A4(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n762), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n384), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(new_n757), .B2(G68), .ZN(new_n788));
  INV_X1    g0588(.A(new_n781), .ZN(new_n789));
  INV_X1    g0589(.A(new_n771), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n258), .B1(new_n789), .B2(new_n201), .C1(new_n358), .C2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(G87), .B2(new_n760), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n769), .A2(G97), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n774), .A2(G159), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT32), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n795), .B1(G58), .B2(new_n778), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n788), .A2(new_n792), .A3(new_n793), .A4(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n747), .B1(new_n785), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n743), .A2(new_n746), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n695), .A2(new_n258), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(G45), .B2(new_n217), .ZN(new_n801));
  INV_X1    g0601(.A(new_n241), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n801), .B1(G45), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n695), .A2(new_n271), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(G355), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(G116), .B2(new_n211), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n803), .B1(KEYINPUT90), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(KEYINPUT90), .B2(new_n806), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n738), .B(new_n798), .C1(new_n799), .C2(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n740), .B1(new_n745), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(G396));
  NAND2_X1  g0611(.A1(new_n652), .A2(new_n679), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n400), .A2(new_n678), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n405), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n402), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(KEYINPUT95), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT95), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n812), .A2(new_n815), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NOR3_X1   g0620(.A1(new_n702), .A2(new_n820), .A3(KEYINPUT96), .ZN(new_n821));
  INV_X1    g0621(.A(new_n816), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n821), .B1(new_n702), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(KEYINPUT96), .B1(new_n702), .B2(new_n820), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n730), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT97), .Z(new_n828));
  AOI21_X1  g0628(.A(new_n739), .B1(new_n825), .B2(new_n826), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(G283), .ZN(new_n831));
  INV_X1    g0631(.A(new_n760), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n756), .A2(new_n831), .B1(new_n384), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(G87), .B2(new_n762), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n271), .B1(new_n790), .B2(new_n495), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(G311), .B2(new_n774), .ZN(new_n836));
  AOI22_X1  g0636(.A1(G294), .A2(new_n778), .B1(new_n781), .B2(G303), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n834), .A2(new_n793), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT94), .Z(new_n839));
  AOI22_X1  g0639(.A1(new_n771), .A2(G159), .B1(new_n781), .B2(G137), .ZN(new_n840));
  INV_X1    g0640(.A(G143), .ZN(new_n841));
  INV_X1    g0641(.A(G150), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n840), .B1(new_n841), .B2(new_n779), .C1(new_n756), .C2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT34), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n769), .A2(G58), .ZN(new_n846));
  INV_X1    g0646(.A(G132), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n258), .B1(new_n773), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n786), .A2(new_n203), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n848), .B(new_n849), .C1(G50), .C2(new_n760), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n845), .A2(new_n846), .A3(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n843), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n851), .B1(KEYINPUT34), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n746), .B1(new_n839), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n746), .A2(new_n741), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n738), .B1(new_n358), .B2(new_n855), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n854), .B(new_n856), .C1(new_n742), .C2(new_n822), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n830), .A2(new_n857), .ZN(G384));
  AOI211_X1 g0658(.A(new_n495), .B(new_n216), .C1(new_n617), .C2(KEYINPUT35), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(KEYINPUT35), .B2(new_n617), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT36), .ZN(new_n861));
  OAI21_X1  g0661(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n862), .A2(new_n217), .B1(G50), .B2(new_n203), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n863), .A2(G1), .A3(new_n735), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n865), .B(KEYINPUT98), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n710), .B1(new_n472), .B2(new_n473), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n655), .ZN(new_n868));
  XOR2_X1   g0668(.A(new_n868), .B(KEYINPUT103), .Z(new_n869));
  INV_X1    g0669(.A(KEYINPUT38), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n318), .A2(new_n321), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n331), .A2(G68), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT16), .B1(new_n872), .B2(new_n280), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n871), .B1(new_n291), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n676), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(KEYINPUT37), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n350), .A2(new_n352), .B1(new_n277), .B2(new_n874), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n877), .B1(new_n878), .B2(KEYINPUT101), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n275), .A2(new_n276), .ZN(new_n880));
  INV_X1    g0680(.A(new_n262), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n874), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT101), .B1(new_n346), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT37), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n875), .B1(new_n304), .B2(new_n327), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n346), .A2(new_n646), .A3(new_n886), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n879), .A2(new_n884), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n344), .A2(new_n345), .ZN(new_n889));
  NOR3_X1   g0689(.A1(new_n341), .A2(new_n347), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT17), .B1(new_n350), .B2(new_n352), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n648), .A2(new_n328), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n876), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n888), .B1(new_n894), .B2(KEYINPUT100), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT100), .ZN(new_n896));
  AOI211_X1 g0696(.A(new_n896), .B(new_n876), .C1(new_n892), .C2(new_n893), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n870), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n887), .A2(new_n885), .ZN(new_n899));
  OAI211_X1 g0699(.A(KEYINPUT101), .B(new_n882), .C1(new_n341), .C2(new_n889), .ZN(new_n900));
  INV_X1    g0700(.A(new_n877), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n899), .B1(new_n902), .B2(new_n883), .ZN(new_n903));
  INV_X1    g0703(.A(new_n876), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n343), .B2(new_n354), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n903), .B1(new_n905), .B2(new_n896), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n894), .A2(KEYINPUT100), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n906), .A2(KEYINPUT38), .A3(new_n907), .ZN(new_n908));
  AND3_X1   g0708(.A1(new_n898), .A2(KEYINPUT39), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n645), .A2(new_n892), .A3(new_n649), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT102), .ZN(new_n911));
  INV_X1    g0711(.A(new_n886), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n911), .B1(new_n910), .B2(new_n912), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n346), .A2(new_n886), .A3(new_n644), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT37), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n887), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n346), .A2(new_n886), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n919), .A2(KEYINPUT88), .A3(KEYINPUT37), .A4(new_n646), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n914), .A2(new_n915), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n908), .B1(new_n922), .B2(KEYINPUT38), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT39), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n909), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n468), .A2(new_n463), .A3(new_n469), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n460), .A2(KEYINPUT14), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n427), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n928), .A2(new_n678), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n925), .A2(new_n929), .ZN(new_n930));
  AOI211_X1 g0730(.A(new_n678), .B(new_n816), .C1(new_n659), .C2(new_n666), .ZN(new_n931));
  INV_X1    g0731(.A(new_n812), .ZN(new_n932));
  OAI21_X1  g0732(.A(KEYINPUT99), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n702), .A2(new_n822), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT99), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n934), .A2(new_n935), .A3(new_n812), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n427), .A2(new_n678), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n928), .A2(new_n651), .A3(new_n938), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n427), .B(new_n678), .C1(new_n470), .C2(new_n459), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n895), .A2(new_n870), .A3(new_n897), .ZN(new_n943));
  AOI21_X1  g0743(.A(KEYINPUT38), .B1(new_n906), .B2(new_n907), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n650), .A2(new_n875), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n930), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n869), .B(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT40), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n822), .B1(new_n711), .B2(new_n727), .ZN(new_n952));
  AOI211_X1 g0752(.A(new_n951), .B(new_n952), .C1(new_n939), .C2(new_n940), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n952), .B1(new_n939), .B2(new_n940), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n943), .B2(new_n944), .ZN(new_n955));
  XNOR2_X1  g0755(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n923), .A2(new_n953), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n474), .A2(new_n728), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(new_n959), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n960), .A2(G330), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n950), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n207), .B2(new_n736), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n950), .A2(new_n962), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n866), .B1(new_n964), .B2(new_n965), .ZN(G367));
  NAND2_X1  g0766(.A1(new_n550), .A2(new_n551), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n678), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n664), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n560), .B2(new_n968), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT106), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n658), .B1(new_n620), .B2(new_n679), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n640), .B2(new_n679), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n692), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(KEYINPUT42), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n974), .B(KEYINPUT105), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n977), .A2(new_n687), .B1(new_n636), .B2(new_n663), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n976), .B1(new_n978), .B2(new_n678), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n975), .A2(KEYINPUT42), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n972), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n981), .B(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n690), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n977), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n983), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n983), .A2(new_n986), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n696), .B(KEYINPUT41), .Z(new_n989));
  NAND2_X1  g0789(.A1(new_n693), .A2(new_n974), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT45), .Z(new_n991));
  NOR2_X1   g0791(.A1(new_n693), .A2(new_n974), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT44), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n984), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n691), .B(new_n689), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n683), .B(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n732), .A2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n991), .A2(new_n690), .A3(new_n993), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n995), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n989), .B1(new_n1001), .B2(new_n732), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n737), .B(KEYINPUT107), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n987), .B(new_n988), .C1(new_n1002), .C2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n800), .A2(new_n233), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n743), .B(new_n746), .C1(new_n695), .C2(new_n554), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n738), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n757), .A2(G159), .B1(G77), .B2(new_n762), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n768), .A2(new_n203), .ZN(new_n1010));
  INV_X1    g0810(.A(G137), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n258), .B1(new_n773), .B2(new_n1011), .C1(new_n790), .C2(new_n201), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1010), .B(new_n1012), .C1(G150), .C2(new_n778), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n760), .A2(G58), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n783), .A2(G143), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1009), .A2(new_n1013), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n786), .A2(new_n493), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n258), .B1(new_n774), .B2(G317), .ZN(new_n1018));
  INV_X1    g0818(.A(G303), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1018), .B1(new_n779), .B2(new_n1019), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n1017), .B(new_n1020), .C1(new_n757), .C2(G294), .ZN(new_n1021));
  AOI21_X1  g0821(.A(KEYINPUT109), .B1(new_n760), .B2(G116), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT46), .ZN(new_n1023));
  INV_X1    g0823(.A(G311), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1021), .B(new_n1023), .C1(new_n1024), .C2(new_n782), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n768), .A2(new_n384), .B1(new_n790), .B2(new_n831), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT108), .Z(new_n1027));
  OAI21_X1  g0827(.A(new_n1016), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT47), .Z(new_n1029));
  OAI221_X1 g0829(.A(new_n1008), .B1(new_n744), .B2(new_n970), .C1(new_n1029), .C2(new_n747), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1005), .A2(new_n1030), .ZN(G387));
  NOR2_X1   g0831(.A1(new_n689), .A2(new_n744), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n698), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n804), .A2(new_n1033), .B1(new_n384), .B2(new_n695), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n230), .A2(new_n533), .ZN(new_n1035));
  AOI21_X1  g0835(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1036));
  AND3_X1   g0836(.A1(new_n313), .A2(KEYINPUT50), .A3(new_n201), .ZN(new_n1037));
  AOI21_X1  g0837(.A(KEYINPUT50), .B1(new_n313), .B2(new_n201), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n698), .B(new_n1036), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n800), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1034), .B1(new_n1035), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n799), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n739), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n757), .A2(new_n313), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n258), .B1(new_n773), .B2(new_n842), .ZN(new_n1045));
  INV_X1    g0845(.A(G159), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n201), .A2(new_n779), .B1(new_n789), .B2(new_n1046), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n1045), .B(new_n1047), .C1(G68), .C2(new_n771), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1017), .B1(G77), .B2(new_n760), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n769), .A2(new_n554), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1044), .A2(new_n1048), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n258), .B1(new_n774), .B2(G326), .ZN(new_n1052));
  INV_X1    g0852(.A(G294), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n832), .A2(new_n1053), .B1(new_n831), .B2(new_n768), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G303), .A2(new_n771), .B1(new_n778), .B2(G317), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1055), .B1(new_n776), .B2(new_n782), .C1(new_n756), .C2(new_n1024), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT48), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1054), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n1057), .B2(new_n1056), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT49), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1052), .B1(new_n495), .B2(new_n786), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1051), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1032), .B(new_n1043), .C1(new_n1063), .C2(new_n746), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n997), .B2(new_n1004), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n998), .A2(new_n696), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n732), .A2(new_n997), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1065), .B1(new_n1066), .B2(new_n1067), .ZN(G393));
  NAND3_X1  g0868(.A1(new_n995), .A2(new_n1000), .A3(new_n1004), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n238), .A2(new_n800), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n799), .B1(new_n493), .B2(new_n211), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n739), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n757), .A2(G50), .B1(G68), .B2(new_n760), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n258), .B1(new_n773), .B2(new_n841), .C1(new_n790), .C2(new_n306), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(G87), .B2(new_n762), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n842), .A2(new_n789), .B1(new_n779), .B2(new_n1046), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT51), .ZN(new_n1077));
  OR2_X1    g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1076), .A2(new_n1077), .B1(G77), .B2(new_n769), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1073), .A2(new_n1075), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n757), .A2(G303), .B1(G116), .B2(new_n769), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT110), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n271), .B1(new_n773), .B2(new_n776), .C1(new_n790), .C2(new_n1053), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n1084), .B(new_n787), .C1(G283), .C2(new_n760), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G311), .A2(new_n778), .B1(new_n781), .B2(G317), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT52), .Z(new_n1087));
  NAND3_X1  g0887(.A1(new_n1083), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1080), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT111), .Z(new_n1091));
  AOI21_X1  g0891(.A(new_n1072), .B1(new_n1091), .B2(new_n746), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n977), .B2(new_n744), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1069), .A2(new_n1093), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n1001), .A2(new_n696), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n995), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1000), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n998), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1094), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(G390));
  NOR2_X1   g0900(.A1(new_n952), .A2(new_n729), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n941), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n929), .B1(new_n937), .B2(new_n941), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n910), .A2(new_n912), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n921), .B1(new_n1105), .B2(KEYINPUT102), .ZN(new_n1106));
  AOI21_X1  g0906(.A(KEYINPUT38), .B1(new_n1106), .B2(new_n913), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n924), .B1(new_n1107), .B2(new_n943), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n945), .A2(KEYINPUT39), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1104), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n708), .A2(new_n666), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1111), .A2(new_n679), .A3(new_n815), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n812), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n941), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n929), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n923), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1103), .B1(new_n1110), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n923), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1102), .B(new_n1118), .C1(new_n925), .C2(new_n1104), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1117), .A2(new_n1119), .A3(new_n1004), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT113), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n730), .B1(new_n472), .B2(new_n473), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n867), .A2(new_n655), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n932), .B1(new_n709), .B2(new_n815), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n820), .B(G330), .C1(new_n711), .C2(new_n727), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1126), .A2(new_n939), .A3(new_n940), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1102), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(KEYINPUT112), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT112), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1102), .A2(new_n1125), .A3(new_n1130), .A4(new_n1127), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n941), .A2(new_n1101), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n937), .B1(new_n1103), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1124), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1122), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1117), .A2(new_n1135), .A3(new_n1119), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1137), .A2(new_n696), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n855), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n739), .B1(new_n313), .B2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT114), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n757), .A2(G107), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n271), .B1(new_n773), .B2(new_n1053), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n495), .A2(new_n779), .B1(new_n789), .B2(new_n831), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1144), .B(new_n1145), .C1(G97), .C2(new_n771), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n769), .A2(G77), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n849), .B1(G87), .B2(new_n760), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1143), .A2(new_n1146), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(G125), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT54), .B(G143), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n258), .B1(new_n773), .B2(new_n1150), .C1(new_n790), .C2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(new_n757), .B2(G137), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n1153), .B1(new_n201), .B2(new_n786), .C1(new_n1046), .C2(new_n768), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n760), .A2(G150), .ZN(new_n1155));
  XOR2_X1   g0955(.A(new_n1155), .B(KEYINPUT53), .Z(new_n1156));
  AOI22_X1  g0956(.A1(G128), .A2(new_n781), .B1(new_n778), .B2(G132), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT115), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1149), .B1(new_n1154), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1142), .B1(new_n1160), .B2(new_n746), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n925), .B2(new_n742), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1121), .A2(new_n1139), .A3(new_n1162), .ZN(G378));
  INV_X1    g0963(.A(KEYINPUT118), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n955), .A2(new_n956), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n953), .B1(new_n1107), .B2(new_n943), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1165), .A2(new_n1166), .A3(G330), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(KEYINPUT117), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT117), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1165), .A2(new_n1166), .A3(new_n1169), .A4(G330), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n372), .A2(new_n676), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n414), .B(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1172), .B(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1168), .A2(new_n1170), .A3(new_n1174), .ZN(new_n1175));
  AND2_X1   g0975(.A1(new_n930), .A2(new_n948), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1174), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1167), .A2(KEYINPUT117), .A3(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1175), .A2(new_n1176), .A3(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1176), .B1(new_n1178), .B2(new_n1175), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1164), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1169), .B1(new_n957), .B2(G330), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1170), .A2(new_n1174), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1178), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n949), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1187), .A2(KEYINPUT118), .A3(new_n1179), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1182), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1174), .A2(new_n741), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n739), .B1(G50), .B2(new_n1140), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n832), .A2(new_n1151), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n757), .B2(G132), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n790), .A2(new_n1011), .B1(new_n789), .B2(new_n1150), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G128), .B2(new_n778), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1193), .B(new_n1195), .C1(new_n842), .C2(new_n768), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(KEYINPUT59), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n762), .A2(G159), .ZN(new_n1198));
  AOI211_X1 g0998(.A(G33), .B(G41), .C1(new_n774), .C2(G124), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1196), .A2(KEYINPUT59), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n762), .A2(G58), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n258), .A2(G41), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G283), .B2(new_n774), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1202), .B(new_n1204), .C1(new_n832), .C2(new_n358), .ZN(new_n1205));
  XOR2_X1   g1005(.A(new_n1205), .B(KEYINPUT116), .Z(new_n1206));
  AOI22_X1  g1006(.A1(new_n554), .A2(new_n771), .B1(new_n778), .B2(G107), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n495), .B2(new_n789), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1010), .B(new_n1208), .C1(new_n757), .C2(G97), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1206), .A2(new_n1209), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1200), .A2(new_n1201), .B1(KEYINPUT58), .B2(new_n1210), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1203), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(KEYINPUT58), .C2(new_n1210), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1191), .B1(new_n1213), .B2(new_n746), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n1189), .A2(new_n1004), .B1(new_n1190), .B2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1124), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1138), .A2(new_n1216), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1187), .A2(new_n1217), .A3(KEYINPUT57), .A4(new_n1179), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n696), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(KEYINPUT119), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT119), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1218), .A2(new_n1221), .A3(new_n696), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1220), .A2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(KEYINPUT57), .B1(new_n1189), .B2(new_n1217), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1215), .B1(new_n1223), .B2(new_n1224), .ZN(G375));
  INV_X1    g1025(.A(new_n989), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1132), .A2(new_n1124), .A3(new_n1134), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1136), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1003), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n939), .A2(new_n741), .A3(new_n940), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n739), .B1(G68), .B2(new_n1140), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1202), .B1(new_n1046), .B2(new_n832), .C1(new_n756), .C2(new_n1151), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n258), .B1(new_n790), .B2(new_n842), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(G128), .B2(new_n774), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(G132), .A2(new_n781), .B1(new_n778), .B2(G137), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1234), .B(new_n1235), .C1(new_n201), .C2(new_n768), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(G77), .A2(new_n762), .B1(new_n760), .B2(G97), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n756), .B2(new_n495), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n271), .B1(new_n790), .B2(new_n384), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(G303), .B2(new_n774), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(G283), .A2(new_n778), .B1(new_n781), .B2(G294), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1240), .A2(new_n1050), .A3(new_n1241), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n1232), .A2(new_n1236), .B1(new_n1238), .B2(new_n1242), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1243), .A2(KEYINPUT120), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n747), .B1(new_n1243), .B2(KEYINPUT120), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1231), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1229), .B1(new_n1230), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1228), .A2(new_n1247), .ZN(G381));
  NOR2_X1   g1048(.A1(G375), .A2(G378), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1005), .A2(new_n1099), .A3(new_n1030), .ZN(new_n1251));
  INV_X1    g1051(.A(G384), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(G393), .A2(G396), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  OR4_X1    g1054(.A1(G381), .A2(new_n1250), .A3(new_n1251), .A4(new_n1254), .ZN(G407));
  OAI211_X1 g1055(.A(G407), .B(G213), .C1(G343), .C2(new_n1250), .ZN(G409));
  AND2_X1   g1056(.A1(G393), .A2(G396), .ZN(new_n1257));
  OAI21_X1  g1057(.A(KEYINPUT125), .B1(new_n1257), .B2(new_n1253), .ZN(new_n1258));
  AND2_X1   g1058(.A1(new_n1251), .A2(new_n1258), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1257), .A2(new_n1253), .A3(KEYINPUT125), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(G387), .A2(G390), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1259), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1261), .B1(new_n1259), .B2(new_n1262), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT62), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G378), .B(new_n1215), .C1(new_n1223), .C2(new_n1224), .ZN(new_n1267));
  INV_X1    g1067(.A(G378), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1189), .A2(new_n1226), .A3(new_n1217), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1187), .A2(new_n1004), .A3(new_n1179), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1214), .A2(new_n1190), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(KEYINPUT121), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT121), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1270), .A2(new_n1274), .A3(new_n1271), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1273), .A2(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1268), .B1(new_n1269), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1267), .A2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n677), .A2(G213), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT60), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1227), .B1(new_n1135), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(KEYINPUT122), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT122), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1283), .B(new_n1227), .C1(new_n1135), .C2(new_n1280), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1227), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n697), .B1(new_n1285), .B2(KEYINPUT60), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1282), .A2(new_n1284), .A3(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1287), .A2(G384), .A3(new_n1247), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(G384), .B1(new_n1287), .B2(new_n1247), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  AND4_X1   g1091(.A1(new_n1266), .A2(new_n1278), .A3(new_n1279), .A4(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1279), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1293), .B1(new_n1267), .B2(new_n1277), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1266), .B1(new_n1294), .B2(new_n1291), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1292), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT61), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1287), .A2(new_n1247), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1252), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT123), .ZN(new_n1300));
  INV_X1    g1100(.A(G2897), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1279), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1302), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1303));
  AND3_X1   g1103(.A1(new_n1299), .A2(new_n1288), .A3(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1293), .A2(G2897), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1305), .B1(new_n1299), .B2(new_n1288), .ZN(new_n1306));
  OAI21_X1  g1106(.A(KEYINPUT124), .B1(new_n1304), .B2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT124), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1299), .A2(new_n1288), .A3(new_n1303), .ZN(new_n1309));
  OAI211_X1 g1109(.A(new_n1308), .B(new_n1309), .C1(new_n1291), .C2(new_n1305), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1307), .A2(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1297), .B1(new_n1294), .B2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT126), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1265), .B1(new_n1296), .B2(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1313), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1316));
  OAI211_X1 g1116(.A(new_n1316), .B(new_n1297), .C1(new_n1294), .C2(new_n1311), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1278), .A2(new_n1279), .A3(new_n1291), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT63), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1294), .A2(KEYINPUT63), .A3(new_n1291), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1317), .B1(new_n1322), .B2(new_n1265), .ZN(new_n1323));
  OAI21_X1  g1123(.A(KEYINPUT127), .B1(new_n1315), .B2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1265), .ZN(new_n1325));
  AND2_X1   g1125(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1318), .A2(KEYINPUT62), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1294), .A2(new_n1266), .A3(new_n1291), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1325), .B1(new_n1326), .B2(new_n1329), .ZN(new_n1330));
  AND3_X1   g1130(.A1(new_n1294), .A2(KEYINPUT63), .A3(new_n1291), .ZN(new_n1331));
  AOI21_X1  g1131(.A(KEYINPUT63), .B1(new_n1294), .B2(new_n1291), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1265), .B1(new_n1331), .B2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1317), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT127), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1330), .A2(new_n1335), .A3(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1324), .A2(new_n1337), .ZN(G405));
  XNOR2_X1  g1138(.A(G375), .B(G378), .ZN(new_n1339));
  XNOR2_X1  g1139(.A(new_n1339), .B(new_n1291), .ZN(new_n1340));
  XNOR2_X1  g1140(.A(new_n1340), .B(new_n1265), .ZN(G402));
endmodule


