

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581;

  NOR2_X2 U321 ( .A1(n517), .A2(n447), .ZN(n559) );
  XNOR2_X1 U322 ( .A(n419), .B(n418), .ZN(n555) );
  XNOR2_X1 U323 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n289) );
  INV_X1 U324 ( .A(G134GAT), .ZN(n404) );
  XNOR2_X1 U325 ( .A(n405), .B(n404), .ZN(n406) );
  NOR2_X1 U326 ( .A1(n486), .A2(n445), .ZN(n561) );
  XNOR2_X1 U327 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U328 ( .A(KEYINPUT101), .B(KEYINPUT36), .ZN(n423) );
  XNOR2_X1 U329 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U330 ( .A(n536), .B(n423), .ZN(n579) );
  INV_X1 U331 ( .A(G190GAT), .ZN(n453) );
  XNOR2_X1 U332 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U333 ( .A(n456), .B(n455), .ZN(G1351GAT) );
  XOR2_X1 U334 ( .A(G15GAT), .B(G127GAT), .Z(n348) );
  XOR2_X1 U335 ( .A(KEYINPUT87), .B(G190GAT), .Z(n291) );
  XNOR2_X1 U336 ( .A(G43GAT), .B(G99GAT), .ZN(n290) );
  XNOR2_X1 U337 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U338 ( .A(n348), .B(n292), .Z(n294) );
  NAND2_X1 U339 ( .A1(G227GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U340 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U341 ( .A(n295), .B(KEYINPUT88), .Z(n299) );
  XOR2_X1 U342 ( .A(G120GAT), .B(KEYINPUT0), .Z(n297) );
  XNOR2_X1 U343 ( .A(G113GAT), .B(G134GAT), .ZN(n296) );
  XNOR2_X1 U344 ( .A(n297), .B(n296), .ZN(n334) );
  XNOR2_X1 U345 ( .A(n334), .B(KEYINPUT83), .ZN(n298) );
  XNOR2_X1 U346 ( .A(n299), .B(n298), .ZN(n309) );
  XOR2_X1 U347 ( .A(KEYINPUT17), .B(KEYINPUT85), .Z(n301) );
  XNOR2_X1 U348 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n300) );
  XNOR2_X1 U349 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U350 ( .A(n302), .B(KEYINPUT86), .Z(n304) );
  XNOR2_X1 U351 ( .A(G169GAT), .B(G183GAT), .ZN(n303) );
  XNOR2_X1 U352 ( .A(n304), .B(n303), .ZN(n440) );
  XOR2_X1 U353 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n306) );
  XNOR2_X1 U354 ( .A(G176GAT), .B(G71GAT), .ZN(n305) );
  XNOR2_X1 U355 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U356 ( .A(n440), .B(n307), .Z(n308) );
  XNOR2_X1 U357 ( .A(n309), .B(n308), .ZN(n517) );
  XOR2_X1 U358 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n311) );
  XNOR2_X1 U359 ( .A(G204GAT), .B(KEYINPUT89), .ZN(n310) );
  XNOR2_X1 U360 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U361 ( .A(KEYINPUT24), .B(KEYINPUT92), .Z(n313) );
  XOR2_X1 U362 ( .A(G141GAT), .B(G22GAT), .Z(n369) );
  XOR2_X1 U363 ( .A(G50GAT), .B(G162GAT), .Z(n413) );
  XNOR2_X1 U364 ( .A(n369), .B(n413), .ZN(n312) );
  XNOR2_X1 U365 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U366 ( .A(n315), .B(n314), .Z(n317) );
  NAND2_X1 U367 ( .A1(G228GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U368 ( .A(n317), .B(n316), .ZN(n320) );
  XOR2_X1 U369 ( .A(G155GAT), .B(KEYINPUT2), .Z(n319) );
  XNOR2_X1 U370 ( .A(KEYINPUT3), .B(KEYINPUT91), .ZN(n318) );
  XNOR2_X1 U371 ( .A(n319), .B(n318), .ZN(n333) );
  XOR2_X1 U372 ( .A(n320), .B(n333), .Z(n326) );
  XOR2_X1 U373 ( .A(KEYINPUT90), .B(G218GAT), .Z(n322) );
  XNOR2_X1 U374 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n321) );
  XNOR2_X1 U375 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U376 ( .A(G197GAT), .B(n323), .Z(n439) );
  XNOR2_X1 U377 ( .A(G106GAT), .B(G78GAT), .ZN(n324) );
  XNOR2_X1 U378 ( .A(n324), .B(G148GAT), .ZN(n385) );
  XNOR2_X1 U379 ( .A(n439), .B(n385), .ZN(n325) );
  XNOR2_X1 U380 ( .A(n326), .B(n325), .ZN(n463) );
  XOR2_X1 U381 ( .A(KEYINPUT94), .B(KEYINPUT6), .Z(n328) );
  XNOR2_X1 U382 ( .A(G1GAT), .B(G57GAT), .ZN(n327) );
  XNOR2_X1 U383 ( .A(n328), .B(n327), .ZN(n344) );
  XOR2_X1 U384 ( .A(G162GAT), .B(G148GAT), .Z(n330) );
  XNOR2_X1 U385 ( .A(G141GAT), .B(G127GAT), .ZN(n329) );
  XNOR2_X1 U386 ( .A(n330), .B(n329), .ZN(n332) );
  XOR2_X1 U387 ( .A(G29GAT), .B(G85GAT), .Z(n331) );
  XNOR2_X1 U388 ( .A(n332), .B(n331), .ZN(n340) );
  XNOR2_X1 U389 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U390 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n336) );
  XNOR2_X1 U391 ( .A(KEYINPUT1), .B(KEYINPUT93), .ZN(n335) );
  XNOR2_X1 U392 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U393 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U394 ( .A(n340), .B(n339), .ZN(n342) );
  NAND2_X1 U395 ( .A1(G225GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U396 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U397 ( .A(n344), .B(n343), .ZN(n486) );
  XOR2_X1 U398 ( .A(KEYINPUT47), .B(KEYINPUT109), .Z(n422) );
  XOR2_X1 U399 ( .A(KEYINPUT13), .B(KEYINPUT72), .Z(n346) );
  XNOR2_X1 U400 ( .A(G71GAT), .B(KEYINPUT71), .ZN(n345) );
  XNOR2_X1 U401 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U402 ( .A(G57GAT), .B(n347), .Z(n398) );
  XOR2_X1 U403 ( .A(G78GAT), .B(n348), .Z(n351) );
  XNOR2_X1 U404 ( .A(G8GAT), .B(G1GAT), .ZN(n349) );
  XNOR2_X1 U405 ( .A(n349), .B(KEYINPUT70), .ZN(n380) );
  XNOR2_X1 U406 ( .A(n380), .B(G183GAT), .ZN(n350) );
  XNOR2_X1 U407 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U408 ( .A(n398), .B(n352), .ZN(n365) );
  XOR2_X1 U409 ( .A(G64GAT), .B(G155GAT), .Z(n354) );
  XNOR2_X1 U410 ( .A(G22GAT), .B(G211GAT), .ZN(n353) );
  XNOR2_X1 U411 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U412 ( .A(KEYINPUT15), .B(KEYINPUT81), .Z(n356) );
  XNOR2_X1 U413 ( .A(KEYINPUT80), .B(KEYINPUT79), .ZN(n355) );
  XNOR2_X1 U414 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U415 ( .A(n358), .B(n357), .Z(n363) );
  XOR2_X1 U416 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n360) );
  NAND2_X1 U417 ( .A1(G231GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U418 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U419 ( .A(KEYINPUT78), .B(n361), .ZN(n362) );
  XNOR2_X1 U420 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U421 ( .A(n365), .B(n364), .ZN(n572) );
  XOR2_X1 U422 ( .A(G15GAT), .B(G50GAT), .Z(n367) );
  XNOR2_X1 U423 ( .A(G169GAT), .B(G36GAT), .ZN(n366) );
  XNOR2_X1 U424 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U425 ( .A(n369), .B(n368), .Z(n371) );
  NAND2_X1 U426 ( .A1(G229GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U427 ( .A(n371), .B(n370), .ZN(n384) );
  XOR2_X1 U428 ( .A(KEYINPUT29), .B(KEYINPUT68), .Z(n373) );
  XNOR2_X1 U429 ( .A(KEYINPUT67), .B(KEYINPUT69), .ZN(n372) );
  XNOR2_X1 U430 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U431 ( .A(KEYINPUT66), .B(KEYINPUT30), .Z(n375) );
  XNOR2_X1 U432 ( .A(G113GAT), .B(G197GAT), .ZN(n374) );
  XNOR2_X1 U433 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U434 ( .A(n377), .B(n376), .Z(n382) );
  XOR2_X1 U435 ( .A(G29GAT), .B(G43GAT), .Z(n379) );
  XNOR2_X1 U436 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n378) );
  XNOR2_X1 U437 ( .A(n379), .B(n378), .ZN(n407) );
  XNOR2_X1 U438 ( .A(n407), .B(n380), .ZN(n381) );
  XNOR2_X1 U439 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U440 ( .A(n384), .B(n383), .Z(n544) );
  XOR2_X1 U441 ( .A(G99GAT), .B(G85GAT), .Z(n401) );
  XOR2_X1 U442 ( .A(KEYINPUT31), .B(n401), .Z(n387) );
  XNOR2_X1 U443 ( .A(G120GAT), .B(n385), .ZN(n386) );
  XNOR2_X1 U444 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U445 ( .A(KEYINPUT73), .B(KEYINPUT32), .Z(n389) );
  NAND2_X1 U446 ( .A1(G230GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U447 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U448 ( .A(n391), .B(n390), .Z(n396) );
  XOR2_X1 U449 ( .A(KEYINPUT74), .B(G64GAT), .Z(n393) );
  XNOR2_X1 U450 ( .A(G176GAT), .B(G92GAT), .ZN(n392) );
  XNOR2_X1 U451 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U452 ( .A(G204GAT), .B(n394), .Z(n437) );
  XNOR2_X1 U453 ( .A(n437), .B(KEYINPUT33), .ZN(n395) );
  XNOR2_X1 U454 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U455 ( .A(n398), .B(n397), .ZN(n568) );
  XNOR2_X1 U456 ( .A(KEYINPUT41), .B(n568), .ZN(n549) );
  NOR2_X1 U457 ( .A1(n544), .A2(n549), .ZN(n399) );
  XNOR2_X1 U458 ( .A(n399), .B(KEYINPUT46), .ZN(n400) );
  NOR2_X1 U459 ( .A1(n572), .A2(n400), .ZN(n420) );
  XOR2_X1 U460 ( .A(G36GAT), .B(G190GAT), .Z(n434) );
  XOR2_X1 U461 ( .A(KEYINPUT76), .B(n434), .Z(n403) );
  XNOR2_X1 U462 ( .A(G218GAT), .B(n401), .ZN(n402) );
  XOR2_X1 U463 ( .A(n403), .B(n402), .Z(n409) );
  NAND2_X1 U464 ( .A1(G232GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U465 ( .A(n409), .B(n408), .ZN(n419) );
  XOR2_X1 U466 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n411) );
  XNOR2_X1 U467 ( .A(G106GAT), .B(KEYINPUT64), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U469 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U470 ( .A(KEYINPUT77), .B(KEYINPUT75), .Z(n415) );
  XNOR2_X1 U471 ( .A(KEYINPUT9), .B(G92GAT), .ZN(n414) );
  XNOR2_X1 U472 ( .A(n415), .B(n414), .ZN(n416) );
  NAND2_X1 U473 ( .A1(n420), .A2(n555), .ZN(n421) );
  XNOR2_X1 U474 ( .A(n422), .B(n421), .ZN(n429) );
  INV_X1 U475 ( .A(n555), .ZN(n536) );
  INV_X1 U476 ( .A(n572), .ZN(n552) );
  NOR2_X1 U477 ( .A1(n579), .A2(n552), .ZN(n424) );
  XNOR2_X1 U478 ( .A(KEYINPUT45), .B(n424), .ZN(n426) );
  INV_X1 U479 ( .A(n568), .ZN(n425) );
  NAND2_X1 U480 ( .A1(n426), .A2(n425), .ZN(n427) );
  INV_X1 U481 ( .A(n544), .ZN(n564) );
  NOR2_X1 U482 ( .A1(n427), .A2(n564), .ZN(n428) );
  NOR2_X1 U483 ( .A1(n429), .A2(n428), .ZN(n430) );
  XNOR2_X1 U484 ( .A(KEYINPUT48), .B(n430), .ZN(n542) );
  XOR2_X1 U485 ( .A(KEYINPUT95), .B(KEYINPUT97), .Z(n432) );
  XNOR2_X1 U486 ( .A(G8GAT), .B(KEYINPUT96), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U488 ( .A(n434), .B(n433), .Z(n436) );
  NAND2_X1 U489 ( .A1(G226GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n438) );
  XOR2_X1 U491 ( .A(n438), .B(n437), .Z(n442) );
  XNOR2_X1 U492 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U493 ( .A(n442), .B(n441), .ZN(n514) );
  XOR2_X1 U494 ( .A(KEYINPUT117), .B(n514), .Z(n443) );
  NOR2_X1 U495 ( .A1(n542), .A2(n443), .ZN(n444) );
  XOR2_X1 U496 ( .A(KEYINPUT54), .B(n444), .Z(n445) );
  NAND2_X1 U497 ( .A1(n463), .A2(n561), .ZN(n446) );
  XOR2_X1 U498 ( .A(KEYINPUT55), .B(n446), .Z(n447) );
  INV_X1 U499 ( .A(n549), .ZN(n528) );
  NAND2_X1 U500 ( .A1(n559), .A2(n528), .ZN(n452) );
  XOR2_X1 U501 ( .A(KEYINPUT121), .B(KEYINPUT120), .Z(n449) );
  XNOR2_X1 U502 ( .A(KEYINPUT119), .B(KEYINPUT57), .ZN(n448) );
  XNOR2_X1 U503 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U504 ( .A(n450), .B(n289), .ZN(n451) );
  XNOR2_X1 U505 ( .A(n452), .B(n451), .ZN(G1349GAT) );
  NAND2_X1 U506 ( .A1(n559), .A2(n536), .ZN(n456) );
  XOR2_X1 U507 ( .A(KEYINPUT122), .B(KEYINPUT58), .Z(n454) );
  NOR2_X1 U508 ( .A1(n544), .A2(n568), .ZN(n484) );
  XOR2_X1 U509 ( .A(KEYINPUT82), .B(KEYINPUT16), .Z(n458) );
  NAND2_X1 U510 ( .A1(n572), .A2(n555), .ZN(n457) );
  XNOR2_X1 U511 ( .A(n458), .B(n457), .ZN(n470) );
  XNOR2_X1 U512 ( .A(n463), .B(KEYINPUT65), .ZN(n459) );
  XNOR2_X1 U513 ( .A(n459), .B(KEYINPUT28), .ZN(n504) );
  XOR2_X1 U514 ( .A(n514), .B(KEYINPUT27), .Z(n461) );
  NAND2_X1 U515 ( .A1(n461), .A2(n486), .ZN(n541) );
  NOR2_X1 U516 ( .A1(n504), .A2(n541), .ZN(n523) );
  NAND2_X1 U517 ( .A1(n523), .A2(n517), .ZN(n469) );
  INV_X1 U518 ( .A(n517), .ZN(n524) );
  NOR2_X1 U519 ( .A1(n463), .A2(n524), .ZN(n460) );
  XNOR2_X1 U520 ( .A(n460), .B(KEYINPUT26), .ZN(n562) );
  NAND2_X1 U521 ( .A1(n562), .A2(n461), .ZN(n466) );
  INV_X1 U522 ( .A(n514), .ZN(n490) );
  NAND2_X1 U523 ( .A1(n524), .A2(n490), .ZN(n462) );
  NAND2_X1 U524 ( .A1(n463), .A2(n462), .ZN(n464) );
  XOR2_X1 U525 ( .A(KEYINPUT25), .B(n464), .Z(n465) );
  NAND2_X1 U526 ( .A1(n466), .A2(n465), .ZN(n467) );
  INV_X1 U527 ( .A(n486), .ZN(n511) );
  NAND2_X1 U528 ( .A1(n467), .A2(n511), .ZN(n468) );
  NAND2_X1 U529 ( .A1(n469), .A2(n468), .ZN(n482) );
  AND2_X1 U530 ( .A1(n470), .A2(n482), .ZN(n499) );
  NAND2_X1 U531 ( .A1(n484), .A2(n499), .ZN(n471) );
  XOR2_X1 U532 ( .A(KEYINPUT98), .B(n471), .Z(n479) );
  NAND2_X1 U533 ( .A1(n479), .A2(n486), .ZN(n474) );
  XOR2_X1 U534 ( .A(G1GAT), .B(KEYINPUT99), .Z(n472) );
  XNOR2_X1 U535 ( .A(KEYINPUT34), .B(n472), .ZN(n473) );
  XNOR2_X1 U536 ( .A(n474), .B(n473), .ZN(G1324GAT) );
  NAND2_X1 U537 ( .A1(n479), .A2(n490), .ZN(n475) );
  XNOR2_X1 U538 ( .A(n475), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U539 ( .A(KEYINPUT100), .B(KEYINPUT35), .Z(n477) );
  NAND2_X1 U540 ( .A1(n524), .A2(n479), .ZN(n476) );
  XNOR2_X1 U541 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U542 ( .A(G15GAT), .B(n478), .ZN(G1326GAT) );
  NAND2_X1 U543 ( .A1(n479), .A2(n504), .ZN(n480) );
  XNOR2_X1 U544 ( .A(n480), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT102), .B(KEYINPUT39), .Z(n488) );
  NOR2_X1 U546 ( .A1(n572), .A2(n579), .ZN(n481) );
  NAND2_X1 U547 ( .A1(n482), .A2(n481), .ZN(n483) );
  XNOR2_X1 U548 ( .A(KEYINPUT37), .B(n483), .ZN(n508) );
  NAND2_X1 U549 ( .A1(n508), .A2(n484), .ZN(n485) );
  XOR2_X1 U550 ( .A(KEYINPUT38), .B(n485), .Z(n495) );
  NAND2_X1 U551 ( .A1(n495), .A2(n486), .ZN(n487) );
  XNOR2_X1 U552 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U553 ( .A(G29GAT), .B(n489), .ZN(G1328GAT) );
  XOR2_X1 U554 ( .A(G36GAT), .B(KEYINPUT103), .Z(n492) );
  NAND2_X1 U555 ( .A1(n495), .A2(n490), .ZN(n491) );
  XNOR2_X1 U556 ( .A(n492), .B(n491), .ZN(G1329GAT) );
  NAND2_X1 U557 ( .A1(n495), .A2(n524), .ZN(n493) );
  XNOR2_X1 U558 ( .A(n493), .B(KEYINPUT40), .ZN(n494) );
  XNOR2_X1 U559 ( .A(G43GAT), .B(n494), .ZN(G1330GAT) );
  NAND2_X1 U560 ( .A1(n495), .A2(n504), .ZN(n496) );
  XNOR2_X1 U561 ( .A(n496), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT105), .B(KEYINPUT42), .Z(n498) );
  XNOR2_X1 U563 ( .A(G57GAT), .B(KEYINPUT104), .ZN(n497) );
  XNOR2_X1 U564 ( .A(n498), .B(n497), .ZN(n501) );
  NOR2_X1 U565 ( .A1(n549), .A2(n564), .ZN(n509) );
  NAND2_X1 U566 ( .A1(n509), .A2(n499), .ZN(n505) );
  NOR2_X1 U567 ( .A1(n511), .A2(n505), .ZN(n500) );
  XOR2_X1 U568 ( .A(n501), .B(n500), .Z(G1332GAT) );
  NOR2_X1 U569 ( .A1(n514), .A2(n505), .ZN(n502) );
  XOR2_X1 U570 ( .A(G64GAT), .B(n502), .Z(G1333GAT) );
  NOR2_X1 U571 ( .A1(n517), .A2(n505), .ZN(n503) );
  XOR2_X1 U572 ( .A(G71GAT), .B(n503), .Z(G1334GAT) );
  INV_X1 U573 ( .A(n504), .ZN(n519) );
  NOR2_X1 U574 ( .A1(n519), .A2(n505), .ZN(n507) );
  XNOR2_X1 U575 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n506) );
  XNOR2_X1 U576 ( .A(n507), .B(n506), .ZN(G1335GAT) );
  NAND2_X1 U577 ( .A1(n509), .A2(n508), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n510), .B(KEYINPUT106), .ZN(n520) );
  NOR2_X1 U579 ( .A1(n511), .A2(n520), .ZN(n512) );
  XNOR2_X1 U580 ( .A(G85GAT), .B(n512), .ZN(n513) );
  XNOR2_X1 U581 ( .A(n513), .B(KEYINPUT107), .ZN(G1336GAT) );
  NOR2_X1 U582 ( .A1(n514), .A2(n520), .ZN(n515) );
  XOR2_X1 U583 ( .A(KEYINPUT108), .B(n515), .Z(n516) );
  XNOR2_X1 U584 ( .A(G92GAT), .B(n516), .ZN(G1337GAT) );
  NOR2_X1 U585 ( .A1(n520), .A2(n517), .ZN(n518) );
  XOR2_X1 U586 ( .A(G99GAT), .B(n518), .Z(G1338GAT) );
  NOR2_X1 U587 ( .A1(n520), .A2(n519), .ZN(n521) );
  XOR2_X1 U588 ( .A(KEYINPUT44), .B(n521), .Z(n522) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n522), .ZN(G1339GAT) );
  NAND2_X1 U590 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X1 U591 ( .A1(n542), .A2(n525), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n564), .A2(n537), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n526), .B(KEYINPUT110), .ZN(n527) );
  XNOR2_X1 U594 ( .A(G113GAT), .B(n527), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT49), .B(KEYINPUT112), .Z(n530) );
  NAND2_X1 U596 ( .A1(n537), .A2(n528), .ZN(n529) );
  XNOR2_X1 U597 ( .A(n530), .B(n529), .ZN(n532) );
  XOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT111), .Z(n531) );
  XNOR2_X1 U599 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT113), .B(KEYINPUT50), .Z(n534) );
  NAND2_X1 U601 ( .A1(n537), .A2(n572), .ZN(n533) );
  XNOR2_X1 U602 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n539) );
  NAND2_X1 U605 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U607 ( .A(G134GAT), .B(n540), .ZN(G1343GAT) );
  NOR2_X1 U608 ( .A1(n542), .A2(n541), .ZN(n543) );
  NAND2_X1 U609 ( .A1(n543), .A2(n562), .ZN(n554) );
  NOR2_X1 U610 ( .A1(n544), .A2(n554), .ZN(n546) );
  XNOR2_X1 U611 ( .A(G141GAT), .B(KEYINPUT115), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(G1344GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n548) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n551) );
  NOR2_X1 U616 ( .A1(n549), .A2(n554), .ZN(n550) );
  XOR2_X1 U617 ( .A(n551), .B(n550), .Z(G1345GAT) );
  NOR2_X1 U618 ( .A1(n552), .A2(n554), .ZN(n553) );
  XOR2_X1 U619 ( .A(G155GAT), .B(n553), .Z(G1346GAT) );
  NOR2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U621 ( .A(G162GAT), .B(n556), .Z(G1347GAT) );
  NAND2_X1 U622 ( .A1(n564), .A2(n559), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(KEYINPUT118), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G169GAT), .B(n558), .ZN(G1348GAT) );
  NAND2_X1 U625 ( .A1(n559), .A2(n572), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n566) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(KEYINPUT123), .ZN(n577) );
  NAND2_X1 U630 ( .A1(n577), .A2(n564), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(n567), .ZN(G1352GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n570) );
  NAND2_X1 U634 ( .A1(n577), .A2(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(G204GAT), .B(n571), .ZN(G1353GAT) );
  XOR2_X1 U637 ( .A(G211GAT), .B(KEYINPUT125), .Z(n574) );
  NAND2_X1 U638 ( .A1(n577), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1354GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n576) );
  XNOR2_X1 U641 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n581) );
  INV_X1 U643 ( .A(n577), .ZN(n578) );
  NOR2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U645 ( .A(n581), .B(n580), .Z(G1355GAT) );
endmodule

