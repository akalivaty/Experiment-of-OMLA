//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 1 0 1 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 1 1 0 1 1 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n209), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  OR2_X1    g0016(.A1(new_n216), .A2(KEYINPUT1), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT65), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n209), .A2(G13), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n219), .B(G250), .C1(G257), .C2(G264), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT0), .ZN(new_n221));
  AND2_X1   g0021(.A1(KEYINPUT64), .A2(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(KEYINPUT64), .A2(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n201), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n221), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n218), .B(new_n230), .C1(KEYINPUT1), .C2(new_n216), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G58), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  AND2_X1   g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  NOR2_X1   g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  OAI211_X1 g0048(.A(G232), .B(G1698), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G1698), .ZN(new_n250));
  OAI211_X1 g0050(.A(G226), .B(new_n250), .C1(new_n247), .C2(new_n248), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G97), .ZN(new_n253));
  OAI211_X1 g0053(.A(new_n249), .B(new_n251), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G1), .A3(G13), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G41), .ZN(new_n259));
  INV_X1    g0059(.A(G45), .ZN(new_n260));
  AOI21_X1  g0060(.A(G1), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AND3_X1   g0061(.A1(new_n261), .A2(new_n256), .A3(G274), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n257), .A2(new_n261), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n262), .B1(G238), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT13), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n258), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n265), .B1(new_n258), .B2(new_n264), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G169), .ZN(new_n270));
  OAI21_X1  g0070(.A(KEYINPUT14), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT14), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n272), .B(G169), .C1(new_n267), .C2(new_n268), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT72), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n274), .B1(new_n269), .B2(G179), .ZN(new_n275));
  INV_X1    g0075(.A(G179), .ZN(new_n276));
  NOR4_X1   g0076(.A1(new_n267), .A2(new_n268), .A3(KEYINPUT72), .A4(new_n276), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n271), .B(new_n273), .C1(new_n275), .C2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G68), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(new_n282), .B(KEYINPUT12), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n279), .A2(new_n225), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT68), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n286), .B1(new_n207), .B2(G1), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n206), .A2(KEYINPUT68), .A3(G20), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OR2_X1    g0089(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n283), .B1(new_n290), .B2(new_n281), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n284), .A2(new_n225), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT64), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n207), .ZN(new_n295));
  NAND2_X1  g0095(.A1(KEYINPUT64), .A2(G20), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n295), .A2(G33), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT67), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n295), .A2(KEYINPUT67), .A3(G33), .A4(new_n296), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n299), .A2(G77), .A3(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(G20), .A2(G33), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n302), .A2(G50), .B1(G20), .B2(new_n281), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n293), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n291), .B1(KEYINPUT11), .B2(new_n304), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n304), .A2(KEYINPUT11), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n278), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n268), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n309), .A2(G190), .A3(new_n266), .ZN(new_n310));
  OAI21_X1  g0110(.A(G200), .B1(new_n267), .B2(new_n268), .ZN(new_n311));
  AND4_X1   g0111(.A1(new_n306), .A2(new_n310), .A3(new_n311), .A4(new_n305), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  OR2_X1    g0113(.A1(KEYINPUT3), .A2(G33), .ZN(new_n314));
  NAND2_X1  g0114(.A1(KEYINPUT3), .A2(G33), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n316), .A2(G232), .A3(new_n250), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(G238), .A3(G1698), .ZN(new_n318));
  INV_X1    g0118(.A(G107), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n317), .B(new_n318), .C1(new_n319), .C2(new_n316), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n257), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n262), .B1(G244), .B2(new_n263), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G190), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n325), .B1(G200), .B2(new_n323), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n279), .A2(G77), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n290), .B1(new_n224), .B2(new_n293), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n327), .B1(new_n328), .B2(G77), .ZN(new_n329));
  XOR2_X1   g0129(.A(KEYINPUT15), .B(G87), .Z(new_n330));
  NAND3_X1  g0130(.A1(new_n299), .A2(new_n300), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G58), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT8), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT8), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G58), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n302), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n293), .B1(new_n331), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT70), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n329), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n340), .B1(new_n329), .B2(new_n339), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n326), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n323), .A2(G179), .ZN(new_n345));
  AOI21_X1  g0145(.A(G169), .B1(new_n321), .B2(new_n322), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n341), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n347), .B1(new_n348), .B2(new_n342), .ZN(new_n349));
  AND4_X1   g0149(.A1(new_n308), .A2(new_n313), .A3(new_n344), .A4(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n332), .A2(KEYINPUT66), .A3(KEYINPUT8), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT66), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n333), .A2(new_n335), .A3(new_n352), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n351), .B(new_n353), .C1(new_n285), .C2(new_n289), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n351), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n279), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT73), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n354), .A2(new_n356), .A3(KEYINPUT73), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n332), .A2(new_n281), .ZN(new_n362));
  OAI21_X1  g0162(.A(G20), .B1(new_n362), .B2(new_n201), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n302), .A2(G159), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n314), .A2(new_n207), .A3(new_n315), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n281), .B1(new_n367), .B2(KEYINPUT7), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n247), .A2(new_n248), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT7), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n224), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n366), .B(KEYINPUT16), .C1(new_n369), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n292), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n295), .A2(new_n296), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT7), .B1(new_n316), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n370), .A2(new_n371), .A3(new_n207), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(G68), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(KEYINPUT16), .B1(new_n379), .B2(new_n366), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n361), .B1(new_n375), .B2(new_n380), .ZN(new_n381));
  OAI211_X1 g0181(.A(G223), .B(new_n250), .C1(new_n247), .C2(new_n248), .ZN(new_n382));
  OAI211_X1 g0182(.A(G226), .B(G1698), .C1(new_n247), .C2(new_n248), .ZN(new_n383));
  INV_X1    g0183(.A(G87), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n382), .B(new_n383), .C1(new_n252), .C2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n257), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n256), .A2(G274), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n263), .A2(G232), .B1(new_n387), .B2(new_n261), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(new_n388), .A3(G179), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n386), .A2(new_n388), .ZN(new_n390));
  OAI211_X1 g0190(.A(KEYINPUT74), .B(new_n389), .C1(new_n390), .C2(new_n270), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT74), .ZN(new_n392));
  AND3_X1   g0192(.A1(new_n386), .A2(new_n388), .A3(G179), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n270), .B1(new_n386), .B2(new_n388), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n381), .A2(new_n391), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT18), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT18), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n381), .A2(new_n391), .A3(new_n395), .A4(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT17), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n390), .A2(G190), .ZN(new_n401));
  INV_X1    g0201(.A(G200), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n402), .B1(new_n386), .B2(new_n388), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n400), .B1(new_n405), .B2(new_n381), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n365), .B1(new_n372), .B2(new_n368), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n293), .B1(new_n407), .B2(KEYINPUT16), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n379), .A2(new_n366), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT16), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n408), .A2(new_n411), .B1(new_n359), .B2(new_n360), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n403), .B1(G190), .B2(new_n390), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(KEYINPUT17), .A3(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n397), .A2(new_n399), .A3(new_n406), .A4(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n350), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(G1698), .B1(new_n314), .B2(new_n315), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(G222), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n316), .A2(G223), .A3(G1698), .ZN(new_n420));
  INV_X1    g0220(.A(G77), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n419), .B(new_n420), .C1(new_n421), .C2(new_n316), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n257), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n262), .B1(G226), .B2(new_n263), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OR3_X1    g0225(.A1(new_n425), .A2(KEYINPUT69), .A3(G179), .ZN(new_n426));
  OAI21_X1  g0226(.A(KEYINPUT69), .B1(new_n425), .B2(G179), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n355), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n429), .A2(new_n299), .A3(new_n300), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n302), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n293), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n280), .A2(new_n202), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n290), .B2(new_n202), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(G169), .B1(new_n423), .B2(new_n424), .ZN(new_n436));
  NOR3_X1   g0236(.A1(new_n428), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT71), .B1(new_n432), .B2(new_n434), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n432), .A2(KEYINPUT71), .A3(new_n434), .ZN(new_n441));
  OAI21_X1  g0241(.A(KEYINPUT9), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n441), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT9), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(new_n444), .A3(new_n439), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT10), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n425), .A2(new_n324), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n448), .B1(G200), .B2(new_n425), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n446), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n447), .B1(new_n446), .B2(new_n449), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n438), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT75), .B1(new_n417), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n452), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n437), .B1(new_n455), .B2(new_n450), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT75), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n456), .A2(new_n350), .A3(new_n416), .A4(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n206), .A2(G33), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n293), .A2(new_n279), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n330), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT78), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n299), .A2(G97), .A3(new_n300), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT19), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT77), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n465), .A2(KEYINPUT77), .A3(new_n466), .ZN(new_n470));
  NOR2_X1   g0270(.A1(G97), .A2(G107), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n384), .ZN(new_n472));
  NOR3_X1   g0272(.A1(new_n466), .A2(new_n252), .A3(new_n253), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n472), .B1(new_n473), .B2(new_n376), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n316), .A2(new_n224), .A3(G68), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n469), .A2(new_n470), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n292), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n330), .A2(new_n279), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n464), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  AOI211_X1 g0282(.A(KEYINPUT78), .B(new_n480), .C1(new_n478), .C2(new_n292), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n463), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OR2_X1    g0284(.A1(new_n250), .A2(G244), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n316), .B(new_n485), .C1(G238), .C2(G1698), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G116), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n256), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n260), .A2(G1), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n387), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n256), .B(G250), .C1(G1), .C2(new_n260), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n276), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(G169), .B2(new_n493), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n461), .A2(new_n384), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n476), .B1(new_n467), .B2(new_n468), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n293), .B1(new_n498), .B2(new_n470), .ZN(new_n499));
  OAI21_X1  g0299(.A(KEYINPUT78), .B1(new_n499), .B2(new_n480), .ZN(new_n500));
  AND3_X1   g0300(.A1(new_n465), .A2(KEYINPUT77), .A3(new_n466), .ZN(new_n501));
  AOI21_X1  g0301(.A(KEYINPUT77), .B1(new_n465), .B2(new_n466), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n501), .A2(new_n502), .A3(new_n476), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n464), .B(new_n481), .C1(new_n503), .C2(new_n293), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n497), .B1(new_n500), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n493), .A2(new_n324), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n506), .B1(G200), .B2(new_n493), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n484), .A2(new_n496), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G33), .A2(G283), .ZN(new_n509));
  OAI211_X1 g0309(.A(G250), .B(G1698), .C1(new_n247), .C2(new_n248), .ZN(new_n510));
  OAI211_X1 g0310(.A(G244), .B(new_n250), .C1(new_n247), .C2(new_n248), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT4), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n509), .B(new_n510), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(KEYINPUT4), .B1(new_n418), .B2(G244), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n257), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  XNOR2_X1  g0315(.A(KEYINPUT5), .B(G41), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n516), .A2(G274), .A3(new_n256), .A4(new_n489), .ZN(new_n517));
  AND2_X1   g0317(.A1(KEYINPUT5), .A2(G41), .ZN(new_n518));
  NOR2_X1   g0318(.A1(KEYINPUT5), .A2(G41), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n489), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n520), .A2(G257), .A3(new_n256), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n515), .A2(new_n517), .A3(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT76), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n515), .A2(KEYINPUT76), .A3(new_n517), .A4(new_n521), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n524), .A2(G200), .A3(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n515), .A2(G190), .A3(new_n517), .A4(new_n521), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n371), .B1(new_n224), .B2(new_n370), .ZN(new_n528));
  NOR4_X1   g0328(.A1(new_n247), .A2(new_n248), .A3(KEYINPUT7), .A4(G20), .ZN(new_n529));
  NOR3_X1   g0329(.A1(new_n528), .A2(new_n529), .A3(new_n319), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n302), .A2(G77), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT6), .ZN(new_n532));
  NOR3_X1   g0332(.A1(new_n532), .A2(new_n253), .A3(G107), .ZN(new_n533));
  XNOR2_X1  g0333(.A(G97), .B(G107), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n533), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n531), .B1(new_n535), .B2(new_n224), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n292), .B1(new_n530), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n279), .A2(G97), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(new_n462), .B2(G97), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n527), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n270), .A2(new_n522), .B1(new_n537), .B2(new_n539), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n515), .A2(new_n521), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n542), .A2(new_n276), .A3(new_n517), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n526), .A2(new_n540), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n316), .A2(G257), .A3(G1698), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n316), .A2(G250), .A3(new_n250), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G294), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n257), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n520), .A2(G264), .A3(new_n256), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n517), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n553), .A2(new_n324), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n551), .B1(new_n257), .B2(new_n548), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n555), .A2(new_n402), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n280), .A2(KEYINPUT25), .A3(new_n319), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(KEYINPUT25), .B1(new_n280), .B2(new_n319), .ZN(new_n560));
  OAI22_X1  g0360(.A1(new_n559), .A2(new_n560), .B1(new_n461), .B2(new_n319), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n295), .B(new_n296), .C1(new_n247), .C2(new_n248), .ZN(new_n563));
  OAI21_X1  g0363(.A(KEYINPUT22), .B1(new_n563), .B2(new_n384), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT22), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n316), .A2(new_n224), .A3(new_n565), .A4(G87), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n568));
  OAI21_X1  g0368(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n569));
  OR2_X1    g0369(.A1(KEYINPUT23), .A2(G107), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n568), .B(new_n569), .C1(new_n224), .C2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT82), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n574), .A2(KEYINPUT24), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n293), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n571), .B1(new_n564), .B2(new_n566), .ZN(new_n577));
  XOR2_X1   g0377(.A(KEYINPUT82), .B(KEYINPUT24), .Z(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT83), .B1(new_n576), .B2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n575), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n292), .B1(new_n577), .B2(new_n582), .ZN(new_n583));
  AOI211_X1 g0383(.A(new_n578), .B(new_n571), .C1(new_n564), .C2(new_n566), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT83), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n557), .B(new_n562), .C1(new_n581), .C2(new_n586), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n544), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n585), .B1(new_n583), .B2(new_n584), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n573), .A2(new_n575), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n590), .A2(KEYINPUT83), .A3(new_n292), .A4(new_n580), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n561), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  AND4_X1   g0392(.A1(KEYINPUT84), .A2(new_n549), .A3(G179), .A4(new_n552), .ZN(new_n593));
  OAI21_X1  g0393(.A(KEYINPUT84), .B1(new_n555), .B2(new_n270), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n555), .A2(G179), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n520), .A2(G270), .A3(new_n256), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n517), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT79), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n598), .A2(KEYINPUT79), .A3(new_n517), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n316), .A2(G264), .A3(G1698), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n316), .A2(G257), .A3(new_n250), .ZN(new_n604));
  INV_X1    g0404(.A(G303), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n603), .B(new_n604), .C1(new_n605), .C2(new_n316), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n601), .A2(new_n602), .B1(new_n257), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n252), .A2(G97), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n295), .A2(new_n608), .A3(new_n296), .A4(new_n509), .ZN(new_n609));
  INV_X1    g0409(.A(G116), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n284), .A2(new_n225), .B1(G20), .B2(new_n610), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n609), .A2(KEYINPUT20), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT20), .B1(new_n609), .B2(new_n611), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n206), .A2(new_n610), .A3(G13), .A4(G20), .ZN(new_n615));
  XNOR2_X1  g0415(.A(new_n615), .B(KEYINPUT80), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n616), .B1(new_n610), .B2(new_n461), .ZN(new_n617));
  OAI21_X1  g0417(.A(G169), .B1(new_n614), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(KEYINPUT81), .B1(new_n607), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(KEYINPUT21), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT21), .ZN(new_n621));
  OAI211_X1 g0421(.A(KEYINPUT81), .B(new_n621), .C1(new_n607), .C2(new_n618), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n607), .B(G179), .C1(new_n614), .C2(new_n617), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n620), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n607), .A2(G190), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n614), .A2(new_n617), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n625), .B(new_n626), .C1(new_n402), .C2(new_n607), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NOR3_X1   g0428(.A1(new_n597), .A2(new_n624), .A3(new_n628), .ZN(new_n629));
  AND4_X1   g0429(.A1(new_n459), .A2(new_n508), .A3(new_n588), .A4(new_n629), .ZN(G372));
  INV_X1    g0430(.A(new_n497), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n631), .B(new_n507), .C1(new_n482), .C2(new_n483), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n541), .A2(new_n543), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n500), .A2(new_n504), .B1(new_n330), .B2(new_n462), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n632), .B(new_n634), .C1(new_n635), .C2(new_n495), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT26), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n484), .A2(new_n496), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n639), .A2(KEYINPUT26), .A3(new_n632), .A4(new_n634), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n639), .A2(new_n632), .A3(new_n588), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n562), .B1(new_n581), .B2(new_n586), .ZN(new_n643));
  INV_X1    g0443(.A(new_n596), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(new_n644), .A3(KEYINPUT85), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT85), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n592), .B2(new_n596), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n624), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(KEYINPUT86), .B1(new_n642), .B2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n624), .ZN(new_n650));
  AOI21_X1  g0450(.A(KEYINPUT85), .B1(new_n643), .B2(new_n644), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n592), .A2(new_n646), .A3(new_n596), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT86), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n653), .A2(new_n508), .A3(new_n654), .A4(new_n588), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n641), .A2(new_n649), .A3(new_n639), .A4(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n459), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n406), .A2(new_n414), .ZN(new_n658));
  INV_X1    g0458(.A(new_n349), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n313), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n658), .B1(new_n660), .B2(new_n308), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n393), .A2(new_n394), .ZN(new_n662));
  OAI21_X1  g0462(.A(KEYINPUT18), .B1(new_n412), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n389), .B1(new_n390), .B2(new_n270), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n381), .A2(new_n398), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  OAI22_X1  g0466(.A1(new_n661), .A2(new_n666), .B1(new_n451), .B2(new_n452), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n438), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n657), .A2(new_n669), .ZN(G369));
  NAND3_X1  g0470(.A1(new_n224), .A2(new_n206), .A3(G13), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(G213), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G343), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(new_n626), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n624), .B(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(new_n628), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(G330), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n643), .A2(new_n644), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n682), .A2(new_n587), .ZN(new_n683));
  INV_X1    g0483(.A(new_n676), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n643), .A2(new_n684), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n683), .A2(new_n685), .B1(new_n597), .B2(new_n684), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n681), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n650), .A2(new_n684), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n683), .A2(new_n688), .A3(new_n685), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n645), .A2(new_n647), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n689), .B1(new_n690), .B2(new_n684), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n687), .A2(new_n691), .ZN(G399));
  INV_X1    g0492(.A(new_n219), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(G41), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n472), .A2(G116), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G1), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n229), .B2(new_n695), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT87), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n508), .A2(new_n629), .A3(new_n588), .A4(new_n676), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n607), .A2(G179), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n493), .A2(new_n555), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n703), .A2(KEYINPUT30), .A3(new_n542), .A4(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT30), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n542), .A2(new_n493), .A3(new_n555), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n706), .B1(new_n707), .B2(new_n702), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n493), .A2(new_n555), .A3(G179), .ZN(new_n709));
  INV_X1    g0509(.A(new_n607), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(new_n522), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n705), .A2(new_n708), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n684), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(KEYINPUT31), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT31), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n712), .A2(new_n715), .A3(new_n684), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n701), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n700), .B1(new_n718), .B2(G330), .ZN(new_n719));
  INV_X1    g0519(.A(G330), .ZN(new_n720));
  AOI211_X1 g0520(.A(KEYINPUT87), .B(new_n720), .C1(new_n701), .C2(new_n717), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n653), .A2(new_n508), .A3(new_n588), .ZN(new_n723));
  AOI22_X1  g0523(.A1(KEYINPUT86), .A2(new_n723), .B1(new_n638), .B2(new_n640), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n655), .A2(new_n639), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n684), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(KEYINPUT88), .B1(new_n726), .B2(KEYINPUT29), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n656), .A2(new_n676), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT88), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT29), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n638), .A2(new_n640), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n597), .A2(new_n624), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n639), .B1(new_n642), .B2(new_n734), .ZN(new_n735));
  OAI211_X1 g0535(.A(KEYINPUT29), .B(new_n676), .C1(new_n733), .C2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n722), .B1(new_n732), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n699), .B1(new_n737), .B2(G1), .ZN(G364));
  INV_X1    g0538(.A(new_n681), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n224), .A2(G13), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G45), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n742), .A2(new_n694), .A3(new_n206), .ZN(new_n743));
  OR2_X1    g0543(.A1(new_n743), .A2(KEYINPUT89), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(KEYINPUT89), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n739), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n680), .A2(G330), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G13), .A2(G33), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(new_n679), .B2(new_n628), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n219), .A2(new_n316), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n755), .B1(KEYINPUT90), .B2(G355), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n756), .B1(KEYINPUT90), .B2(G355), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n757), .B1(G116), .B2(new_n219), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n242), .A2(new_n260), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n693), .A2(new_n316), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n229), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n761), .B1(new_n260), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n758), .B1(new_n759), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n225), .B1(G20), .B2(new_n270), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n765), .A2(KEYINPUT91), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(KEYINPUT91), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n753), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n747), .B1(new_n764), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n276), .A2(new_n402), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n376), .A2(G190), .A3(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n276), .A2(G200), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n376), .A2(G190), .A3(new_n774), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n202), .A2(new_n773), .B1(new_n775), .B2(new_n332), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G179), .A2(G200), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n224), .B1(G190), .B2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n776), .B1(G97), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n224), .A2(G190), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n402), .A2(G179), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n784), .A2(KEYINPUT93), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(KEYINPUT93), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n781), .A2(new_n774), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT92), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n788), .A2(new_n789), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n780), .B1(new_n787), .B2(new_n319), .C1(new_n794), .C2(new_n421), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n781), .A2(new_n777), .ZN(new_n796));
  INV_X1    g0596(.A(G159), .ZN(new_n797));
  OR3_X1    g0597(.A1(new_n796), .A2(KEYINPUT32), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n781), .A2(new_n772), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G68), .ZN(new_n801));
  OAI21_X1  g0601(.A(KEYINPUT32), .B1(new_n796), .B2(new_n797), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n782), .A2(G20), .A3(G190), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n384), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n370), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n798), .A2(new_n801), .A3(new_n802), .A4(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n796), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n807), .A2(G329), .B1(new_n779), .B2(G294), .ZN(new_n808));
  XNOR2_X1  g0608(.A(KEYINPUT33), .B(G317), .ZN(new_n809));
  INV_X1    g0609(.A(new_n773), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n800), .A2(new_n809), .B1(G326), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n370), .B1(new_n803), .B2(new_n605), .ZN(new_n812));
  INV_X1    g0612(.A(new_n775), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n812), .B1(new_n813), .B2(G322), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n808), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G311), .ZN(new_n816));
  INV_X1    g0616(.A(G283), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n794), .A2(new_n816), .B1(new_n817), .B2(new_n787), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n795), .A2(new_n806), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n771), .B1(new_n819), .B2(new_n768), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n748), .A2(new_n750), .B1(new_n754), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(G396));
  NAND2_X1  g0622(.A1(new_n349), .A2(KEYINPUT96), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT96), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n347), .B(new_n824), .C1(new_n348), .C2(new_n342), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n826), .A2(new_n344), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n656), .A2(new_n676), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n684), .B1(new_n348), .B2(new_n342), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n823), .A2(new_n344), .A3(new_n829), .A4(new_n825), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n659), .A2(new_n684), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n828), .B1(new_n726), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n722), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT97), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n747), .B1(new_n833), .B2(new_n834), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n768), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n752), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n747), .B1(G77), .B2(new_n840), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT94), .Z(new_n842));
  INV_X1    g0642(.A(new_n787), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(G87), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n610), .B2(new_n794), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n370), .B1(new_n319), .B2(new_n803), .C1(new_n778), .C2(new_n253), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n800), .A2(G283), .B1(G303), .B2(new_n810), .ZN(new_n847));
  INV_X1    g0647(.A(G294), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n847), .B1(new_n848), .B2(new_n775), .C1(new_n816), .C2(new_n796), .ZN(new_n849));
  NOR3_X1   g0649(.A1(new_n845), .A2(new_n846), .A3(new_n849), .ZN(new_n850));
  AOI22_X1  g0650(.A1(G143), .A2(new_n813), .B1(new_n810), .B2(G137), .ZN(new_n851));
  INV_X1    g0651(.A(G150), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n851), .B1(new_n852), .B2(new_n799), .C1(new_n794), .C2(new_n797), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(KEYINPUT34), .ZN(new_n854));
  INV_X1    g0654(.A(new_n803), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n370), .B1(new_n855), .B2(G50), .ZN(new_n856));
  INV_X1    g0656(.A(G132), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n856), .B1(new_n778), .B2(new_n332), .C1(new_n796), .C2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(new_n843), .B2(G68), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n850), .B1(new_n854), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(KEYINPUT95), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n768), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n860), .A2(KEYINPUT95), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n842), .B1(new_n752), .B2(new_n832), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n838), .A2(new_n864), .ZN(G384));
  INV_X1    g0665(.A(new_n535), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n610), .B(new_n227), .C1(KEYINPUT35), .C2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(KEYINPUT35), .B2(new_n866), .ZN(new_n868));
  XOR2_X1   g0668(.A(new_n868), .B(KEYINPUT36), .Z(new_n869));
  OR3_X1    g0669(.A1(new_n229), .A2(new_n421), .A3(new_n362), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n202), .A2(G68), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n871), .B(KEYINPUT98), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n206), .B(G13), .C1(new_n870), .C2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n459), .A2(new_n736), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n668), .B1(new_n732), .B2(new_n875), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n876), .B(KEYINPUT103), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n381), .A2(new_n664), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n381), .A2(new_n675), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n412), .A2(new_n413), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT37), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT37), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n396), .A2(new_n879), .A3(new_n880), .A4(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(KEYINPUT101), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n406), .A2(new_n663), .A3(new_n414), .A4(new_n665), .ZN(new_n887));
  INV_X1    g0687(.A(new_n879), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT102), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT101), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n882), .A2(new_n891), .A3(new_n884), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT102), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n887), .A2(new_n893), .A3(new_n888), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n886), .A2(new_n890), .A3(new_n892), .A4(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT38), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT39), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n366), .B1(new_n369), .B2(new_n373), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n410), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n408), .A2(new_n900), .B1(new_n354), .B2(new_n356), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n901), .A2(new_n674), .ZN(new_n902));
  OAI22_X1  g0702(.A1(new_n381), .A2(new_n405), .B1(new_n901), .B2(new_n662), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT37), .B1(new_n903), .B2(new_n902), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n415), .A2(new_n902), .B1(new_n904), .B2(new_n884), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT38), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n897), .A2(new_n898), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n415), .A2(new_n902), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n904), .A2(new_n884), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT99), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n908), .A2(new_n909), .A3(new_n910), .A4(KEYINPUT38), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(KEYINPUT38), .B2(new_n905), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n910), .B1(new_n905), .B2(KEYINPUT38), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT39), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n907), .A2(new_n914), .A3(KEYINPUT100), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n308), .A2(new_n684), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT100), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n917), .B(KEYINPUT39), .C1(new_n912), .C2(new_n913), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n915), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n666), .A2(new_n674), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n676), .B1(new_n305), .B2(new_n306), .ZN(new_n923));
  AOI211_X1 g0723(.A(new_n923), .B(new_n312), .C1(new_n278), .C2(new_n307), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n278), .A2(new_n923), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n912), .A2(new_n913), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n826), .A2(new_n684), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  AOI211_X1 g0730(.A(new_n927), .B(new_n928), .C1(new_n828), .C2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n922), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n877), .B(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT40), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n718), .A2(new_n926), .A3(new_n832), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n935), .B1(new_n928), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n897), .A2(new_n906), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n832), .B1(new_n924), .B2(new_n925), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n701), .B2(new_n717), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n938), .A2(KEYINPUT40), .A3(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n937), .A2(new_n941), .A3(G330), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n720), .B1(new_n701), .B2(new_n717), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n459), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT104), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n937), .A2(new_n941), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n459), .A2(new_n718), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n934), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n206), .B2(new_n740), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n934), .A2(new_n949), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n874), .B1(new_n951), .B2(new_n952), .ZN(G367));
  OR3_X1    g0753(.A1(new_n639), .A2(new_n505), .A3(new_n676), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n508), .B1(new_n505), .B2(new_n676), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n954), .A2(new_n955), .A3(KEYINPUT105), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(KEYINPUT105), .B2(new_n954), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n753), .ZN(new_n958));
  AOI22_X1  g0758(.A1(G150), .A2(new_n813), .B1(new_n810), .B2(G143), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n281), .B2(new_n778), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n370), .B1(new_n855), .B2(G58), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n783), .B2(new_n421), .ZN(new_n962));
  INV_X1    g0762(.A(G137), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n963), .A2(new_n796), .B1(new_n799), .B2(new_n797), .ZN(new_n964));
  NOR3_X1   g0764(.A1(new_n960), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n202), .B2(new_n794), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n794), .A2(new_n817), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n803), .A2(new_n610), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT46), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n775), .A2(new_n605), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n773), .A2(new_n816), .ZN(new_n971));
  NOR4_X1   g0771(.A1(new_n969), .A2(new_n316), .A3(new_n970), .A4(new_n971), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n807), .A2(G317), .B1(new_n784), .B2(G97), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n800), .A2(G294), .B1(new_n779), .B2(G107), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n966), .B1(new_n967), .B2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n839), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n976), .B2(new_n977), .ZN(new_n979));
  INV_X1    g0779(.A(new_n330), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n769), .B1(new_n219), .B2(new_n980), .C1(new_n761), .C2(new_n238), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n958), .A2(new_n747), .A3(new_n979), .A4(new_n981), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n537), .A2(new_n539), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n544), .B1(new_n983), .B2(new_n676), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n634), .A2(new_n684), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n689), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT42), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT43), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n633), .B1(new_n984), .B2(new_n682), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT106), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n992), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n993), .A2(new_n676), .A3(new_n994), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n989), .A2(new_n990), .A3(new_n957), .A4(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT107), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n957), .B(KEYINPUT43), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n989), .A2(new_n995), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n687), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1001), .B1(new_n1002), .B2(new_n987), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n997), .A2(new_n687), .A3(new_n986), .A4(new_n1000), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n742), .A2(new_n206), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n686), .B1(new_n650), .B2(new_n684), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n689), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(new_n681), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n691), .A2(new_n987), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT44), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n691), .A2(KEYINPUT44), .A3(new_n987), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n689), .B(new_n986), .C1(new_n690), .C2(new_n684), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT45), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1016), .B(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n687), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1015), .A2(new_n1018), .A3(new_n1002), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n737), .B1(new_n1010), .B2(new_n1022), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n694), .B(KEYINPUT41), .Z(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1007), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n982), .B1(new_n1005), .B2(new_n1026), .ZN(G387));
  OAI22_X1  g0827(.A1(new_n778), .A2(new_n817), .B1(new_n848), .B2(new_n803), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n800), .A2(G311), .B1(G317), .B2(new_n813), .ZN(new_n1029));
  INV_X1    g0829(.A(G322), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1029), .B1(new_n1030), .B2(new_n773), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(G303), .B2(new_n793), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1028), .B1(new_n1032), .B2(KEYINPUT48), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT111), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(KEYINPUT48), .B2(new_n1032), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT49), .Z(new_n1036));
  AOI21_X1  g0836(.A(new_n316), .B1(new_n807), .B2(G326), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n610), .B2(new_n783), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n794), .A2(new_n281), .B1(new_n253), .B2(new_n787), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n316), .B1(new_n421), .B2(new_n803), .C1(new_n799), .C2(new_n355), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n202), .A2(new_n775), .B1(new_n773), .B2(new_n797), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n796), .A2(new_n852), .B1(new_n778), .B2(new_n980), .ZN(new_n1043));
  NOR4_X1   g0843(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n768), .B1(new_n1039), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT109), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n260), .B1(new_n281), .B2(new_n421), .C1(new_n696), .C2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(G50), .B1(new_n333), .B2(new_n335), .ZN(new_n1048));
  XOR2_X1   g0848(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n1049));
  OR2_X1    g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1049), .A2(new_n202), .A3(new_n336), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n696), .A2(new_n1046), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n760), .B1(new_n1047), .B2(new_n1053), .C1(new_n235), .C2(new_n260), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1054), .B1(G107), .B2(new_n219), .C1(new_n696), .C2(new_n755), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n746), .B1(new_n1055), .B2(new_n769), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1045), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(new_n686), .B2(new_n753), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1010), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1058), .B1(new_n1007), .B2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n695), .B1(new_n737), .B2(new_n1059), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n737), .B2(new_n1059), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1062), .ZN(G393));
  NAND3_X1  g0863(.A1(new_n1020), .A2(KEYINPUT112), .A3(new_n1021), .ZN(new_n1064));
  OR3_X1    g0864(.A1(new_n1019), .A2(KEYINPUT112), .A3(new_n687), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n1007), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n316), .B1(new_n803), .B2(new_n281), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n807), .B2(G143), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n844), .A2(new_n1069), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n1070), .A2(KEYINPUT113), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(KEYINPUT113), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n852), .A2(new_n773), .B1(new_n775), .B2(new_n797), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT51), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n799), .A2(new_n202), .B1(new_n778), .B2(new_n421), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n793), .B2(new_n336), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1071), .A2(new_n1072), .A3(new_n1074), .A4(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n807), .A2(G322), .B1(new_n779), .B2(G116), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n316), .B1(new_n855), .B2(G283), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(new_n605), .C2(new_n799), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n843), .B2(G107), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G311), .A2(new_n813), .B1(new_n810), .B2(G317), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n793), .A2(G294), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1081), .B(new_n1084), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n839), .B1(new_n1077), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n769), .B1(new_n253), .B2(new_n219), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n245), .B2(new_n760), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n1086), .A2(new_n746), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n753), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1089), .B1(new_n1090), .B2(new_n986), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n737), .A2(new_n1059), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1092), .A2(new_n1065), .A3(new_n1064), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n737), .A2(new_n1059), .A3(new_n1021), .A4(new_n1020), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n694), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1067), .B(new_n1091), .C1(new_n1094), .C2(new_n1096), .ZN(G390));
  AOI21_X1  g0897(.A(new_n729), .B1(new_n728), .B2(new_n730), .ZN(new_n1098));
  AOI211_X1 g0898(.A(KEYINPUT88), .B(KEYINPUT29), .C1(new_n656), .C2(new_n676), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n875), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1100), .A2(new_n669), .A3(new_n944), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(KEYINPUT116), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n676), .B1(new_n733), .B2(new_n735), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n827), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n930), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n926), .B1(new_n943), .B2(new_n832), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n832), .ZN(new_n1108));
  NOR3_X1   g0908(.A1(new_n719), .A2(new_n721), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(KEYINPUT115), .B1(new_n1109), .B2(new_n926), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n718), .A2(G330), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(KEYINPUT87), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n943), .A2(new_n700), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1112), .A2(new_n1113), .A3(new_n832), .A4(new_n926), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT115), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1107), .B1(new_n1110), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n943), .A2(new_n832), .A3(new_n926), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n1109), .B2(new_n926), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n828), .A2(new_n930), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT116), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1100), .A2(new_n1123), .A3(new_n669), .A4(new_n944), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1102), .A2(new_n1122), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n915), .A2(new_n918), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n927), .B1(new_n828), .B2(new_n930), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1126), .B1(new_n1127), .B2(new_n916), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n722), .A2(KEYINPUT115), .A3(new_n832), .A4(new_n926), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1105), .A2(new_n926), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n916), .B1(new_n897), .B2(new_n906), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1128), .A2(new_n1131), .A3(new_n1134), .ZN(new_n1135));
  AND2_X1   g0935(.A1(new_n1128), .A2(new_n1134), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1135), .B1(new_n1136), .B2(new_n1118), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n695), .B1(new_n1125), .B2(new_n1137), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n1128), .A2(new_n1131), .A3(new_n1134), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1118), .B1(new_n1128), .B2(new_n1134), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1141), .A2(new_n1124), .A3(new_n1102), .A4(new_n1122), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1138), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1141), .A2(new_n1007), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n747), .B1(new_n429), .B2(new_n840), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n793), .A2(G97), .B1(G107), .B2(new_n800), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT118), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n316), .B(new_n804), .C1(new_n779), .C2(G77), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n807), .A2(G294), .B1(G116), .B2(new_n813), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1148), .B(new_n1149), .C1(new_n817), .C2(new_n773), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(G68), .B2(new_n843), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n316), .B1(new_n783), .B2(new_n202), .ZN(new_n1152));
  XOR2_X1   g0952(.A(new_n1152), .B(KEYINPUT117), .Z(new_n1153));
  OR3_X1    g0953(.A1(new_n803), .A2(KEYINPUT53), .A3(new_n852), .ZN(new_n1154));
  OAI21_X1  g0954(.A(KEYINPUT53), .B1(new_n803), .B2(new_n852), .ZN(new_n1155));
  INV_X1    g0955(.A(G125), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1154), .B(new_n1155), .C1(new_n1156), .C2(new_n796), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n779), .A2(G159), .B1(new_n813), .B2(G132), .ZN(new_n1158));
  INV_X1    g0958(.A(G128), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1158), .B1(new_n1159), .B2(new_n773), .C1(new_n963), .C2(new_n799), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(KEYINPUT54), .B(G143), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1157), .B(new_n1160), .C1(new_n793), .C2(new_n1162), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1147), .A2(new_n1151), .B1(new_n1153), .B2(new_n1163), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n1164), .A2(KEYINPUT119), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n839), .B1(new_n1164), .B2(KEYINPUT119), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1145), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1126), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1167), .B1(new_n1168), .B2(new_n752), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n1144), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1143), .A2(new_n1170), .ZN(G378));
  INV_X1    g0971(.A(KEYINPUT123), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n674), .B1(new_n443), .B2(new_n439), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n456), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n453), .A2(new_n1173), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1177), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n942), .A2(new_n1181), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1180), .A2(G330), .A3(new_n937), .A4(new_n941), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1184), .A2(new_n922), .A3(new_n932), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1183), .B(new_n1182), .C1(new_n921), .C2(new_n931), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1172), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  AND2_X1   g0987(.A1(new_n1186), .A2(new_n1172), .ZN(new_n1188));
  OAI21_X1  g0988(.A(KEYINPUT57), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1102), .A2(new_n1124), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n1141), .B2(new_n1122), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n694), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1124), .B(new_n1102), .C1(new_n1137), .C2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1195));
  AOI21_X1  g0995(.A(KEYINPUT57), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  OR2_X1    g0996(.A1(new_n1192), .A2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n747), .B1(G50), .B2(new_n840), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n316), .A2(G41), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(G33), .A2(G41), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1199), .A2(G50), .A3(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n783), .A2(new_n332), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1199), .B1(new_n421), .B2(new_n803), .C1(new_n778), .C2(new_n281), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1202), .B(new_n1203), .C1(G283), .C2(new_n807), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n319), .A2(new_n775), .B1(new_n773), .B2(new_n610), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(G97), .B2(new_n800), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1204), .B(new_n1206), .C1(new_n980), .C2(new_n794), .ZN(new_n1207));
  XOR2_X1   g1007(.A(new_n1207), .B(KEYINPUT58), .Z(new_n1208));
  AOI22_X1  g1008(.A1(new_n793), .A2(G137), .B1(G132), .B2(new_n800), .ZN(new_n1209));
  XOR2_X1   g1009(.A(new_n1209), .B(KEYINPUT120), .Z(new_n1210));
  NOR2_X1   g1010(.A1(new_n773), .A2(new_n1156), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n775), .A2(new_n1159), .B1(new_n803), .B2(new_n1161), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(G150), .C2(new_n779), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1210), .A2(new_n1213), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1214), .A2(KEYINPUT59), .ZN(new_n1215));
  INV_X1    g1015(.A(G124), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1200), .B1(new_n796), .B2(new_n1216), .C1(new_n797), .C2(new_n783), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n1214), .B2(KEYINPUT59), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1201), .B(new_n1208), .C1(new_n1215), .C2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT121), .ZN(new_n1220));
  OR2_X1    g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n839), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1198), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n1181), .B2(new_n752), .ZN(new_n1224));
  XOR2_X1   g1024(.A(new_n1224), .B(KEYINPUT122), .Z(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n1195), .B2(new_n1007), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1197), .A2(new_n1226), .ZN(G375));
  OAI22_X1  g1027(.A1(new_n796), .A2(new_n1159), .B1(new_n857), .B2(new_n773), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n370), .B(new_n1202), .C1(G159), .C2(new_n855), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1229), .B1(new_n963), .B2(new_n775), .C1(new_n799), .C2(new_n1161), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n1228), .B(new_n1230), .C1(G50), .C2(new_n779), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n793), .A2(G150), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n370), .B1(new_n253), .B2(new_n803), .C1(new_n778), .C2(new_n980), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n796), .A2(new_n605), .B1(new_n817), .B2(new_n775), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n799), .A2(new_n610), .B1(new_n848), .B2(new_n773), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n843), .A2(G77), .B1(G107), .B2(new_n793), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1231), .A2(new_n1232), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n747), .B1(G68), .B2(new_n840), .C1(new_n1238), .C2(new_n839), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1239), .B(KEYINPUT124), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(new_n751), .B2(new_n927), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1122), .B2(new_n1007), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1125), .A2(new_n1025), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1122), .B1(new_n1102), .B2(new_n1124), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1242), .B1(new_n1243), .B2(new_n1244), .ZN(G381));
  NAND2_X1  g1045(.A1(new_n1144), .A2(new_n1169), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(new_n1138), .B2(new_n1142), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1197), .A2(new_n1247), .A3(new_n1226), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(G393), .A2(G396), .ZN(new_n1249));
  INV_X1    g1049(.A(G384), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1067), .A2(new_n1091), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1096), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1251), .B1(new_n1252), .B2(new_n1093), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1249), .A2(new_n1250), .A3(new_n1253), .ZN(new_n1254));
  OR4_X1    g1054(.A1(G387), .A2(new_n1248), .A3(G381), .A4(new_n1254), .ZN(G407));
  OAI211_X1 g1055(.A(G407), .B(G213), .C1(G343), .C2(new_n1248), .ZN(G409));
  AOI21_X1  g1056(.A(new_n1244), .B1(KEYINPUT60), .B2(new_n1125), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1123), .B1(new_n876), .B2(new_n944), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1124), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1193), .B(KEYINPUT60), .C1(new_n1258), .C2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n694), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1242), .B1(new_n1257), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1250), .ZN(new_n1263));
  OAI211_X1 g1063(.A(G384), .B(new_n1242), .C1(new_n1257), .C2(new_n1261), .ZN(new_n1264));
  INV_X1    g1064(.A(G213), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1265), .A2(G343), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(G2897), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1263), .A2(new_n1264), .A3(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1267), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  OAI211_X1 g1070(.A(G378), .B(new_n1226), .C1(new_n1192), .C2(new_n1196), .ZN(new_n1271));
  AND3_X1   g1071(.A1(new_n1194), .A2(new_n1025), .A3(new_n1195), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1007), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1224), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1247), .B1(new_n1272), .B2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1266), .B1(new_n1271), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT61), .B1(new_n1270), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT62), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1125), .A2(KEYINPUT60), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1190), .A2(new_n1193), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1282), .A2(new_n694), .A3(new_n1260), .ZN(new_n1283));
  AOI21_X1  g1083(.A(G384), .B1(new_n1283), .B2(new_n1242), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1264), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1276), .A2(new_n1279), .A3(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1271), .A2(new_n1275), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1266), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1288), .A2(new_n1286), .A3(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(KEYINPUT62), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1278), .A2(new_n1287), .A3(new_n1291), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(G393), .B(G396), .ZN(new_n1293));
  AND2_X1   g1093(.A1(G387), .A2(new_n1253), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(G387), .A2(new_n1253), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1293), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n821), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1249), .A2(new_n1297), .ZN(new_n1298));
  OAI211_X1 g1098(.A(G390), .B(new_n982), .C1(new_n1026), .C2(new_n1005), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(G387), .A2(new_n1253), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1298), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1296), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT126), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1292), .A2(new_n1307), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1263), .A2(KEYINPUT63), .A3(new_n1264), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1276), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1302), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(KEYINPUT63), .B1(new_n1276), .B2(new_n1286), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(KEYINPUT125), .B1(new_n1314), .B2(new_n1278), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT63), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1290), .A2(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1302), .B1(new_n1276), .B2(new_n1309), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT125), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT61), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1267), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1322), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1263), .A2(new_n1264), .A3(new_n1267), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1321), .B1(new_n1325), .B2(new_n1276), .ZN(new_n1326));
  NOR3_X1   g1126(.A1(new_n1319), .A2(new_n1320), .A3(new_n1326), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1308), .B1(new_n1315), .B2(new_n1327), .ZN(G405));
  INV_X1    g1128(.A(KEYINPUT127), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1306), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1329), .B1(new_n1330), .B2(new_n1304), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1305), .A2(KEYINPUT127), .A3(new_n1306), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(G375), .A2(new_n1247), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(new_n1271), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1334), .A2(new_n1286), .ZN(new_n1335));
  OAI211_X1 g1135(.A(new_n1333), .B(new_n1271), .C1(new_n1284), .C2(new_n1285), .ZN(new_n1336));
  NAND4_X1  g1136(.A1(new_n1331), .A2(new_n1332), .A3(new_n1335), .A4(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1338), .A2(new_n1329), .A3(new_n1307), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1337), .A2(new_n1339), .ZN(G402));
endmodule


