//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 0 0 0 0 1 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n546, new_n547, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n560, new_n564, new_n565, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n598, new_n601, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1163, new_n1164, new_n1165, new_n1166;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  XOR2_X1   g012(.A(KEYINPUT66), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT67), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  OR4_X1    g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  AOI21_X1  g035(.A(KEYINPUT70), .B1(new_n460), .B2(KEYINPUT3), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT69), .B(KEYINPUT3), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n461), .B1(new_n462), .B2(new_n460), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT69), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(KEYINPUT69), .ZN(new_n467));
  OAI211_X1 g042(.A(KEYINPUT70), .B(G2104), .C1(new_n465), .C2(new_n467), .ZN(new_n468));
  AOI21_X1  g043(.A(G2105), .B1(new_n463), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G137), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n466), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n466), .A2(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT68), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n471), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  AND2_X1   g054(.A1(G113), .A2(G2104), .ZN(new_n480));
  OAI21_X1  g055(.A(G2105), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n460), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G101), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT71), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n470), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G160));
  OAI21_X1  g061(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G112), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(new_n488), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G2105), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n490), .B1(new_n463), .B2(new_n468), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G124), .ZN(new_n492));
  XNOR2_X1  g067(.A(new_n492), .B(KEYINPUT72), .ZN(new_n493));
  AOI211_X1 g068(.A(new_n489), .B(new_n493), .C1(G136), .C2(new_n469), .ZN(G162));
  NAND2_X1  g069(.A1(new_n475), .A2(new_n478), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n490), .A2(G138), .ZN(new_n496));
  OR2_X1    g071(.A1(KEYINPUT73), .A2(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT73), .A2(KEYINPUT4), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n496), .B1(new_n463), .B2(new_n468), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(G114), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n504), .B1(new_n505), .B2(G2105), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n506), .B1(new_n491), .B2(G126), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G50), .ZN(new_n512));
  XNOR2_X1  g087(.A(new_n512), .B(KEYINPUT74), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT5), .B(G543), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n510), .A2(new_n514), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n515), .A2(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n513), .A2(new_n519), .ZN(G166));
  NAND2_X1  g095(.A1(new_n510), .A2(G543), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT75), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n522), .A2(G51), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT76), .B(G89), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n510), .A2(new_n526), .B1(G63), .B2(G651), .ZN(new_n527));
  XOR2_X1   g102(.A(KEYINPUT5), .B(G543), .Z(new_n528));
  OAI21_X1  g103(.A(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n523), .A2(new_n529), .ZN(G168));
  NAND2_X1  g105(.A1(G77), .A2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G64), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n528), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G651), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n535), .B2(new_n517), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n536), .B1(new_n522), .B2(G52), .ZN(G171));
  NAND2_X1  g112(.A1(new_n522), .A2(G43), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n516), .ZN(new_n540));
  INV_X1    g115(.A(G81), .ZN(new_n541));
  OAI211_X1 g116(.A(new_n538), .B(new_n540), .C1(new_n541), .C2(new_n517), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND4_X1  g122(.A1(G319), .A2(G483), .A3(G661), .A4(new_n547), .ZN(G188));
  XNOR2_X1  g123(.A(new_n514), .B(KEYINPUT77), .ZN(new_n549));
  INV_X1    g124(.A(G65), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AND2_X1   g126(.A1(G78), .A2(G543), .ZN(new_n552));
  OAI21_X1  g127(.A(G651), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(G53), .ZN(new_n554));
  OR3_X1    g129(.A1(new_n521), .A2(KEYINPUT9), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g130(.A(KEYINPUT9), .B1(new_n521), .B2(new_n554), .ZN(new_n556));
  AND2_X1   g131(.A1(new_n510), .A2(new_n514), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n555), .A2(new_n556), .B1(G91), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n553), .A2(new_n558), .ZN(G299));
  NAND2_X1  g134(.A1(new_n522), .A2(G52), .ZN(new_n560));
  OAI211_X1 g135(.A(new_n560), .B(new_n534), .C1(new_n535), .C2(new_n517), .ZN(G301));
  INV_X1    g136(.A(G168), .ZN(G286));
  INV_X1    g137(.A(G166), .ZN(G303));
  NAND2_X1  g138(.A1(new_n557), .A2(G87), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n511), .A2(G49), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT78), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(G288));
  INV_X1    g144(.A(G86), .ZN(new_n570));
  INV_X1    g145(.A(G48), .ZN(new_n571));
  OAI22_X1  g146(.A1(new_n517), .A2(new_n570), .B1(new_n521), .B2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n514), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n573), .A2(new_n516), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G305));
  AOI22_X1  g151(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n577), .A2(new_n516), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT79), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n580), .B1(G85), .B2(new_n557), .ZN(new_n581));
  AOI22_X1  g156(.A1(G47), .A2(new_n522), .B1(new_n578), .B2(new_n579), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n557), .A2(G92), .ZN(new_n585));
  XOR2_X1   g160(.A(new_n585), .B(KEYINPUT10), .Z(new_n586));
  INV_X1    g161(.A(G66), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n549), .A2(new_n587), .ZN(new_n588));
  AND2_X1   g163(.A1(G79), .A2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n522), .A2(G54), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n586), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n584), .B1(new_n593), .B2(G868), .ZN(G284));
  OAI21_X1  g169(.A(new_n584), .B1(new_n593), .B2(G868), .ZN(G321));
  INV_X1    g170(.A(G868), .ZN(new_n596));
  NOR2_X1   g171(.A1(G286), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g172(.A(G299), .B(KEYINPUT80), .Z(new_n598));
  AOI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(new_n596), .ZN(G297));
  AOI21_X1  g174(.A(new_n597), .B1(new_n598), .B2(new_n596), .ZN(G280));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n593), .B1(new_n601), .B2(G860), .ZN(G148));
  NAND2_X1  g177(.A1(new_n542), .A2(new_n596), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n592), .A2(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(new_n596), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g181(.A1(new_n495), .A2(new_n482), .ZN(new_n607));
  XNOR2_X1  g182(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT13), .ZN(new_n610));
  INV_X1    g185(.A(G2100), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n491), .A2(G123), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n469), .A2(G135), .ZN(new_n614));
  OAI21_X1  g189(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT82), .ZN(new_n616));
  INV_X1    g191(.A(G111), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n615), .A2(new_n616), .B1(new_n617), .B2(G2105), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(new_n616), .B2(new_n615), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n613), .A2(new_n614), .A3(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(G2096), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n612), .A2(new_n622), .ZN(G156));
  XNOR2_X1  g198(.A(G2427), .B(G2438), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2430), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT15), .B(G2435), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n627), .A2(KEYINPUT14), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2443), .B(G2446), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G1341), .B(G1348), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G2451), .B(G2454), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT83), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n633), .A2(new_n636), .ZN(new_n638));
  AND3_X1   g213(.A1(new_n637), .A2(G14), .A3(new_n638), .ZN(G401));
  INV_X1    g214(.A(KEYINPUT18), .ZN(new_n640));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  XNOR2_X1  g216(.A(G2067), .B(G2678), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(KEYINPUT17), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n641), .A2(new_n642), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n640), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(new_n611), .ZN(new_n647));
  XOR2_X1   g222(.A(G2072), .B(G2078), .Z(new_n648));
  AOI21_X1  g223(.A(new_n648), .B1(new_n643), .B2(KEYINPUT18), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(new_n621), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(new_n650), .ZN(G227));
  XOR2_X1   g226(.A(G1971), .B(G1976), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT19), .ZN(new_n653));
  XOR2_X1   g228(.A(G1956), .B(G2474), .Z(new_n654));
  XOR2_X1   g229(.A(G1961), .B(G1966), .Z(new_n655));
  AND2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT20), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n654), .A2(new_n655), .ZN(new_n659));
  NOR3_X1   g234(.A1(new_n653), .A2(new_n656), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n660), .B1(new_n653), .B2(new_n659), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1981), .B(G1986), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT84), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n664), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1991), .B(G1996), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G229));
  NOR2_X1   g244(.A1(G29), .A2(G35), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(G162), .B2(G29), .ZN(new_n671));
  INV_X1    g246(.A(G2090), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT97), .B(KEYINPUT29), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(G16), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(G20), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT23), .Z(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(G299), .B2(G16), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(G1956), .Z(new_n680));
  INV_X1    g255(.A(G2078), .ZN(new_n681));
  INV_X1    g256(.A(G29), .ZN(new_n682));
  NOR2_X1   g257(.A1(G164), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(G27), .B2(new_n682), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n680), .B1(new_n681), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(G5), .A2(G16), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(G171), .B2(G16), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT96), .ZN(new_n688));
  OAI221_X1 g263(.A(new_n685), .B1(new_n681), .B2(new_n684), .C1(new_n688), .C2(G1961), .ZN(new_n689));
  INV_X1    g264(.A(G19), .ZN(new_n690));
  OR3_X1    g265(.A1(new_n690), .A2(KEYINPUT91), .A3(G16), .ZN(new_n691));
  OAI21_X1  g266(.A(KEYINPUT91), .B1(new_n690), .B2(G16), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n691), .B(new_n692), .C1(new_n543), .C2(new_n676), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1341), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT90), .B(G1348), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT89), .ZN(new_n696));
  NOR2_X1   g271(.A1(G4), .A2(G16), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT88), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(new_n592), .B2(new_n676), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n694), .B1(new_n696), .B2(new_n699), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n699), .A2(new_n696), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n688), .A2(G1961), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n676), .A2(G21), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G168), .B2(new_n676), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(G1966), .ZN(new_n705));
  INV_X1    g280(.A(G28), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n706), .A2(KEYINPUT30), .ZN(new_n707));
  AOI21_X1  g282(.A(G29), .B1(new_n706), .B2(KEYINPUT30), .ZN(new_n708));
  OR2_X1    g283(.A1(KEYINPUT31), .A2(G11), .ZN(new_n709));
  NAND2_X1  g284(.A1(KEYINPUT31), .A2(G11), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n707), .A2(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n620), .B2(new_n682), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n705), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g288(.A1(new_n700), .A2(new_n701), .A3(new_n702), .A4(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n689), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT24), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n682), .B1(new_n716), .B2(G34), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(KEYINPUT95), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n717), .A2(KEYINPUT95), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n716), .B2(G34), .ZN(new_n720));
  AOI22_X1  g295(.A1(G160), .A2(G29), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G2084), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n682), .A2(G26), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT28), .Z(new_n724));
  NAND2_X1  g299(.A1(new_n469), .A2(G140), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n491), .A2(G128), .ZN(new_n726));
  OR2_X1    g301(.A1(G104), .A2(G2105), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n727), .B(G2104), .C1(G116), .C2(new_n490), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT92), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n725), .A2(new_n726), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n724), .B1(new_n730), .B2(G29), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G2067), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT93), .B(KEYINPUT25), .Z(new_n733));
  NAND3_X1  g308(.A1(new_n490), .A2(G103), .A3(G2104), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n495), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n736));
  AND3_X1   g311(.A1(new_n469), .A2(KEYINPUT94), .A3(G139), .ZN(new_n737));
  AOI21_X1  g312(.A(KEYINPUT94), .B1(new_n469), .B2(G139), .ZN(new_n738));
  OAI221_X1 g313(.A(new_n735), .B1(new_n490), .B2(new_n736), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  MUX2_X1   g314(.A(G33), .B(new_n739), .S(G29), .Z(new_n740));
  OAI21_X1  g315(.A(new_n732), .B1(new_n740), .B2(G2072), .ZN(new_n741));
  AOI211_X1 g316(.A(new_n722), .B(new_n741), .C1(G2072), .C2(new_n740), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n682), .A2(G32), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n469), .A2(G141), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n491), .A2(G129), .ZN(new_n745));
  NAND3_X1  g320(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT26), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n746), .A2(new_n747), .ZN(new_n749));
  AOI22_X1  g324(.A1(new_n748), .A2(new_n749), .B1(G105), .B2(new_n482), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n744), .A2(new_n745), .A3(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n743), .B1(new_n752), .B2(new_n682), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT27), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1996), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n675), .A2(new_n715), .A3(new_n742), .A4(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n469), .A2(G131), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT85), .Z(new_n758));
  OR2_X1    g333(.A1(G95), .A2(G2105), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n759), .B(G2104), .C1(G107), .C2(new_n490), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT86), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G119), .B2(new_n491), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n758), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n763), .A2(G29), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G25), .B2(G29), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT35), .B(G1991), .Z(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n676), .A2(G24), .ZN(new_n769));
  INV_X1    g344(.A(G290), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n769), .B1(new_n770), .B2(new_n676), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G1986), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n676), .A2(G23), .ZN(new_n774));
  INV_X1    g349(.A(new_n567), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(new_n676), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT33), .B(G1976), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n676), .A2(G22), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G166), .B2(new_n676), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n778), .B1(new_n780), .B2(G1971), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G1971), .B2(new_n780), .ZN(new_n782));
  NOR2_X1   g357(.A1(G6), .A2(G16), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n575), .B2(G16), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT32), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1981), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n767), .B(new_n773), .C1(new_n788), .C2(KEYINPUT34), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT87), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n788), .A2(KEYINPUT34), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n792), .A2(KEYINPUT36), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(KEYINPUT36), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n756), .B1(new_n793), .B2(new_n794), .ZN(G311));
  INV_X1    g370(.A(G311), .ZN(G150));
  NAND2_X1  g371(.A1(new_n593), .A2(G559), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT38), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n522), .A2(G55), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n800), .A2(new_n516), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n799), .B1(KEYINPUT98), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(KEYINPUT98), .ZN(new_n803));
  INV_X1    g378(.A(G93), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(new_n517), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(new_n543), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n542), .B1(new_n802), .B2(new_n805), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n798), .B(new_n809), .Z(new_n810));
  OR2_X1    g385(.A1(new_n810), .A2(KEYINPUT39), .ZN(new_n811));
  INV_X1    g386(.A(G860), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(KEYINPUT39), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n806), .A2(new_n812), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT37), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n814), .A2(new_n816), .ZN(G145));
  INV_X1    g392(.A(new_n507), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n503), .A2(KEYINPUT99), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT99), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n500), .B(new_n820), .C1(new_n501), .C2(new_n502), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n818), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(new_n730), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(new_n739), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n824), .A2(new_n751), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n751), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n491), .A2(G130), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n490), .A2(G118), .ZN(new_n829));
  OAI21_X1  g404(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(G142), .B2(new_n469), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(new_n609), .ZN(new_n833));
  INV_X1    g408(.A(new_n763), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n827), .A2(new_n836), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n620), .B(new_n485), .Z(new_n838));
  XNOR2_X1  g413(.A(G162), .B(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n825), .A2(new_n835), .A3(new_n826), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n837), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT101), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT100), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n846), .A2(new_n840), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n837), .A2(new_n845), .A3(new_n841), .ZN(new_n848));
  AOI21_X1  g423(.A(G37), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n844), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g426(.A(new_n809), .B(new_n604), .Z(new_n852));
  OR2_X1    g427(.A1(new_n592), .A2(G299), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n592), .A2(G299), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n855), .B(KEYINPUT41), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n857), .B1(new_n859), .B2(new_n852), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n860), .A2(KEYINPUT103), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT102), .ZN(new_n862));
  NAND2_X1  g437(.A1(G290), .A2(new_n567), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(G166), .B(G305), .ZN(new_n865));
  NOR2_X1   g440(.A1(G290), .A2(new_n567), .ZN(new_n866));
  OR4_X1    g441(.A1(new_n862), .A2(new_n864), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n862), .B1(new_n864), .B2(new_n866), .ZN(new_n868));
  INV_X1    g443(.A(new_n866), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n869), .A2(KEYINPUT102), .A3(new_n863), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n868), .A2(new_n870), .A3(new_n865), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n861), .B1(KEYINPUT42), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(KEYINPUT42), .B2(new_n873), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n860), .A2(KEYINPUT103), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n875), .B(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(G868), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(G868), .B2(new_n806), .ZN(G295));
  OAI21_X1  g454(.A(new_n878), .B1(G868), .B2(new_n806), .ZN(G331));
  INV_X1    g455(.A(KEYINPUT44), .ZN(new_n881));
  NAND2_X1  g456(.A1(G301), .A2(KEYINPUT104), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT104), .ZN(new_n883));
  NAND2_X1  g458(.A1(G171), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n882), .A2(new_n884), .A3(G168), .ZN(new_n885));
  NAND3_X1  g460(.A1(G286), .A2(KEYINPUT104), .A3(G301), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n809), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n885), .A2(new_n886), .A3(new_n808), .A4(new_n807), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n856), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n887), .A2(KEYINPUT105), .A3(new_n809), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT105), .B1(new_n887), .B2(new_n809), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n889), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n890), .B1(new_n894), .B2(new_n858), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(new_n873), .ZN(new_n896));
  INV_X1    g471(.A(G37), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n895), .A2(new_n873), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n898), .A2(new_n899), .A3(KEYINPUT43), .ZN(new_n900));
  AOI21_X1  g475(.A(G37), .B1(new_n895), .B2(new_n873), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT105), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n888), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n891), .ZN(new_n904));
  INV_X1    g479(.A(new_n889), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n905), .A2(new_n855), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n888), .A2(new_n889), .ZN(new_n907));
  AOI22_X1  g482(.A1(new_n904), .A2(new_n906), .B1(new_n858), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT106), .B1(new_n908), .B2(new_n873), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT106), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n858), .A2(new_n907), .ZN(new_n911));
  AOI211_X1 g486(.A(new_n855), .B(new_n905), .C1(new_n903), .C2(new_n891), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n910), .B(new_n872), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n901), .A2(new_n909), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT43), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n900), .B1(new_n915), .B2(KEYINPUT107), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT107), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n914), .A2(new_n917), .A3(KEYINPUT43), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n881), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  OR2_X1    g494(.A1(new_n914), .A2(KEYINPUT43), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT43), .B1(new_n898), .B2(new_n899), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(new_n881), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT108), .B1(new_n919), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT108), .ZN(new_n925));
  INV_X1    g500(.A(new_n918), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n917), .B1(new_n914), .B2(KEYINPUT43), .ZN(new_n927));
  NOR3_X1   g502(.A1(new_n926), .A2(new_n927), .A3(new_n900), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n925), .B(new_n922), .C1(new_n928), .C2(new_n881), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n924), .A2(new_n929), .ZN(G397));
  INV_X1    g505(.A(KEYINPUT45), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(new_n822), .B2(G1384), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n470), .A2(new_n481), .A3(G40), .A4(new_n484), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n936), .A2(G1986), .A3(G290), .ZN(new_n937));
  OR2_X1    g512(.A1(new_n937), .A2(KEYINPUT48), .ZN(new_n938));
  INV_X1    g513(.A(new_n936), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n763), .B(new_n766), .ZN(new_n940));
  XOR2_X1   g515(.A(new_n730), .B(G2067), .Z(new_n941));
  INV_X1    g516(.A(G1996), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n751), .B(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n939), .B1(new_n940), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n938), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n946), .B1(KEYINPUT48), .B2(new_n937), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n936), .A2(G1996), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(KEYINPUT46), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n936), .B1(new_n752), .B2(new_n941), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n951), .B(KEYINPUT47), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n763), .A2(new_n766), .ZN(new_n953));
  OAI22_X1  g528(.A1(new_n953), .A2(new_n944), .B1(G2067), .B2(new_n730), .ZN(new_n954));
  AOI211_X1 g529(.A(new_n947), .B(new_n952), .C1(new_n939), .C2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT51), .ZN(new_n956));
  INV_X1    g531(.A(G1966), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n932), .A2(KEYINPUT115), .A3(new_n935), .ZN(new_n958));
  AOI21_X1  g533(.A(G1384), .B1(new_n503), .B2(new_n507), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT45), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT116), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n960), .B(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n958), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT115), .B1(new_n932), .B2(new_n935), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n957), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G2084), .ZN(new_n966));
  INV_X1    g541(.A(G1384), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n508), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n968), .A2(KEYINPUT111), .A3(KEYINPUT50), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT50), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n970), .B1(new_n959), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n934), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT110), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n819), .A2(new_n821), .ZN(new_n975));
  AOI21_X1  g550(.A(G1384), .B1(new_n975), .B2(new_n507), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n974), .B1(new_n976), .B2(new_n971), .ZN(new_n977));
  NOR4_X1   g552(.A1(new_n822), .A2(KEYINPUT110), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n966), .B(new_n973), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT117), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n496), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT70), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n476), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n466), .A2(KEYINPUT69), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n984), .B1(new_n987), .B2(G2104), .ZN(new_n988));
  AOI211_X1 g563(.A(new_n983), .B(new_n460), .C1(new_n985), .C2(new_n986), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n982), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT4), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n820), .B1(new_n991), .B2(new_n500), .ZN(new_n992));
  INV_X1    g567(.A(new_n821), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n507), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n994), .A2(new_n971), .A3(new_n967), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT110), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n976), .A2(new_n974), .A3(new_n971), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n998), .A2(KEYINPUT117), .A3(new_n966), .A4(new_n973), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n965), .A2(new_n981), .A3(G168), .A4(new_n999), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n1000), .A2(G8), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n965), .A2(new_n981), .A3(new_n999), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(G286), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n956), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1000), .A2(G8), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1005), .A2(KEYINPUT51), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT62), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1003), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT51), .B1(new_n1008), .B2(new_n1005), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT62), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1001), .A2(new_n956), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G8), .ZN(new_n1013));
  NOR2_X1   g588(.A1(G166), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(KEYINPUT112), .A2(KEYINPUT55), .ZN(new_n1015));
  AND2_X1   g590(.A1(KEYINPUT112), .A2(KEYINPUT55), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1017), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT50), .B1(new_n822), .B2(G1384), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n934), .B1(new_n959), .B2(new_n971), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1019), .A2(new_n672), .A3(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n935), .B1(new_n959), .B2(KEYINPUT45), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1022), .B1(new_n976), .B2(KEYINPUT45), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1021), .B1(new_n1023), .B2(G1971), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1018), .B1(new_n1024), .B2(G8), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n994), .A2(new_n967), .A3(new_n935), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n775), .A2(G1976), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1026), .A2(G8), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT52), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1013), .B1(new_n976), .B2(new_n935), .ZN(new_n1030));
  INV_X1    g605(.A(G1976), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT52), .B1(G288), .B2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1030), .A2(new_n1027), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(G305), .A2(G1981), .ZN(new_n1034));
  INV_X1    g609(.A(G1981), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n575), .A2(new_n1035), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n1034), .A2(KEYINPUT49), .A3(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT49), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1030), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1029), .A2(new_n1033), .A3(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1025), .A2(new_n1041), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n672), .B(new_n973), .C1(new_n977), .C2(new_n978), .ZN(new_n1043));
  INV_X1    g618(.A(G1971), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n994), .A2(KEYINPUT45), .A3(new_n967), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1044), .B1(new_n1046), .B2(new_n1022), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1043), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1048), .A2(G8), .A3(new_n1018), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1042), .A2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n973), .B1(new_n977), .B2(new_n978), .ZN(new_n1051));
  INV_X1    g626(.A(G1961), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n932), .A2(new_n935), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT115), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(new_n962), .A3(new_n958), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n681), .A2(KEYINPUT53), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1053), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n934), .B1(new_n968), .B2(new_n931), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1045), .A2(new_n681), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT123), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1062), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(G171), .B1(new_n1059), .B2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1050), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1007), .A2(new_n1012), .A3(new_n1068), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n1039), .A2(G1976), .A3(G288), .ZN(new_n1070));
  XOR2_X1   g645(.A(new_n1036), .B(KEYINPUT114), .Z(new_n1071));
  OAI21_X1  g646(.A(new_n1030), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AOI22_X1  g647(.A1(new_n1028), .A2(KEYINPUT52), .B1(new_n1030), .B2(new_n1039), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1073), .A2(KEYINPUT113), .A3(new_n1033), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT113), .B1(new_n1073), .B2(new_n1033), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1072), .B1(new_n1076), .B2(new_n1049), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT118), .ZN(new_n1078));
  NOR2_X1   g653(.A1(G286), .A2(new_n1013), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1042), .A2(new_n1002), .A3(new_n1049), .A4(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT63), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1078), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1013), .B1(new_n1043), .B2(new_n1047), .ZN(new_n1083));
  OAI22_X1  g658(.A1(new_n1074), .A2(new_n1075), .B1(new_n1083), .B2(new_n1018), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1002), .A2(new_n1079), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1049), .A2(KEYINPUT63), .ZN(new_n1086));
  NOR3_X1   g661(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1082), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1080), .A2(new_n1078), .A3(new_n1081), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1077), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1069), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT125), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1045), .A2(KEYINPUT53), .A3(new_n681), .ZN(new_n1094));
  OAI22_X1  g669(.A1(new_n1064), .A2(new_n1065), .B1(new_n1054), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT124), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1096), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1051), .A2(new_n1096), .A3(new_n1052), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1095), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1093), .B1(new_n1100), .B2(G301), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1094), .A2(new_n1054), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT123), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1102), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1099), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1106), .B1(new_n1107), .B2(new_n1097), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1108), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1059), .A2(new_n1066), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1110), .B1(new_n1111), .B2(G301), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1101), .A2(new_n1109), .A3(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1067), .B1(new_n1108), .B2(G171), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1050), .B1(new_n1114), .B2(new_n1110), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1092), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT126), .ZN(new_n1117));
  OR2_X1    g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT57), .ZN(new_n1119));
  OAI21_X1  g694(.A(G299), .B1(KEYINPUT119), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(KEYINPUT119), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1120), .B(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT120), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT56), .B(G2072), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1023), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1126), .B1(new_n1127), .B2(G1956), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1124), .B1(new_n1023), .B2(new_n1125), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1123), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1026), .A2(G2067), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1131), .B1(new_n1051), .B2(new_n695), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1130), .B1(new_n592), .B2(new_n1132), .ZN(new_n1133));
  OR2_X1    g708(.A1(new_n1127), .A2(G1956), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1129), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1134), .A2(new_n1135), .A3(new_n1122), .A4(new_n1126), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1023), .A2(new_n942), .ZN(new_n1138));
  XOR2_X1   g713(.A(KEYINPUT58), .B(G1341), .Z(new_n1139));
  NAND2_X1  g714(.A1(new_n1026), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n542), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT121), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(KEYINPUT59), .ZN(new_n1143));
  XOR2_X1   g718(.A(new_n1143), .B(KEYINPUT122), .Z(new_n1144));
  XNOR2_X1  g719(.A(new_n1141), .B(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1132), .A2(KEYINPUT60), .A3(new_n592), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  OR2_X1    g722(.A1(new_n1132), .A2(KEYINPUT60), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n592), .B1(new_n1132), .B2(KEYINPUT60), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1130), .A2(new_n1136), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT61), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  AOI22_X1  g728(.A1(new_n1116), .A2(new_n1117), .B1(new_n1137), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1091), .B1(new_n1118), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n937), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n939), .A2(G1986), .A3(G290), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  XOR2_X1   g733(.A(new_n1158), .B(KEYINPUT109), .Z(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(new_n945), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n955), .B1(new_n1155), .B2(new_n1160), .ZN(G329));
  assign    G231 = 1'b0;
  OR4_X1    g736(.A1(new_n458), .A2(G229), .A3(G401), .A4(G227), .ZN(new_n1163));
  AOI21_X1  g737(.A(new_n1163), .B1(new_n920), .B2(new_n921), .ZN(new_n1164));
  AND3_X1   g738(.A1(new_n850), .A2(new_n1164), .A3(KEYINPUT127), .ZN(new_n1165));
  AOI21_X1  g739(.A(KEYINPUT127), .B1(new_n850), .B2(new_n1164), .ZN(new_n1166));
  NOR2_X1   g740(.A1(new_n1165), .A2(new_n1166), .ZN(G308));
  NAND2_X1  g741(.A1(new_n850), .A2(new_n1164), .ZN(G225));
endmodule


