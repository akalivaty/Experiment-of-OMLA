//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1 1 0 0 1 0 1 1 0 0 1 1 0 1 0 0 1 1 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(KEYINPUT64), .ZN(new_n203));
  NAND2_X1  g0003(.A1(G1), .A2(G20), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n203), .B1(new_n204), .B2(G13), .ZN(new_n205));
  INV_X1    g0005(.A(G13), .ZN(new_n206));
  NAND4_X1  g0006(.A1(new_n206), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  AOI22_X1  g0010(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G50), .A2(G226), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n213), .B1(G77), .B2(G244), .ZN(new_n214));
  AND2_X1   g0014(.A1(KEYINPUT66), .A2(G68), .ZN(new_n215));
  NOR2_X1   g0015(.A1(KEYINPUT66), .A2(G68), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G238), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G58), .A2(G232), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G97), .A2(G257), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n214), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n204), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(G58), .A2(G68), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT65), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n210), .B(new_n227), .C1(new_n230), .C2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XOR2_X1   g0037(.A(G238), .B(G244), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT69), .B(G226), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT70), .B(G250), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n241), .B(new_n245), .Z(G358));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G107), .B(G116), .Z(new_n250));
  XNOR2_X1  g0050(.A(G87), .B(G97), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(G274), .ZN(new_n254));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT71), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT71), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G41), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G45), .ZN(new_n260));
  AOI211_X1 g0060(.A(G1), .B(new_n254), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT3), .B(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G1698), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G222), .ZN(new_n264));
  INV_X1    g0064(.A(G223), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n262), .B(new_n264), .C1(new_n265), .C2(new_n263), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(G77), .B2(new_n262), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n268), .B(KEYINPUT72), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n268), .ZN(new_n271));
  INV_X1    g0071(.A(G1), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n272), .B1(G41), .B2(G45), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  AOI211_X1 g0075(.A(new_n261), .B(new_n270), .C1(G226), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G190), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT74), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT10), .ZN(new_n279));
  INV_X1    g0079(.A(G200), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n277), .B(new_n279), .C1(new_n280), .C2(new_n276), .ZN(new_n281));
  INV_X1    g0081(.A(G50), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n229), .B1(new_n231), .B2(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G20), .A2(G33), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n283), .B1(G150), .B2(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT73), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G58), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n289), .A2(KEYINPUT73), .A3(KEYINPUT8), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n229), .A2(G33), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n285), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n228), .ZN(new_n295));
  NOR3_X1   g0095(.A1(new_n206), .A2(new_n229), .A3(G1), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n293), .A2(new_n295), .B1(new_n282), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n295), .B1(new_n272), .B2(G20), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n297), .B1(new_n282), .B2(new_n299), .ZN(new_n300));
  XOR2_X1   g0100(.A(new_n300), .B(KEYINPUT9), .Z(new_n301));
  NOR2_X1   g0101(.A1(new_n281), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n302), .B1(new_n278), .B2(KEYINPUT10), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n278), .A2(KEYINPUT10), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n304), .B1(new_n281), .B2(new_n301), .ZN(new_n305));
  INV_X1    g0105(.A(G179), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n276), .A2(new_n306), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n307), .B(new_n300), .C1(G169), .C2(new_n276), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n303), .A2(new_n305), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G238), .A2(G1698), .ZN(new_n310));
  INV_X1    g0110(.A(G232), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n262), .B(new_n310), .C1(new_n311), .C2(G1698), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(G107), .B2(new_n262), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n313), .A2(new_n269), .ZN(new_n314));
  AOI211_X1 g0114(.A(new_n261), .B(new_n314), .C1(G244), .C2(new_n275), .ZN(new_n315));
  OR2_X1    g0115(.A1(new_n315), .A2(G169), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G20), .A2(G77), .ZN(new_n317));
  INV_X1    g0117(.A(new_n284), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT15), .B(G87), .ZN(new_n319));
  OAI221_X1 g0119(.A(new_n317), .B1(new_n286), .B2(new_n318), .C1(new_n292), .C2(new_n319), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n320), .A2(new_n295), .B1(G77), .B2(new_n298), .ZN(new_n321));
  INV_X1    g0121(.A(new_n296), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n321), .B1(G77), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n315), .A2(new_n306), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n316), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n309), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n275), .A2(G238), .ZN(new_n328));
  INV_X1    g0128(.A(new_n259), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n272), .B(G274), .C1(new_n329), .C2(G45), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G33), .A2(G97), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n311), .A2(G1698), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n262), .B(new_n333), .C1(G226), .C2(G1698), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n269), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT13), .B1(new_n331), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n269), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n334), .A2(new_n332), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT13), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n339), .A2(new_n340), .A3(new_n330), .A4(new_n328), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n336), .A2(new_n341), .A3(KEYINPUT75), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT75), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n343), .B(KEYINPUT13), .C1(new_n331), .C2(new_n335), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n342), .A2(G200), .A3(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n322), .A2(new_n217), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT12), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n346), .B1(KEYINPUT76), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(KEYINPUT76), .B2(new_n347), .ZN(new_n349));
  OAI21_X1  g0149(.A(G68), .B1(new_n349), .B2(new_n298), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n349), .B1(KEYINPUT12), .B2(new_n322), .ZN(new_n351));
  OAI22_X1  g0151(.A1(new_n217), .A2(new_n229), .B1(new_n282), .B2(new_n318), .ZN(new_n352));
  INV_X1    g0152(.A(G77), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n292), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n295), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n355), .B(KEYINPUT11), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n350), .A2(new_n351), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n336), .A2(new_n341), .A3(G190), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n345), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT77), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n345), .A2(new_n358), .A3(KEYINPUT77), .A4(new_n359), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n342), .A2(G169), .A3(new_n344), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(KEYINPUT14), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT14), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n342), .A2(new_n367), .A3(G169), .A4(new_n344), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n336), .A2(new_n341), .A3(G179), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n366), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n357), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n323), .B1(new_n315), .B2(G190), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(new_n280), .B2(new_n315), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n364), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n291), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n299), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n291), .A2(new_n322), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G159), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n318), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n217), .A2(G58), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n232), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n380), .B1(new_n382), .B2(G20), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT7), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n262), .A2(new_n384), .A3(G20), .ZN(new_n385));
  INV_X1    g0185(.A(G33), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT3), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT3), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(G33), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT7), .B1(new_n390), .B2(new_n229), .ZN(new_n391));
  OAI21_X1  g0191(.A(G68), .B1(new_n385), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n383), .A2(KEYINPUT16), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n295), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n384), .B1(new_n262), .B2(G20), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n390), .A2(KEYINPUT7), .A3(new_n229), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT78), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n390), .A2(KEYINPUT78), .A3(KEYINPUT7), .A4(new_n229), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(new_n217), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(KEYINPUT16), .B1(new_n400), .B2(new_n383), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n378), .B1(new_n394), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G33), .A2(G87), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n265), .A2(new_n263), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n262), .B(new_n404), .C1(G226), .C2(new_n263), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n269), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n330), .B1(new_n274), .B2(new_n311), .ZN(new_n407));
  OAI21_X1  g0207(.A(G169), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n405), .A2(new_n403), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n337), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n261), .B1(new_n275), .B2(G232), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(new_n411), .A3(G179), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n402), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT18), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n400), .A2(new_n383), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT16), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n295), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n231), .B1(new_n217), .B2(G58), .ZN(new_n420));
  OAI22_X1  g0220(.A1(new_n420), .A2(new_n229), .B1(new_n379), .B2(new_n318), .ZN(new_n421));
  INV_X1    g0221(.A(G68), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n422), .B1(new_n395), .B2(new_n396), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n419), .B1(new_n424), .B2(KEYINPUT16), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n418), .A2(new_n425), .B1(new_n376), .B2(new_n377), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n280), .B1(new_n410), .B2(new_n411), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n410), .A2(new_n411), .A3(G190), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n426), .A2(KEYINPUT17), .A3(new_n428), .A4(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT17), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n378), .B(new_n429), .C1(new_n394), .C2(new_n401), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n431), .B1(new_n432), .B2(new_n427), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT18), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n402), .A2(new_n434), .A3(new_n413), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n415), .A2(new_n430), .A3(new_n433), .A4(new_n435), .ZN(new_n436));
  XOR2_X1   g0236(.A(new_n436), .B(KEYINPUT79), .Z(new_n437));
  NAND3_X1  g0237(.A1(new_n327), .A2(new_n374), .A3(new_n437), .ZN(new_n438));
  OR2_X1    g0238(.A1(new_n438), .A2(KEYINPUT80), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(KEYINPUT80), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT5), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n256), .A2(new_n258), .A3(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n260), .A2(G1), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT81), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n255), .A2(KEYINPUT5), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT81), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n443), .A2(new_n448), .A3(new_n444), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n446), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(G270), .A3(new_n271), .ZN(new_n451));
  INV_X1    g0251(.A(G303), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n390), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G264), .A2(G1698), .ZN(new_n454));
  INV_X1    g0254(.A(G257), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n262), .B(new_n454), .C1(new_n455), .C2(G1698), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n337), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n268), .A2(new_n254), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n446), .A2(new_n447), .A3(new_n449), .A4(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n451), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G200), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT85), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G33), .A2(G283), .ZN(new_n463));
  INV_X1    g0263(.A(G97), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n463), .B(new_n229), .C1(G33), .C2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G116), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G20), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n465), .A2(new_n295), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n462), .B1(new_n468), .B2(KEYINPUT20), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n469), .B1(KEYINPUT20), .B2(new_n468), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n465), .A2(new_n295), .A3(new_n467), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT20), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n471), .A2(new_n462), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n272), .A2(G33), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n322), .A2(G116), .A3(new_n419), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n296), .A2(new_n466), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n473), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n470), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n451), .A2(new_n457), .A3(G190), .A4(new_n459), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n461), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(G169), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n482), .B1(new_n470), .B2(new_n477), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n460), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT21), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n451), .A2(new_n459), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n487), .A2(G179), .A3(new_n457), .A4(new_n478), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n460), .A2(new_n483), .A3(KEYINPUT21), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n481), .A2(new_n486), .A3(new_n488), .A4(new_n489), .ZN(new_n490));
  XNOR2_X1  g0290(.A(new_n490), .B(KEYINPUT86), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n450), .A2(G257), .A3(new_n271), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n459), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT82), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT4), .ZN(new_n495));
  INV_X1    g0295(.A(G244), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n495), .B1(new_n390), .B2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n262), .A2(KEYINPUT4), .A3(G244), .A4(new_n263), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n497), .A2(new_n498), .A3(new_n463), .ZN(new_n499));
  OAI21_X1  g0299(.A(KEYINPUT4), .B1(new_n390), .B2(new_n223), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G1698), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n269), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT82), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n492), .A2(new_n504), .A3(new_n459), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n494), .A2(G179), .A3(new_n503), .A4(new_n505), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n492), .A2(new_n504), .A3(new_n459), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n504), .B1(new_n492), .B2(new_n459), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n507), .A2(new_n508), .A3(new_n502), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n506), .B1(new_n509), .B2(new_n482), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n398), .A2(G107), .A3(new_n399), .ZN(new_n511));
  INV_X1    g0311(.A(G107), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(KEYINPUT6), .A3(G97), .ZN(new_n513));
  XOR2_X1   g0313(.A(G97), .B(G107), .Z(new_n514));
  OAI21_X1  g0314(.A(new_n513), .B1(new_n514), .B2(KEYINPUT6), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n515), .A2(G20), .B1(G77), .B2(new_n284), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n419), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n322), .A2(new_n419), .A3(new_n474), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n518), .A2(new_n464), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n322), .A2(G97), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n517), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  XNOR2_X1  g0321(.A(new_n521), .B(KEYINPUT83), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n510), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n262), .A2(new_n229), .A3(G87), .ZN(new_n524));
  XNOR2_X1  g0324(.A(new_n524), .B(KEYINPUT22), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n229), .A2(G107), .ZN(new_n526));
  XNOR2_X1  g0326(.A(new_n526), .B(KEYINPUT23), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n229), .A2(G33), .A3(G116), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n525), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT24), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n525), .A2(KEYINPUT24), .A3(new_n527), .A4(new_n528), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n531), .A2(new_n295), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT87), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT25), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n534), .B(new_n535), .C1(new_n322), .C2(G107), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n296), .B(new_n512), .C1(KEYINPUT87), .C2(KEYINPUT25), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n536), .B(new_n537), .C1(new_n534), .C2(new_n535), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n533), .A2(new_n538), .ZN(new_n539));
  OR2_X1    g0339(.A1(new_n518), .A2(new_n512), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n390), .B1(new_n455), .B2(G1698), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(G250), .B2(G1698), .ZN(new_n542));
  INV_X1    g0342(.A(G294), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n542), .B1(new_n386), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n337), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n450), .A2(G264), .A3(new_n271), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n546), .A3(new_n459), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(G200), .ZN(new_n548));
  INV_X1    g0348(.A(G190), .ZN(new_n549));
  OR2_X1    g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n539), .A2(new_n540), .A3(new_n548), .A4(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n494), .A2(new_n503), .A3(new_n505), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G200), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n494), .A2(G190), .A3(new_n503), .A4(new_n505), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(new_n521), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n523), .A2(new_n551), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n533), .A2(new_n540), .A3(new_n538), .ZN(new_n557));
  OR2_X1    g0357(.A1(new_n547), .A2(G179), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n547), .A2(new_n482), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT19), .ZN(new_n561));
  NOR2_X1   g0361(.A1(G97), .A2(G107), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n222), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n332), .A2(new_n229), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n561), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NOR3_X1   g0365(.A1(new_n292), .A2(KEYINPUT19), .A3(new_n464), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n262), .A2(new_n229), .ZN(new_n567));
  OAI22_X1  g0367(.A1(new_n565), .A2(new_n566), .B1(new_n567), .B2(new_n422), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT84), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT84), .ZN(new_n570));
  OAI221_X1 g0370(.A(new_n570), .B1(new_n567), .B2(new_n422), .C1(new_n565), .C2(new_n566), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n571), .A3(new_n295), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n319), .A2(new_n296), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n572), .B(new_n573), .C1(new_n319), .C2(new_n518), .ZN(new_n574));
  NOR2_X1   g0374(.A1(G238), .A2(G1698), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n575), .B1(new_n496), .B2(G1698), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n576), .A2(new_n262), .B1(G33), .B2(G116), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n269), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n444), .A2(G250), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n260), .A2(G1), .A3(G274), .ZN(new_n580));
  NOR3_X1   g0380(.A1(new_n579), .A2(new_n268), .A3(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n306), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n574), .B(new_n583), .C1(G169), .C2(new_n582), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n572), .A2(new_n573), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n518), .A2(new_n222), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n582), .A2(G190), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n587), .B(new_n588), .C1(new_n280), .C2(new_n582), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n560), .A2(new_n584), .A3(new_n589), .ZN(new_n590));
  NOR3_X1   g0390(.A1(new_n491), .A2(new_n556), .A3(new_n590), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n441), .A2(new_n591), .ZN(G372));
  INV_X1    g0392(.A(new_n560), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n486), .A2(new_n488), .A3(new_n489), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n578), .A2(KEYINPUT88), .ZN(new_n596));
  XNOR2_X1  g0396(.A(new_n581), .B(KEYINPUT89), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT88), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(new_n269), .B2(new_n577), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n596), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(G200), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n587), .A2(new_n601), .A3(new_n588), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(new_n482), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n603), .A2(new_n583), .A3(new_n574), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n523), .A2(new_n551), .A3(new_n555), .A4(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT90), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n595), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n553), .A2(new_n554), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n609), .A2(new_n521), .B1(new_n510), .B2(new_n522), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n610), .A2(KEYINPUT90), .A3(new_n551), .A4(new_n605), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n589), .A2(new_n584), .ZN(new_n613));
  OAI21_X1  g0413(.A(KEYINPUT26), .B1(new_n523), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n552), .A2(G169), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n521), .B1(new_n615), .B2(new_n506), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT26), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(new_n617), .A3(new_n605), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n604), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n612), .A2(new_n614), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n441), .A2(new_n621), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n303), .A2(new_n305), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n430), .A2(new_n433), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n364), .A2(new_n326), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n625), .B1(new_n626), .B2(new_n371), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n415), .A2(new_n435), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n623), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n630), .A2(new_n308), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n622), .A2(new_n631), .ZN(G369));
  NOR2_X1   g0432(.A1(new_n206), .A2(G20), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  OR3_X1    g0434(.A1(new_n634), .A2(KEYINPUT27), .A3(G1), .ZN(new_n635));
  OAI21_X1  g0435(.A(KEYINPUT27), .B1(new_n634), .B2(G1), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(G213), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(G343), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n479), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n594), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n642), .B1(new_n491), .B2(new_n641), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(G330), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n560), .A2(new_n639), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n557), .A2(new_n639), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n551), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n647), .B1(new_n649), .B2(new_n560), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n594), .A2(new_n640), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n647), .B1(new_n650), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n651), .A2(new_n654), .ZN(G399));
  INV_X1    g0455(.A(new_n208), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n656), .A2(new_n329), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n563), .A2(G116), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(G1), .A3(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(new_n233), .B2(new_n658), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n661), .B(KEYINPUT28), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n621), .A2(new_n640), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT29), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n589), .A2(new_n584), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n666), .A2(new_n617), .A3(new_n510), .A4(new_n522), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n616), .A2(new_n605), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n667), .B(new_n604), .C1(new_n668), .C2(new_n617), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n606), .A2(new_n595), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n640), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(KEYINPUT29), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n460), .A2(new_n306), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT92), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT30), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n545), .A2(new_n546), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n509), .A2(new_n582), .A3(new_n674), .A4(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n675), .A2(new_n676), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n494), .A2(new_n582), .A3(new_n503), .A4(new_n505), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n685), .A2(new_n674), .A3(new_n681), .A4(new_n679), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n600), .A2(new_n460), .A3(new_n306), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n552), .A2(new_n547), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT91), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n552), .A2(KEYINPUT91), .A3(new_n547), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n688), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OAI211_X1 g0493(.A(KEYINPUT31), .B(new_n639), .C1(new_n687), .C2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT93), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n639), .B1(new_n687), .B2(new_n693), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT31), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n688), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n552), .A2(KEYINPUT91), .A3(new_n547), .ZN(new_n701));
  AOI21_X1  g0501(.A(KEYINPUT91), .B1(new_n552), .B2(new_n547), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(new_n683), .A3(new_n686), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n704), .A2(KEYINPUT93), .A3(KEYINPUT31), .A4(new_n639), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n523), .A2(new_n551), .A3(new_n555), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT86), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n490), .B(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n590), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n706), .A2(new_n708), .A3(new_n709), .A4(new_n640), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n696), .A2(new_n699), .A3(new_n705), .A4(new_n710), .ZN(new_n711));
  AOI22_X1  g0511(.A1(new_n665), .A2(new_n673), .B1(G330), .B2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n662), .B1(new_n712), .B2(G1), .ZN(G364));
  NOR2_X1   g0513(.A1(new_n643), .A2(G330), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT94), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n272), .B1(new_n633), .B2(G45), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n657), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n715), .B(new_n719), .C1(new_n645), .C2(new_n644), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n228), .B1(G20), .B2(new_n482), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n229), .A2(G190), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n280), .A2(G179), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(G283), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n229), .A2(new_n306), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n727), .A2(new_n549), .A3(G200), .ZN(new_n728));
  INV_X1    g0528(.A(G317), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n728), .B1(KEYINPUT33), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(KEYINPUT33), .B2(new_n729), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n727), .A2(G190), .A3(G200), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n262), .B1(new_n733), .B2(G326), .ZN(new_n734));
  NOR2_X1   g0534(.A1(G179), .A2(G200), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G190), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G20), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n731), .B(new_n734), .C1(new_n543), .C2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n229), .A2(new_n549), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n306), .A2(G200), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT95), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n742), .A2(new_n743), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n739), .B1(G322), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n740), .A2(new_n723), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n722), .A2(new_n735), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI22_X1  g0553(.A1(G303), .A2(new_n751), .B1(new_n753), .B2(G329), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n722), .A2(new_n741), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n726), .B(new_n755), .C1(G311), .C2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n751), .A2(G87), .ZN(new_n759));
  OAI221_X1 g0559(.A(new_n759), .B1(new_n282), .B2(new_n732), .C1(new_n353), .C2(new_n756), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT32), .ZN(new_n761));
  XNOR2_X1  g0561(.A(KEYINPUT96), .B(G159), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n761), .B1(new_n763), .B2(new_n752), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n753), .A2(KEYINPUT32), .A3(new_n762), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n760), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n728), .ZN(new_n767));
  INV_X1    g0567(.A(new_n724), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n767), .A2(G68), .B1(new_n768), .B2(G107), .ZN(new_n769));
  OAI211_X1 g0569(.A(new_n766), .B(new_n769), .C1(new_n464), .C2(new_n738), .ZN(new_n770));
  AOI211_X1 g0570(.A(new_n390), .B(new_n770), .C1(G58), .C2(new_n748), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n721), .B1(new_n758), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n234), .A2(new_n260), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n656), .A2(new_n262), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n773), .B(new_n774), .C1(new_n249), .C2(new_n260), .ZN(new_n775));
  INV_X1    g0575(.A(G355), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n208), .A2(new_n262), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n775), .B1(G116), .B2(new_n208), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G13), .A2(G33), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n721), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n719), .B1(new_n778), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n781), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n772), .B(new_n783), .C1(new_n643), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n720), .A2(new_n785), .ZN(G396));
  NAND2_X1  g0586(.A1(new_n323), .A2(new_n639), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n373), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n325), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n326), .A2(new_n640), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n621), .A2(new_n640), .A3(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n619), .B1(new_n608), .B2(new_n611), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n639), .B1(new_n794), .B2(new_n614), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n791), .B(KEYINPUT99), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n793), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n711), .A2(G330), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n797), .B(new_n798), .Z(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(new_n719), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n738), .A2(new_n464), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n390), .B1(new_n747), .B2(new_n543), .ZN(new_n802));
  XNOR2_X1  g0602(.A(KEYINPUT97), .B(G283), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n801), .B(new_n802), .C1(new_n767), .C2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(G311), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n756), .A2(new_n466), .B1(new_n752), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(G303), .B2(new_n733), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n804), .B(new_n807), .C1(new_n512), .C2(new_n750), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n724), .A2(new_n222), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n767), .A2(G150), .B1(new_n733), .B2(G137), .ZN(new_n810));
  INV_X1    g0610(.A(G143), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n810), .B1(new_n756), .B2(new_n763), .C1(new_n747), .C2(new_n811), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n812), .B(KEYINPUT34), .Z(new_n813));
  NOR2_X1   g0613(.A1(new_n738), .A2(new_n289), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n262), .B1(new_n724), .B2(new_n422), .C1(new_n282), .C2(new_n750), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n814), .B(new_n815), .C1(G132), .C2(new_n753), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT98), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n808), .A2(new_n809), .B1(new_n813), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n719), .B1(new_n818), .B2(new_n721), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n721), .A2(new_n779), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n819), .B1(G77), .B2(new_n821), .C1(new_n792), .C2(new_n780), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n800), .A2(new_n822), .ZN(G384));
  INV_X1    g0623(.A(new_n790), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(new_n795), .B2(new_n792), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n358), .A2(new_n640), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(new_n364), .B2(new_n371), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n364), .A2(new_n371), .A3(new_n827), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(KEYINPUT101), .B1(new_n825), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n793), .A2(new_n790), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT101), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n834), .A2(new_n835), .A3(new_n831), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n418), .A2(new_n425), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n837), .A2(new_n378), .A3(new_n428), .A4(new_n429), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n408), .A2(new_n412), .A3(new_n637), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n402), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT37), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n838), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT103), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n838), .A2(new_n840), .A3(KEYINPUT103), .A4(new_n841), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n417), .B1(new_n421), .B2(new_n423), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n393), .A2(new_n847), .A3(new_n295), .ZN(new_n848));
  AND3_X1   g0648(.A1(new_n848), .A2(KEYINPUT102), .A3(new_n378), .ZN(new_n849));
  INV_X1    g0649(.A(new_n839), .ZN(new_n850));
  AOI21_X1  g0650(.A(KEYINPUT102), .B1(new_n848), .B2(new_n378), .ZN(new_n851));
  NOR3_X1   g0651(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n838), .ZN(new_n853));
  OAI21_X1  g0653(.A(KEYINPUT37), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n846), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n637), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n849), .A2(new_n851), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n436), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT38), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n855), .A2(KEYINPUT38), .A3(new_n858), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n833), .A2(new_n836), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n629), .A2(new_n637), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT39), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n838), .A2(new_n840), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n846), .B1(new_n841), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n436), .A2(new_n402), .A3(new_n856), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT104), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n436), .A2(KEYINPUT104), .A3(new_n402), .A4(new_n856), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n869), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n860), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n637), .B1(new_n628), .B2(new_n624), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n876), .A2(new_n857), .B1(new_n846), .B2(new_n854), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT105), .B1(new_n877), .B2(KEYINPUT38), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT105), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n862), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n875), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n867), .B1(new_n866), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n371), .A2(new_n639), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n864), .A2(new_n865), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n831), .A2(new_n792), .ZN(new_n886));
  AOI22_X1  g0686(.A1(KEYINPUT106), .A2(new_n699), .B1(new_n591), .B2(new_n640), .ZN(new_n887));
  INV_X1    g0687(.A(new_n694), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT106), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT31), .B1(new_n704), .B2(new_n639), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n886), .B1(new_n887), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT40), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n877), .A2(KEYINPUT105), .A3(KEYINPUT38), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n862), .A2(new_n879), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n893), .B1(new_n896), .B2(new_n875), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n791), .B1(new_n829), .B2(new_n830), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n710), .B1(new_n890), .B2(new_n889), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n697), .A2(new_n889), .A3(new_n698), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n694), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n863), .B(new_n898), .C1(new_n899), .C2(new_n901), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n892), .A2(new_n897), .B1(new_n902), .B2(new_n893), .ZN(new_n903));
  INV_X1    g0703(.A(new_n674), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n684), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n681), .B1(new_n905), .B2(new_n679), .ZN(new_n906));
  NOR4_X1   g0706(.A1(new_n684), .A2(new_n904), .A3(new_n678), .A4(new_n682), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n640), .B1(new_n908), .B2(new_n703), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT106), .B1(new_n909), .B2(KEYINPUT31), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n910), .A2(new_n694), .A3(new_n710), .A4(new_n900), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n903), .A2(new_n441), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n441), .A2(G330), .A3(new_n911), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n902), .A2(new_n893), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n881), .A2(new_n911), .A3(KEYINPUT40), .A4(new_n898), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n915), .A2(new_n916), .A3(G330), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n912), .B1(new_n914), .B2(new_n918), .ZN(new_n919));
  XOR2_X1   g0719(.A(new_n885), .B(new_n919), .Z(new_n920));
  NAND3_X1  g0720(.A1(new_n441), .A2(new_n665), .A3(new_n673), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n631), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n920), .B(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n272), .B2(new_n633), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n515), .B(KEYINPUT100), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n466), .B1(new_n925), .B2(KEYINPUT35), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n926), .B(new_n230), .C1(KEYINPUT35), .C2(new_n925), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT36), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n381), .A2(G50), .A3(G77), .A4(new_n232), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(G50), .B2(new_n422), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n930), .A2(G1), .A3(new_n206), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n924), .A2(new_n928), .A3(new_n931), .ZN(G367));
  AOI21_X1  g0732(.A(new_n262), .B1(new_n757), .B2(new_n803), .ZN(new_n933));
  OAI221_X1 g0733(.A(new_n933), .B1(new_n512), .B2(new_n738), .C1(new_n543), .C2(new_n728), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n751), .A2(G116), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT109), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT46), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n768), .A2(G97), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n729), .B2(new_n752), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n937), .B1(new_n935), .B2(new_n936), .ZN(new_n942));
  NOR4_X1   g0742(.A1(new_n934), .A2(new_n939), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n943), .B1(new_n452), .B2(new_n747), .C1(new_n805), .C2(new_n732), .ZN(new_n944));
  OAI221_X1 g0744(.A(new_n262), .B1(new_n750), .B2(new_n289), .C1(new_n811), .C2(new_n732), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n737), .A2(G68), .ZN(new_n946));
  INV_X1    g0746(.A(G137), .ZN(new_n947));
  OAI221_X1 g0747(.A(new_n946), .B1(new_n947), .B2(new_n752), .C1(new_n728), .C2(new_n763), .ZN(new_n948));
  AOI211_X1 g0748(.A(new_n945), .B(new_n948), .C1(G77), .C2(new_n768), .ZN(new_n949));
  INV_X1    g0749(.A(G150), .ZN(new_n950));
  OAI221_X1 g0750(.A(new_n949), .B1(new_n282), .B2(new_n756), .C1(new_n950), .C2(new_n747), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n944), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT47), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n245), .A2(new_n774), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n208), .A2(new_n319), .ZN(new_n955));
  NOR3_X1   g0755(.A1(new_n955), .A2(new_n721), .A3(new_n781), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n953), .A2(new_n721), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n639), .B1(new_n585), .B2(new_n586), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n605), .A2(new_n958), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n604), .A2(new_n958), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n957), .B(new_n718), .C1(new_n784), .C2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n610), .B1(new_n521), .B2(new_n640), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n616), .A2(new_n639), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n523), .B1(new_n966), .B2(new_n560), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n640), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n650), .A2(new_n610), .A3(new_n653), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT42), .Z(new_n970));
  AOI22_X1  g0770(.A1(new_n968), .A2(new_n970), .B1(KEYINPUT43), .B2(new_n961), .ZN(new_n971));
  OR3_X1    g0771(.A1(new_n971), .A2(KEYINPUT43), .A3(new_n961), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n971), .B1(KEYINPUT43), .B2(new_n961), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n651), .A2(new_n966), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n974), .B(new_n975), .Z(new_n976));
  XNOR2_X1  g0776(.A(new_n650), .B(new_n653), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n646), .B(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n965), .A2(new_n654), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT45), .Z(new_n980));
  NOR2_X1   g0780(.A1(new_n965), .A2(new_n654), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT44), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n651), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(KEYINPUT108), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n712), .B(new_n978), .C1(new_n983), .C2(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n985), .B1(new_n982), .B2(new_n980), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n712), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  XOR2_X1   g0789(.A(KEYINPUT107), .B(KEYINPUT41), .Z(new_n990));
  XNOR2_X1  g0790(.A(new_n657), .B(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n717), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n962), .B1(new_n976), .B2(new_n992), .ZN(G387));
  OR2_X1    g0793(.A1(new_n712), .A2(new_n978), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n712), .A2(new_n978), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n994), .A2(new_n657), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n978), .A2(new_n717), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n756), .A2(new_n422), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n375), .A2(new_n767), .B1(G150), .B2(new_n753), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n999), .B1(new_n282), .B2(new_n747), .C1(new_n353), .C2(new_n750), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n998), .B(new_n1000), .C1(G159), .C2(new_n733), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n738), .A2(new_n319), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n1001), .A2(new_n262), .A3(new_n940), .A4(new_n1003), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n748), .A2(G317), .B1(G303), .B2(new_n757), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n733), .A2(G322), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1005), .B(new_n1006), .C1(new_n805), .C2(new_n728), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT48), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n737), .A2(new_n803), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1008), .B(new_n1009), .C1(new_n543), .C2(new_n750), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT49), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n768), .A2(G116), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n753), .A2(G326), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1012), .A2(new_n390), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  AND2_X1   g0815(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1004), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n721), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n659), .B(KEYINPUT110), .Z(new_n1019));
  NOR2_X1   g0819(.A1(new_n286), .A2(G50), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT50), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(G68), .A2(G77), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1019), .A2(new_n1021), .A3(new_n260), .A4(new_n1022), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n774), .B(new_n1023), .C1(new_n241), .C2(new_n260), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1024), .B1(G107), .B2(new_n208), .C1(new_n659), .C2(new_n777), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n719), .B1(new_n1025), .B2(new_n782), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1018), .B(new_n1026), .C1(new_n650), .C2(new_n784), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n996), .A2(new_n997), .A3(new_n1027), .ZN(G393));
  AOI21_X1  g0828(.A(new_n719), .B1(new_n966), .B2(new_n781), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n774), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n782), .B1(new_n464), .B2(new_n208), .C1(new_n1030), .C2(new_n252), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n747), .A2(new_n379), .B1(new_n950), .B2(new_n732), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT111), .Z(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT51), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n751), .A2(new_n217), .B1(new_n737), .B2(G77), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1034), .B(new_n1035), .C1(new_n811), .C2(new_n752), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n756), .A2(new_n286), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n262), .B1(new_n728), .B2(new_n282), .ZN(new_n1038));
  NOR4_X1   g0838(.A1(new_n1036), .A2(new_n809), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n747), .A2(new_n805), .B1(new_n729), .B2(new_n732), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT52), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n757), .A2(G294), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n753), .A2(G322), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n728), .A2(new_n452), .B1(new_n724), .B2(new_n512), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n262), .B(new_n1044), .C1(G116), .C2(new_n737), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .A4(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(new_n751), .B2(new_n803), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n721), .B1(new_n1039), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1029), .A2(new_n1031), .A3(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n983), .B(new_n984), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1049), .B1(new_n1050), .B2(new_n716), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT112), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1050), .A2(new_n995), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1053), .B(new_n657), .C1(new_n987), .C2(new_n988), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1054), .ZN(G390));
  OAI211_X1 g0855(.A(G330), .B(new_n796), .C1(new_n899), .C2(new_n901), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n832), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n789), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n790), .B1(new_n671), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n711), .A2(G330), .A3(new_n792), .A4(new_n831), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1057), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n645), .B1(new_n887), .B2(new_n891), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n711), .A2(G330), .A3(new_n792), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n1064), .A2(new_n898), .B1(new_n1065), .B2(new_n832), .ZN(new_n1066));
  OAI21_X1  g0866(.A(KEYINPUT113), .B1(new_n1066), .B2(new_n825), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1065), .A2(new_n832), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n911), .A2(G330), .A3(new_n898), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT113), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1070), .A2(new_n1071), .A3(new_n834), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1063), .B1(new_n1067), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n921), .A2(new_n913), .A3(new_n631), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n867), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n894), .A2(new_n895), .B1(new_n860), .B2(new_n874), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1078), .B1(new_n1079), .B2(KEYINPUT39), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n832), .B1(new_n793), .B2(new_n790), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1080), .B1(new_n1081), .B2(new_n883), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n883), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n881), .B(new_n1083), .C1(new_n1060), .C2(new_n832), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1061), .ZN(new_n1085));
  AND3_X1   g0885(.A1(new_n1082), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1069), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1077), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1082), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n883), .B(new_n1079), .C1(new_n1059), .C2(new_n831), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1083), .B1(new_n825), .B2(new_n832), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1092), .B1(new_n1080), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1091), .B1(new_n1094), .B2(new_n1087), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1074), .A2(new_n1095), .A3(new_n1076), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1090), .A2(new_n1096), .A3(new_n657), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n1069), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n716), .B1(new_n1099), .B2(new_n1091), .ZN(new_n1100));
  INV_X1    g0900(.A(G128), .ZN(new_n1101));
  INV_X1    g0901(.A(G125), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n732), .A2(new_n1101), .B1(new_n752), .B2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n262), .B1(new_n724), .B2(new_n282), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT115), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1103), .B(new_n1105), .C1(G132), .C2(new_n748), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n767), .A2(G137), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n750), .A2(new_n950), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT53), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n1108), .A2(new_n1109), .B1(new_n738), .B2(new_n379), .ZN(new_n1111));
  XOR2_X1   g0911(.A(KEYINPUT54), .B(G143), .Z(new_n1112));
  AOI21_X1  g0912(.A(new_n1111), .B1(new_n757), .B2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1106), .A2(new_n1107), .A3(new_n1110), .A4(new_n1113), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n390), .B1(new_n728), .B2(new_n512), .C1(new_n725), .C2(new_n732), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n747), .A2(new_n466), .B1(new_n353), .B2(new_n738), .ZN(new_n1116));
  XOR2_X1   g0916(.A(new_n1116), .B(KEYINPUT116), .Z(new_n1117));
  AOI211_X1 g0917(.A(new_n1115), .B(new_n1117), .C1(G97), .C2(new_n757), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1118), .B(new_n759), .C1(new_n543), .C2(new_n752), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n724), .A2(new_n422), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1114), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n721), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n718), .B1(new_n375), .B2(new_n821), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT114), .Z(new_n1124));
  OAI211_X1 g0924(.A(new_n1122), .B(new_n1124), .C1(new_n882), .C2(new_n780), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT117), .ZN(new_n1126));
  OR3_X1    g0926(.A1(new_n1100), .A2(KEYINPUT118), .A3(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(KEYINPUT118), .B1(new_n1100), .B2(new_n1126), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1097), .A2(new_n1127), .A3(new_n1128), .ZN(G378));
  INV_X1    g0929(.A(KEYINPUT57), .ZN(new_n1130));
  XOR2_X1   g0930(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1131));
  OR2_X1    g0931(.A1(new_n309), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n309), .A2(new_n1131), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n300), .A2(new_n856), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1132), .A2(new_n300), .A3(new_n856), .A4(new_n1133), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n903), .B2(G330), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n915), .A2(new_n916), .A3(new_n1138), .A4(G330), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n885), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1138), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n917), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n1140), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1146), .A2(new_n865), .A3(new_n884), .A4(new_n864), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n1143), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1075), .B1(new_n1074), .B2(new_n1095), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1130), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1076), .B1(new_n1089), .B2(new_n1073), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT119), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1143), .A2(new_n1147), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n885), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1154), .A2(KEYINPUT119), .A3(new_n1146), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1151), .A2(new_n1153), .A3(KEYINPUT57), .A4(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1150), .A2(new_n1156), .A3(new_n657), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1143), .A2(new_n1147), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n717), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n390), .A2(new_n259), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1160), .B(new_n282), .C1(G33), .C2(G41), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n748), .A2(G128), .B1(new_n751), .B2(new_n1112), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n767), .A2(G132), .B1(new_n733), .B2(G125), .ZN(new_n1163));
  AND2_X1   g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1164), .B1(new_n947), .B2(new_n756), .C1(new_n950), .C2(new_n738), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT59), .ZN(new_n1166));
  AOI211_X1 g0966(.A(G33), .B(G41), .C1(new_n753), .C2(G124), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n724), .B2(new_n763), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1161), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n756), .A2(new_n319), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n728), .A2(new_n464), .B1(new_n724), .B2(new_n289), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1170), .B(new_n1171), .C1(new_n748), .C2(G107), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1160), .B1(G77), .B2(new_n751), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n753), .A2(G283), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1172), .A2(new_n946), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(G116), .B2(new_n733), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT58), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n721), .B1(new_n1169), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n719), .B1(new_n282), .B2(new_n820), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1178), .B(new_n1179), .C1(new_n1144), .C2(new_n780), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1157), .A2(new_n1159), .A3(new_n1180), .ZN(G375));
  NAND2_X1  g0981(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1077), .A2(new_n991), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n832), .A2(new_n779), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT120), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n718), .B1(G68), .B2(new_n821), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n750), .A2(new_n464), .B1(new_n724), .B2(new_n353), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n390), .B1(new_n747), .B2(new_n725), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1188), .A2(new_n1002), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n543), .B2(new_n732), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1187), .B(new_n1190), .C1(G116), .C2(new_n767), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1191), .B1(new_n512), .B2(new_n756), .C1(new_n452), .C2(new_n752), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n752), .A2(new_n1101), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n738), .A2(new_n282), .B1(new_n950), .B2(new_n756), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT121), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(G159), .B2(new_n751), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n733), .A2(G132), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n262), .B1(new_n724), .B2(new_n289), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT122), .Z(new_n1199));
  AOI22_X1  g0999(.A1(new_n748), .A2(G137), .B1(new_n767), .B2(new_n1112), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1196), .A2(new_n1197), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1192), .B1(new_n1193), .B2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1186), .B1(new_n1202), .B2(new_n721), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1185), .A2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n1073), .B2(new_n716), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1183), .A2(new_n1206), .ZN(G381));
  NOR2_X1   g1007(.A1(G375), .A2(G378), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  NOR3_X1   g1009(.A1(new_n1209), .A2(G384), .A3(G381), .ZN(new_n1210));
  OR2_X1    g1010(.A1(G390), .A2(G387), .ZN(new_n1211));
  NOR3_X1   g1011(.A1(new_n1211), .A2(G396), .A3(G393), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1210), .A2(new_n1212), .ZN(G407));
  OAI211_X1 g1013(.A(G407), .B(G213), .C1(G343), .C2(new_n1209), .ZN(G409));
  NAND2_X1  g1014(.A1(G390), .A2(G387), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1211), .A2(new_n1215), .ZN(new_n1216));
  XOR2_X1   g1016(.A(G393), .B(G396), .Z(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1217), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1211), .A2(new_n1215), .A3(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1157), .A2(G378), .A3(new_n1159), .A4(new_n1180), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n1097), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1151), .A2(new_n991), .A3(new_n1158), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1153), .A2(new_n717), .A3(new_n1155), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1224), .A2(new_n1225), .A3(new_n1180), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1223), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1222), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n638), .A2(G213), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(G384), .A2(KEYINPUT124), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT124), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n800), .A2(new_n1232), .A3(new_n822), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(KEYINPUT60), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n1182), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1073), .A2(KEYINPUT60), .A3(new_n1075), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1236), .A2(new_n657), .A3(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT123), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1236), .A2(KEYINPUT123), .A3(new_n657), .A4(new_n1237), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1234), .B1(new_n1242), .B2(new_n1206), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n1205), .B(new_n1233), .C1(new_n1240), .C2(new_n1241), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(KEYINPUT125), .B1(new_n1230), .B2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1221), .B1(new_n1246), .B2(KEYINPUT63), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n638), .A2(G213), .A3(G2897), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1233), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1242), .A2(new_n1206), .A3(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1248), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1205), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1251), .B(new_n1252), .C1(new_n1234), .C2(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1230), .A2(new_n1249), .A3(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT61), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT63), .ZN(new_n1258));
  OAI211_X1 g1058(.A(KEYINPUT125), .B(new_n1258), .C1(new_n1230), .C2(new_n1245), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1247), .A2(new_n1257), .A3(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(KEYINPUT62), .B1(new_n1230), .B2(new_n1245), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1251), .B1(new_n1234), .B2(new_n1253), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT62), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1262), .A2(new_n1263), .A3(new_n1229), .A4(new_n1228), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1261), .A2(new_n1255), .A3(new_n1256), .A4(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1221), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1260), .A2(new_n1266), .ZN(G405));
  INV_X1    g1067(.A(KEYINPUT127), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1218), .A2(new_n1268), .A3(new_n1220), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1221), .A2(KEYINPUT127), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(G375), .A2(new_n1223), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1245), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1222), .A2(KEYINPUT126), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1223), .B(G375), .C1(new_n1243), .C2(new_n1244), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1272), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1274), .B1(new_n1272), .B2(new_n1275), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1269), .B(new_n1270), .C1(new_n1276), .C2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1272), .A2(new_n1275), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1273), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1272), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1280), .A2(KEYINPUT127), .A3(new_n1221), .A4(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1278), .A2(new_n1282), .ZN(G402));
endmodule


