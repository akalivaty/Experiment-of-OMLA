//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 0 1 1 0 0 0 1 0 1 0 1 0 0 1 1 1 1 1 1 0 1 1 0 1 0 1 1 1 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0 0 0 1 1 1 0 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n573,
    new_n574, new_n575, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n632,
    new_n633, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1216, new_n1217;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT66), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n455), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OR3_X1    g033(.A1(new_n452), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n457), .B1(new_n452), .B2(new_n458), .ZN(new_n460));
  NAND3_X1  g035(.A1(new_n456), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n463), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n468), .A2(new_n472), .ZN(G160));
  OR2_X1    g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n463), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n463), .A2(G112), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n464), .A2(new_n465), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n480), .B1(G136), .B2(new_n482), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT68), .ZN(G162));
  INV_X1    g059(.A(G138), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n486), .B1(new_n464), .B2(new_n465), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT70), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n486), .B(new_n489), .C1(new_n465), .C2(new_n464), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n488), .A2(KEYINPUT4), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT69), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G114), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(KEYINPUT69), .ZN(new_n495));
  OAI21_X1  g070(.A(G2105), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n496), .A2(new_n498), .B1(new_n476), .B2(G126), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n487), .A2(KEYINPUT70), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n491), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  AND2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G50), .ZN(new_n509));
  XOR2_X1   g084(.A(new_n509), .B(KEYINPUT71), .Z(new_n510));
  NAND2_X1  g085(.A1(G75), .A2(G543), .ZN(new_n511));
  AND3_X1   g086(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n512));
  AOI21_X1  g087(.A(G543), .B1(KEYINPUT72), .B2(KEYINPUT5), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G62), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n511), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n512), .A2(new_n513), .B1(new_n504), .B2(new_n505), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n516), .A2(G651), .B1(new_n518), .B2(G88), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n510), .A2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  INV_X1    g096(.A(KEYINPUT73), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n522), .B1(new_n512), .B2(new_n513), .ZN(new_n523));
  NAND2_X1  g098(.A1(KEYINPUT72), .A2(KEYINPUT5), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(new_n507), .ZN(new_n525));
  NAND3_X1  g100(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n525), .A2(KEYINPUT73), .A3(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n523), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  XNOR2_X1  g104(.A(KEYINPUT6), .B(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n530), .A2(G51), .A3(G543), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT74), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT7), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n536), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(G89), .ZN(new_n539));
  OAI211_X1 g114(.A(new_n533), .B(new_n538), .C1(new_n517), .C2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n525), .A2(new_n526), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n542), .A2(G89), .A3(new_n530), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n533), .B1(new_n543), .B2(new_n538), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n532), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(KEYINPUT75), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT75), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n538), .B1(new_n517), .B2(new_n539), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(KEYINPUT74), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(new_n540), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n547), .B1(new_n550), .B2(new_n532), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n546), .A2(new_n551), .ZN(G286));
  INV_X1    g127(.A(G286), .ZN(G168));
  NAND2_X1  g128(.A1(G77), .A2(G543), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n523), .A2(new_n527), .ZN(new_n555));
  INV_X1    g130(.A(G64), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G651), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n518), .A2(G90), .B1(new_n508), .B2(G52), .ZN(new_n559));
  AND2_X1   g134(.A1(new_n558), .A2(new_n559), .ZN(G171));
  INV_X1    g135(.A(G651), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n523), .A2(new_n527), .A3(G56), .ZN(new_n562));
  NAND2_X1  g137(.A1(G68), .A2(G543), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n530), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G43), .ZN(new_n566));
  INV_X1    g141(.A(G81), .ZN(new_n567));
  OAI22_X1  g142(.A1(new_n565), .A2(new_n566), .B1(new_n517), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(new_n570));
  XOR2_X1   g145(.A(new_n570), .B(KEYINPUT76), .Z(G153));
  NAND4_X1  g146(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT77), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT8), .ZN(new_n575));
  NAND4_X1  g150(.A1(G319), .A2(G483), .A3(G661), .A4(new_n575), .ZN(G188));
  INV_X1    g151(.A(G53), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT9), .B1(new_n565), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT9), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n530), .A2(new_n579), .A3(G53), .A4(G543), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n578), .A2(new_n580), .B1(G91), .B2(new_n518), .ZN(new_n581));
  INV_X1    g156(.A(G65), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT78), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n583), .B1(new_n512), .B2(new_n513), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n525), .A2(KEYINPUT78), .A3(new_n526), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n582), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AND2_X1   g161(.A1(G78), .A2(G543), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n581), .A2(new_n588), .ZN(G299));
  NAND2_X1  g164(.A1(new_n558), .A2(new_n559), .ZN(G301));
  AOI22_X1  g165(.A1(new_n518), .A2(G87), .B1(new_n508), .B2(G49), .ZN(new_n591));
  AOI21_X1  g166(.A(G74), .B1(new_n523), .B2(new_n527), .ZN(new_n592));
  OAI21_X1  g167(.A(KEYINPUT79), .B1(new_n592), .B2(new_n561), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  NOR3_X1   g169(.A1(new_n592), .A2(KEYINPUT79), .A3(new_n561), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n591), .B1(new_n594), .B2(new_n595), .ZN(G288));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G61), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n514), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n599), .A2(G651), .B1(new_n518), .B2(G86), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT80), .ZN(new_n601));
  INV_X1    g176(.A(G48), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n565), .B2(new_n602), .ZN(new_n603));
  NAND4_X1  g178(.A1(new_n530), .A2(KEYINPUT80), .A3(G48), .A4(G543), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n600), .A2(new_n605), .ZN(G305));
  NAND3_X1  g181(.A1(new_n523), .A2(new_n527), .A3(G60), .ZN(new_n607));
  NAND2_X1  g182(.A1(G72), .A2(G543), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n561), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(G47), .ZN(new_n610));
  INV_X1    g185(.A(G85), .ZN(new_n611));
  OAI22_X1  g186(.A1(new_n565), .A2(new_n610), .B1(new_n517), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(G290));
  INV_X1    g189(.A(KEYINPUT10), .ZN(new_n615));
  INV_X1    g190(.A(G92), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n517), .B2(new_n616), .ZN(new_n617));
  NAND4_X1  g192(.A1(new_n542), .A2(KEYINPUT10), .A3(new_n530), .A4(G92), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n617), .A2(new_n618), .B1(G54), .B2(new_n508), .ZN(new_n619));
  INV_X1    g194(.A(G66), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n620), .B1(new_n584), .B2(new_n585), .ZN(new_n621));
  AND2_X1   g196(.A1(G79), .A2(G543), .ZN(new_n622));
  OAI21_X1  g197(.A(G651), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(G868), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G171), .B2(new_n625), .ZN(G284));
  OAI21_X1  g202(.A(new_n626), .B1(G171), .B2(new_n625), .ZN(G321));
  NOR2_X1   g203(.A1(G299), .A2(G868), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n629), .B1(G168), .B2(G868), .ZN(G297));
  XNOR2_X1  g205(.A(G297), .B(KEYINPUT81), .ZN(G280));
  INV_X1    g206(.A(new_n624), .ZN(new_n632));
  INV_X1    g207(.A(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n633), .B2(G860), .ZN(G148));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(G868), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(G868), .B2(new_n569), .ZN(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g213(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT12), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT13), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT82), .B(G2100), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT83), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n641), .A2(new_n642), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT84), .ZN(new_n646));
  AOI22_X1  g221(.A1(new_n482), .A2(G135), .B1(G123), .B2(new_n476), .ZN(new_n647));
  OAI21_X1  g222(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n648));
  INV_X1    g223(.A(G111), .ZN(new_n649));
  AOI22_X1  g224(.A1(new_n648), .A2(KEYINPUT85), .B1(new_n649), .B2(G2105), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(KEYINPUT85), .B2(new_n648), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(KEYINPUT86), .B(G2096), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n644), .A2(new_n646), .A3(new_n654), .ZN(G156));
  XNOR2_X1  g230(.A(G2427), .B(G2438), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2430), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT15), .B(G2435), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n659), .A2(KEYINPUT14), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2451), .B(G2454), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT16), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n661), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2443), .B(G2446), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1341), .B(G1348), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT87), .Z(new_n669));
  OAI21_X1  g244(.A(G14), .B1(new_n666), .B2(new_n667), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT88), .ZN(G401));
  XOR2_X1   g247(.A(KEYINPUT89), .B(KEYINPUT18), .Z(new_n673));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  XNOR2_X1  g249(.A(G2067), .B(G2678), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(KEYINPUT17), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n674), .A2(new_n675), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n673), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G2072), .B(G2078), .Z(new_n680));
  INV_X1    g255(.A(new_n673), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n680), .B1(new_n676), .B2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n679), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G2096), .B(G2100), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G227));
  XOR2_X1   g260(.A(G1971), .B(G1976), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1956), .B(G2474), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1961), .B(G1966), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  NOR3_X1   g266(.A1(new_n687), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n687), .A2(new_n690), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT20), .Z(new_n694));
  AOI211_X1 g269(.A(new_n692), .B(new_n694), .C1(new_n687), .C2(new_n691), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT90), .ZN(new_n696));
  XOR2_X1   g271(.A(G1981), .B(G1986), .Z(new_n697));
  XNOR2_X1  g272(.A(G1991), .B(G1996), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n696), .B(new_n701), .ZN(G229));
  INV_X1    g277(.A(G16), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n703), .A2(G22), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(G303), .B2(G16), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G1971), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT32), .B(G1981), .ZN(new_n707));
  MUX2_X1   g282(.A(G6), .B(G305), .S(G16), .Z(new_n708));
  AND2_X1   g283(.A1(new_n708), .A2(KEYINPUT91), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(KEYINPUT91), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n707), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n703), .A2(G23), .ZN(new_n713));
  INV_X1    g288(.A(new_n591), .ZN(new_n714));
  INV_X1    g289(.A(new_n592), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT79), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n715), .A2(new_n716), .A3(G651), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n714), .B1(new_n717), .B2(new_n593), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n713), .B1(new_n718), .B2(new_n703), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT92), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT33), .B(G1976), .Z(new_n721));
  OR2_X1    g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n720), .A2(new_n721), .ZN(new_n723));
  OR3_X1    g298(.A1(new_n709), .A2(new_n710), .A3(new_n707), .ZN(new_n724));
  NAND4_X1  g299(.A1(new_n712), .A2(new_n722), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n725), .A2(KEYINPUT34), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(KEYINPUT34), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n482), .A2(G131), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n476), .A2(G119), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n463), .A2(G107), .ZN(new_n730));
  OAI21_X1  g305(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n728), .B(new_n729), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  MUX2_X1   g307(.A(G25), .B(new_n732), .S(G29), .Z(new_n733));
  XOR2_X1   g308(.A(KEYINPUT35), .B(G1991), .Z(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n733), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n703), .A2(G24), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n613), .B2(new_n703), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n738), .A2(G1986), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n738), .A2(G1986), .ZN(new_n740));
  NOR3_X1   g315(.A1(new_n736), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n726), .A2(new_n727), .A3(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT93), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(KEYINPUT36), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT94), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n742), .A2(new_n745), .ZN(new_n747));
  INV_X1    g322(.A(G29), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G26), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT96), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT28), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n482), .A2(G140), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n476), .A2(G128), .ZN(new_n753));
  OR2_X1    g328(.A1(G104), .A2(G2105), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n754), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n752), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n751), .B1(new_n757), .B2(new_n748), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G2067), .ZN(new_n759));
  INV_X1    g334(.A(G2078), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n502), .A2(G29), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n748), .A2(G27), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n759), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT30), .B(G28), .ZN(new_n765));
  OR2_X1    g340(.A1(KEYINPUT31), .A2(G11), .ZN(new_n766));
  NAND2_X1  g341(.A1(KEYINPUT31), .A2(G11), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n765), .A2(new_n748), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n748), .A2(G32), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n482), .A2(G141), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n470), .A2(G105), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n476), .A2(G129), .ZN(new_n772));
  NAND3_X1  g347(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT26), .Z(new_n774));
  NAND4_X1  g349(.A1(new_n770), .A2(new_n771), .A3(new_n772), .A4(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n769), .B1(new_n776), .B2(new_n748), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT27), .B(G1996), .Z(new_n778));
  OAI221_X1 g353(.A(new_n768), .B1(new_n748), .B2(new_n652), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n763), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n779), .B1(G2078), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(G4), .A2(G16), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n632), .B2(G16), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n764), .B(new_n781), .C1(G1348), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n703), .A2(G5), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G171), .B2(new_n703), .ZN(new_n786));
  AOI22_X1  g361(.A1(G1961), .A2(new_n786), .B1(new_n783), .B2(G1348), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G1961), .B2(new_n786), .ZN(new_n788));
  NAND2_X1  g363(.A1(G115), .A2(G2104), .ZN(new_n789));
  INV_X1    g364(.A(G127), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n481), .B2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT97), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n463), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n792), .B2(new_n791), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT25), .ZN(new_n795));
  NAND2_X1  g370(.A1(G103), .A2(G2104), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n795), .B1(new_n796), .B2(G2105), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n463), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n482), .A2(G139), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n794), .A2(new_n799), .ZN(new_n800));
  MUX2_X1   g375(.A(G33), .B(new_n800), .S(G29), .Z(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(G2072), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(G2072), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT24), .ZN(new_n804));
  INV_X1    g379(.A(G34), .ZN(new_n805));
  AOI21_X1  g380(.A(G29), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n804), .B2(new_n805), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G160), .B2(new_n748), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n808), .A2(G2084), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n777), .A2(new_n778), .B1(G2084), .B2(new_n808), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n802), .A2(new_n803), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n784), .A2(new_n788), .A3(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(G29), .A2(G35), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G162), .B2(G29), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT29), .Z(new_n815));
  INV_X1    g390(.A(G2090), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT98), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n815), .A2(new_n816), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n703), .A2(G20), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT23), .Z(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(G299), .B2(G16), .ZN(new_n822));
  INV_X1    g397(.A(G1956), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n703), .A2(G19), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT95), .Z(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n569), .B2(new_n703), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G1341), .ZN(new_n828));
  NOR3_X1   g403(.A1(new_n819), .A2(new_n824), .A3(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(G16), .A2(G21), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(G168), .B2(G16), .ZN(new_n831));
  INV_X1    g406(.A(G1966), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  AND4_X1   g408(.A1(new_n812), .A2(new_n818), .A3(new_n829), .A4(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n746), .A2(new_n747), .A3(new_n834), .ZN(G150));
  INV_X1    g410(.A(G150), .ZN(G311));
  NAND2_X1  g411(.A1(new_n632), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT38), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n523), .A2(new_n527), .A3(G67), .ZN(new_n839));
  NAND2_X1  g414(.A1(G80), .A2(G543), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n561), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(G55), .ZN(new_n842));
  INV_X1    g417(.A(G93), .ZN(new_n843));
  OAI22_X1  g418(.A1(new_n565), .A2(new_n842), .B1(new_n517), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n569), .A2(new_n845), .ZN(new_n846));
  OAI22_X1  g421(.A1(new_n564), .A2(new_n568), .B1(new_n841), .B2(new_n844), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n838), .B(new_n849), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n850), .A2(KEYINPUT39), .ZN(new_n851));
  INV_X1    g426(.A(G860), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(KEYINPUT39), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n845), .A2(new_n852), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT37), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(G145));
  XNOR2_X1  g432(.A(new_n800), .B(new_n776), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n476), .A2(G130), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n463), .A2(G118), .ZN(new_n860));
  OAI21_X1  g435(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n862), .B1(G142), .B2(new_n482), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(new_n640), .Z(new_n864));
  XNOR2_X1  g439(.A(new_n858), .B(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n757), .B(new_n502), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n732), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n865), .B(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n652), .B(G160), .ZN(new_n869));
  XNOR2_X1  g444(.A(G162), .B(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(G37), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(new_n870), .B2(new_n868), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g448(.A(new_n848), .B(KEYINPUT99), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n635), .ZN(new_n875));
  NAND2_X1  g450(.A1(G299), .A2(new_n624), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n581), .A2(new_n619), .A3(new_n588), .A4(new_n623), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT41), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n876), .A2(new_n880), .A3(new_n877), .ZN(new_n881));
  XNOR2_X1  g456(.A(KEYINPUT100), .B(KEYINPUT41), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n882), .B1(new_n876), .B2(new_n877), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n879), .B1(new_n875), .B2(new_n885), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n886), .A2(KEYINPUT42), .ZN(new_n887));
  XOR2_X1   g462(.A(G303), .B(G305), .Z(new_n888));
  NAND2_X1  g463(.A1(G288), .A2(new_n613), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n718), .A2(G290), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(G303), .B(G305), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n893), .A2(new_n889), .A3(new_n890), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n886), .A2(KEYINPUT42), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n887), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n896), .B1(new_n887), .B2(new_n897), .ZN(new_n899));
  OAI21_X1  g474(.A(G868), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n625), .B1(new_n841), .B2(new_n844), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(G295));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n901), .ZN(G331));
  NAND2_X1  g478(.A1(new_n545), .A2(KEYINPUT75), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n550), .A2(new_n547), .A3(new_n532), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n904), .A2(G171), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(G171), .B1(new_n904), .B2(new_n905), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n849), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(KEYINPUT101), .ZN(new_n910));
  OAI21_X1  g485(.A(G301), .B1(new_n546), .B2(new_n551), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(new_n906), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT101), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(new_n913), .A3(new_n849), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n911), .A2(new_n848), .A3(new_n906), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n910), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n878), .A2(new_n880), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n878), .A2(new_n882), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n878), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n915), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n909), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n895), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n921), .A2(new_n910), .A3(new_n914), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n909), .A2(new_n915), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n885), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n924), .A2(new_n895), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(G37), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n930));
  NOR3_X1   g505(.A1(new_n923), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n884), .B1(new_n909), .B2(new_n915), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n913), .B1(new_n912), .B2(new_n849), .ZN(new_n933));
  AOI211_X1 g508(.A(KEYINPUT101), .B(new_n848), .C1(new_n911), .C2(new_n906), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n932), .B1(new_n935), .B2(new_n921), .ZN(new_n936));
  AOI21_X1  g511(.A(G37), .B1(new_n936), .B2(new_n895), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n895), .B1(new_n924), .B2(new_n926), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT43), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT44), .B1(new_n931), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n942));
  NOR3_X1   g517(.A1(new_n923), .A2(new_n929), .A3(KEYINPUT43), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n930), .B1(new_n937), .B2(new_n939), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT102), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n941), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n918), .A2(new_n917), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n948), .B1(new_n935), .B2(new_n915), .ZN(new_n949));
  INV_X1    g524(.A(new_n922), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n896), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n951), .A2(new_n937), .A3(KEYINPUT43), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n930), .B1(new_n929), .B2(new_n938), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n942), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n951), .A2(new_n937), .A3(new_n930), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT43), .B1(new_n929), .B2(new_n938), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT44), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT102), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n947), .A2(new_n958), .ZN(G397));
  AND3_X1   g534(.A1(new_n487), .A2(KEYINPUT70), .A3(new_n500), .ZN(new_n960));
  OAI211_X1 g535(.A(G126), .B(G2105), .C1(new_n464), .C2(new_n465), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n494), .A2(KEYINPUT69), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n492), .A2(G114), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n463), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n961), .B1(new_n964), .B2(new_n497), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n960), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(G1384), .B1(new_n966), .B2(new_n491), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT103), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT45), .ZN(new_n969));
  INV_X1    g544(.A(G1384), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n488), .A2(KEYINPUT4), .A3(new_n490), .ZN(new_n971));
  XNOR2_X1  g546(.A(KEYINPUT69), .B(G114), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n498), .B1(new_n972), .B2(new_n463), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n501), .A2(new_n973), .A3(new_n961), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n970), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT103), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n968), .A2(new_n969), .A3(new_n977), .ZN(new_n978));
  XOR2_X1   g553(.A(KEYINPUT104), .B(G40), .Z(new_n979));
  NOR3_X1   g554(.A1(new_n468), .A2(new_n472), .A3(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n756), .B(G2067), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n982), .A2(KEYINPUT106), .A3(new_n983), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n775), .B(G1996), .ZN(new_n988));
  AOI22_X1  g563(.A1(new_n986), .A2(new_n987), .B1(new_n982), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n982), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n732), .B(new_n734), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n982), .A2(G1986), .A3(G290), .ZN(new_n993));
  INV_X1    g568(.A(G1986), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n982), .A2(new_n994), .A3(new_n613), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n996), .B(KEYINPUT105), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n992), .A2(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n998), .B(KEYINPUT107), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT117), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT109), .ZN(new_n1001));
  XOR2_X1   g576(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n1002));
  AOI21_X1  g577(.A(new_n981), .B1(new_n967), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1004), .B1(new_n502), .B2(new_n970), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1003), .A2(new_n816), .A3(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n980), .B1(new_n967), .B2(KEYINPUT45), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n970), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n1001), .B(new_n1007), .C1(new_n1011), .C2(G1971), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n981), .B1(new_n975), .B2(new_n969), .ZN(new_n1013));
  AOI21_X1  g588(.A(G1971), .B1(new_n1013), .B2(new_n1009), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n970), .B(new_n1002), .C1(new_n971), .C2(new_n974), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n980), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n1016), .A2(G2090), .A3(new_n1005), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT109), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1012), .A2(new_n1018), .A3(G8), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT116), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(G303), .A2(G8), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1012), .A2(new_n1018), .A3(KEYINPUT116), .A4(G8), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n1021), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n502), .A2(new_n980), .A3(new_n970), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(G8), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(G305), .A2(G1981), .ZN(new_n1031));
  INV_X1    g606(.A(G1981), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n600), .A2(new_n605), .A3(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(KEYINPUT49), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT49), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT111), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AOI211_X1 g612(.A(KEYINPUT111), .B(KEYINPUT49), .C1(new_n1031), .C2(new_n1033), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1030), .B(new_n1034), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT110), .ZN(new_n1040));
  INV_X1    g615(.A(G1976), .ZN(new_n1041));
  NOR2_X1   g616(.A1(G288), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1040), .B1(new_n1042), .B2(new_n1029), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n718), .A2(G1976), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1030), .A2(KEYINPUT110), .A3(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1043), .A2(KEYINPUT52), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT52), .B1(G288), .B2(new_n1041), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1047), .A2(new_n1030), .A3(new_n1044), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1039), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1024), .A2(new_n1012), .A3(new_n1018), .A4(G8), .ZN(new_n1050));
  NAND2_X1  g625(.A1(G168), .A2(G8), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n980), .B(new_n1015), .C1(new_n967), .C2(new_n1004), .ZN(new_n1052));
  XOR2_X1   g627(.A(KEYINPUT114), .B(G2084), .Z(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT115), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT115), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1053), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1003), .A2(new_n1006), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT113), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT45), .B1(new_n502), .B2(new_n970), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1060), .B1(new_n1061), .B2(new_n981), .ZN(new_n1062));
  OAI211_X1 g637(.A(KEYINPUT113), .B(new_n980), .C1(new_n967), .C2(KEYINPUT45), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1062), .A2(new_n1063), .A3(new_n1009), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(new_n832), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1051), .B1(new_n1059), .B2(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1049), .A2(KEYINPUT63), .A3(new_n1050), .A4(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1000), .B1(new_n1027), .B2(new_n1067), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1066), .A2(KEYINPUT63), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1021), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1069), .A2(new_n1071), .A3(new_n1072), .A4(KEYINPUT117), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT63), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n502), .A2(new_n1004), .A3(new_n970), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1075), .B(new_n980), .C1(new_n967), .C2(new_n1002), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1076), .A2(G2090), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT112), .B1(new_n1077), .B2(new_n1014), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT112), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1002), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n981), .B1(new_n975), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1081), .A2(new_n816), .A3(new_n1075), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1079), .B(new_n1082), .C1(new_n1011), .C2(G1971), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1078), .A2(new_n1083), .A3(G8), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n1025), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1085), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1066), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1074), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1068), .A2(new_n1073), .A3(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1039), .A2(new_n1041), .A3(new_n718), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1029), .B1(new_n1090), .B2(new_n1033), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1050), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1091), .B1(new_n1092), .B2(new_n1049), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n1094));
  XNOR2_X1  g669(.A(G299), .B(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT56), .B(G2072), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1013), .A2(new_n1009), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(G1956), .B1(new_n1081), .B2(new_n1075), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1096), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1028), .A2(G2067), .ZN(new_n1102));
  INV_X1    g677(.A(G1348), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1102), .B1(new_n1052), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1101), .B1(new_n624), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1076), .A2(new_n823), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1106), .A2(new_n1095), .A3(new_n1098), .ZN(new_n1107));
  AND2_X1   g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1101), .A2(new_n1107), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT61), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT120), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1106), .A2(new_n1095), .A3(new_n1113), .A4(new_n1098), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1101), .A2(new_n1114), .A3(KEYINPUT61), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1107), .A2(KEYINPUT119), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1112), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n975), .A2(new_n969), .ZN(new_n1118));
  INV_X1    g693(.A(G1996), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1118), .A2(new_n1119), .A3(new_n980), .A4(new_n1009), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT58), .B(G1341), .Z(new_n1121));
  NAND2_X1  g696(.A1(new_n1028), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n569), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(KEYINPUT118), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT118), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1123), .A2(new_n1127), .A3(new_n569), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1125), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1127), .B1(new_n1123), .B2(new_n569), .ZN(new_n1130));
  INV_X1    g705(.A(new_n569), .ZN(new_n1131));
  AOI211_X1 g706(.A(KEYINPUT118), .B(new_n1131), .C1(new_n1120), .C2(new_n1122), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT59), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1129), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1106), .A2(new_n1098), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1110), .B1(new_n1135), .B2(new_n1096), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1107), .A2(KEYINPUT119), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1136), .A2(new_n1137), .A3(KEYINPUT120), .A4(new_n1114), .ZN(new_n1138));
  AND4_X1   g713(.A1(new_n1111), .A2(new_n1117), .A3(new_n1134), .A4(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1104), .A2(KEYINPUT60), .A3(new_n624), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n1140), .A2(KEYINPUT121), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1104), .A2(KEYINPUT60), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n632), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(KEYINPUT122), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1140), .A2(KEYINPUT121), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1142), .A2(new_n1146), .A3(new_n632), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1141), .A2(new_n1144), .A3(new_n1145), .A4(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1148), .B1(KEYINPUT60), .B2(new_n1104), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1108), .B1(new_n1139), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1010), .B1(new_n1008), .B2(new_n1060), .ZN(new_n1151));
  AOI21_X1  g726(.A(G1966), .B1(new_n1151), .B2(new_n1063), .ZN(new_n1152));
  OAI21_X1  g727(.A(G286), .B1(new_n1152), .B2(new_n1058), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1065), .A2(G168), .A3(new_n1054), .A4(new_n1057), .ZN(new_n1154));
  AND4_X1   g729(.A1(KEYINPUT51), .A2(new_n1153), .A3(G8), .A4(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(KEYINPUT51), .B1(new_n1154), .B2(G8), .ZN(new_n1156));
  OAI21_X1  g731(.A(KEYINPUT123), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  XOR2_X1   g732(.A(KEYINPUT124), .B(KEYINPUT54), .Z(new_n1158));
  NAND3_X1  g733(.A1(new_n1013), .A2(new_n760), .A3(new_n1009), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT53), .ZN(new_n1160));
  INV_X1    g735(.A(G1961), .ZN(new_n1161));
  AOI22_X1  g736(.A1(new_n1159), .A2(new_n1160), .B1(new_n1161), .B2(new_n1052), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT125), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n472), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(KEYINPUT125), .B1(new_n469), .B2(new_n471), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1160), .A2(G2078), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(G40), .ZN(new_n1167));
  NOR4_X1   g742(.A1(new_n1164), .A2(new_n1165), .A3(new_n468), .A4(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n978), .A2(new_n1009), .A3(new_n1168), .ZN(new_n1169));
  AND3_X1   g744(.A1(new_n1162), .A2(G301), .A3(new_n1169), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1062), .A2(new_n1063), .A3(new_n1009), .A4(new_n1166), .ZN(new_n1171));
  AOI21_X1  g746(.A(G301), .B1(new_n1162), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1158), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1052), .A2(new_n1161), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1174), .A2(new_n1169), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(G171), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1162), .A2(G301), .A3(new_n1171), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1177), .A2(KEYINPUT54), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1173), .A2(new_n1179), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1180), .A2(new_n1086), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1154), .A2(G8), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT51), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT123), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1153), .A2(new_n1154), .A3(KEYINPUT51), .A4(G8), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1157), .A2(new_n1181), .A3(new_n1187), .ZN(new_n1188));
  OAI211_X1 g763(.A(new_n1089), .B(new_n1093), .C1(new_n1150), .C2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT62), .ZN(new_n1190));
  AND3_X1   g765(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1185), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1190), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1157), .A2(KEYINPUT62), .A3(new_n1187), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1172), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1086), .A2(new_n1195), .ZN(new_n1196));
  AND3_X1   g771(.A1(new_n1193), .A2(new_n1194), .A3(new_n1196), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n999), .B1(new_n1189), .B2(new_n1197), .ZN(new_n1198));
  XOR2_X1   g773(.A(new_n995), .B(KEYINPUT127), .Z(new_n1199));
  XNOR2_X1  g774(.A(new_n1199), .B(KEYINPUT48), .ZN(new_n1200));
  NOR2_X1   g775(.A1(new_n756), .A2(G2067), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n732), .A2(new_n735), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1201), .B1(new_n989), .B2(new_n1202), .ZN(new_n1203));
  OAI22_X1  g778(.A1(new_n1200), .A2(new_n992), .B1(new_n1203), .B2(new_n990), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n982), .A2(new_n1119), .ZN(new_n1205));
  XNOR2_X1  g780(.A(new_n1205), .B(KEYINPUT46), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n982), .B1(new_n775), .B2(new_n983), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  XOR2_X1   g783(.A(new_n1208), .B(KEYINPUT126), .Z(new_n1209));
  INV_X1    g784(.A(KEYINPUT47), .ZN(new_n1210));
  OR2_X1    g785(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n1204), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1198), .A2(new_n1213), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g789(.A1(new_n671), .A2(G229), .A3(new_n461), .A4(G227), .ZN(new_n1216));
  NAND2_X1  g790(.A1(new_n955), .A2(new_n956), .ZN(new_n1217));
  NAND3_X1  g791(.A1(new_n1216), .A2(new_n872), .A3(new_n1217), .ZN(G225));
  INV_X1    g792(.A(G225), .ZN(G308));
endmodule


