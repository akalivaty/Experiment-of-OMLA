//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 1 1 1 1 1 1 0 1 1 0 0 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 0 0 0 0 0 0 0 0 1 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0002(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n203));
  INV_X1    g0003(.A(G87), .ZN(new_n204));
  INV_X1    g0004(.A(G250), .ZN(new_n205));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G257), .ZN(new_n207));
  OAI221_X1 g0007(.A(new_n203), .B1(new_n204), .B2(new_n205), .C1(new_n206), .C2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(KEYINPUT64), .ZN(new_n209));
  AOI21_X1  g0009(.A(new_n209), .B1(G50), .B2(G226), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G68), .A2(G238), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n208), .A2(KEYINPUT64), .ZN(new_n212));
  AND3_X1   g0012(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G77), .ZN(new_n214));
  INV_X1    g0014(.A(G244), .ZN(new_n215));
  INV_X1    g0015(.A(G116), .ZN(new_n216));
  INV_X1    g0016(.A(G270), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G20), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT1), .Z(new_n221));
  NOR2_X1   g0021(.A1(new_n219), .A2(G13), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT0), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(G58), .A2(G68), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n221), .B(new_n224), .C1(new_n228), .C2(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT65), .Z(G361));
  XNOR2_X1  g0033(.A(KEYINPUT66), .B(G264), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n217), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n237), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  INV_X1    g0049(.A(KEYINPUT69), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n250), .B1(new_n219), .B2(new_n251), .ZN(new_n252));
  NAND4_X1  g0052(.A1(KEYINPUT69), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n252), .A2(new_n225), .A3(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G1), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n254), .B1(new_n255), .B2(G20), .ZN(new_n256));
  OAI21_X1  g0056(.A(G20), .B1(new_n230), .B2(G50), .ZN(new_n257));
  INV_X1    g0057(.A(G150), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n226), .A2(G33), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT8), .B(G58), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n257), .B1(new_n258), .B2(new_n260), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  AOI22_X1  g0063(.A1(G50), .A2(new_n256), .B1(new_n263), .B2(new_n254), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n255), .A2(G13), .A3(G20), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n264), .B1(G50), .B2(new_n265), .ZN(new_n266));
  XNOR2_X1  g0066(.A(new_n266), .B(KEYINPUT9), .ZN(new_n267));
  INV_X1    g0067(.A(G190), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT3), .B(G33), .ZN(new_n269));
  INV_X1    g0069(.A(G1698), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G222), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G223), .A2(G1698), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G41), .ZN(new_n274));
  OAI211_X1 g0074(.A(G1), .B(G13), .C1(new_n251), .C2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n273), .B(new_n276), .C1(G77), .C2(new_n269), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n255), .B1(G41), .B2(G45), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G226), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT67), .B(G45), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n255), .B(G274), .C1(new_n282), .C2(G41), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n277), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  OR2_X1    g0084(.A1(new_n284), .A2(KEYINPUT68), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(KEYINPUT68), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n268), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT70), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n285), .A2(new_n286), .ZN(new_n289));
  INV_X1    g0089(.A(G200), .ZN(new_n290));
  OAI22_X1  g0090(.A1(new_n287), .A2(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n285), .A2(KEYINPUT70), .A3(G200), .A4(new_n286), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n267), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT10), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT10), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n267), .A2(new_n291), .A3(new_n295), .A4(new_n292), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G179), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n289), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G169), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n285), .A2(new_n300), .A3(new_n286), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n299), .A2(new_n266), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n297), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(G238), .A2(G1698), .ZN(new_n304));
  INV_X1    g0104(.A(G232), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n269), .B(new_n304), .C1(new_n305), .C2(G1698), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n306), .B(new_n276), .C1(G107), .C2(new_n269), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n280), .A2(G244), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n307), .A2(new_n283), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n300), .ZN(new_n310));
  OAI22_X1  g0110(.A1(new_n262), .A2(new_n260), .B1(new_n226), .B2(new_n214), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT15), .B(G87), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n312), .A2(new_n261), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n254), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n265), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n214), .ZN(new_n316));
  INV_X1    g0116(.A(new_n256), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n314), .B(new_n316), .C1(new_n317), .C2(new_n214), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n307), .A2(new_n298), .A3(new_n283), .A4(new_n308), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n310), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n303), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n226), .A2(G33), .A3(G77), .ZN(new_n323));
  INV_X1    g0123(.A(G68), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G20), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT72), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n323), .A2(KEYINPUT72), .A3(new_n325), .ZN(new_n329));
  INV_X1    g0129(.A(G50), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n328), .B(new_n329), .C1(new_n330), .C2(new_n260), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n254), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT11), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G13), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n335), .A2(G1), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(G20), .A3(new_n324), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT12), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT73), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n256), .A2(G68), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n331), .A2(KEYINPUT11), .A3(new_n254), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n334), .A2(new_n341), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n338), .A2(KEYINPUT73), .ZN(new_n345));
  NOR3_X1   g0145(.A1(new_n337), .A2(new_n345), .A3(new_n340), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n279), .A2(KEYINPUT71), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT71), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n275), .A2(new_n349), .A3(new_n278), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n348), .A2(G238), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(G33), .A2(G97), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n305), .A2(G1698), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(G226), .B2(G1698), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT3), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(G33), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n352), .B1(new_n354), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n276), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n351), .A2(new_n360), .A3(new_n283), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT13), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT13), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n351), .A2(new_n363), .A3(new_n360), .A4(new_n283), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(G200), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n362), .A2(G190), .A3(new_n364), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n347), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT14), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n370), .B1(new_n365), .B2(G169), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n365), .A2(new_n298), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n365), .A2(new_n370), .A3(G169), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n372), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n347), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n369), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT74), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(new_n356), .B2(G33), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n251), .A2(KEYINPUT74), .A3(KEYINPUT3), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n355), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT7), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n382), .A2(new_n383), .A3(new_n226), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n356), .A2(G33), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT74), .B1(new_n251), .B2(KEYINPUT3), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n379), .A2(new_n356), .A3(G33), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(KEYINPUT7), .B1(new_n388), .B2(G20), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n384), .A2(new_n389), .A3(G68), .ZN(new_n390));
  INV_X1    g0190(.A(G58), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n391), .A2(new_n324), .ZN(new_n392));
  OAI21_X1  g0192(.A(G20), .B1(new_n392), .B2(new_n229), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n259), .A2(G159), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n390), .A2(KEYINPUT16), .A3(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT16), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n383), .B1(new_n269), .B2(G20), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n358), .A2(KEYINPUT7), .A3(new_n226), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n324), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n398), .B1(new_n401), .B2(new_n395), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n397), .A2(new_n254), .A3(new_n402), .ZN(new_n403));
  MUX2_X1   g0203(.A(new_n317), .B(new_n265), .S(new_n262), .Z(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n386), .A2(new_n387), .ZN(new_n406));
  OR2_X1    g0206(.A1(G223), .A2(G1698), .ZN(new_n407));
  OR2_X1    g0207(.A1(new_n270), .A2(G226), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n406), .A2(new_n355), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G33), .A2(G87), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n276), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n275), .A2(G232), .A3(new_n278), .ZN(new_n413));
  AOI21_X1  g0213(.A(KEYINPUT75), .B1(new_n283), .B2(new_n413), .ZN(new_n414));
  AND3_X1   g0214(.A1(new_n283), .A2(KEYINPUT75), .A3(new_n413), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n412), .B(G179), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT76), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n275), .B1(new_n409), .B2(new_n410), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n283), .A2(new_n413), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT75), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n283), .A2(KEYINPUT75), .A3(new_n413), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n418), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n416), .B(new_n417), .C1(new_n300), .C2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n415), .A2(new_n414), .ZN(new_n426));
  OAI21_X1  g0226(.A(G169), .B1(new_n426), .B2(new_n418), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n417), .B1(new_n427), .B2(new_n416), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n405), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT18), .ZN(new_n430));
  INV_X1    g0230(.A(new_n416), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n421), .A2(new_n422), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n300), .B1(new_n432), .B2(new_n412), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT76), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n424), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT18), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(new_n436), .A3(new_n405), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n430), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT78), .ZN(new_n439));
  OAI21_X1  g0239(.A(G200), .B1(new_n426), .B2(new_n418), .ZN(new_n440));
  OR2_X1    g0240(.A1(new_n268), .A2(KEYINPUT77), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n268), .A2(KEYINPUT77), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n432), .A2(new_n412), .A3(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n403), .A2(new_n440), .A3(new_n445), .A4(new_n404), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT17), .ZN(new_n447));
  AND2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n446), .A2(new_n447), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n439), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n403), .A2(new_n445), .A3(new_n404), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n451), .A2(KEYINPUT17), .A3(new_n440), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n446), .A2(new_n447), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n452), .A2(KEYINPUT78), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n438), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n309), .A2(G200), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n309), .A2(new_n268), .ZN(new_n457));
  OR3_X1    g0257(.A1(new_n456), .A2(new_n457), .A3(new_n318), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n322), .A2(new_n378), .A3(new_n455), .A4(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT83), .ZN(new_n460));
  INV_X1    g0260(.A(new_n312), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(new_n265), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n406), .A2(new_n226), .A3(G68), .A4(new_n355), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT19), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n464), .A2(new_n226), .A3(G33), .A4(G97), .ZN(new_n465));
  NOR2_X1   g0265(.A1(G97), .A2(G107), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n466), .A2(new_n204), .B1(new_n352), .B2(new_n226), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n465), .B1(new_n467), .B2(new_n464), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n462), .B1(new_n469), .B2(new_n254), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n265), .B1(G1), .B2(new_n251), .ZN(new_n471));
  NOR3_X1   g0271(.A1(new_n254), .A2(new_n312), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n460), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n254), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n475), .B1(new_n463), .B2(new_n468), .ZN(new_n476));
  NOR4_X1   g0276(.A1(new_n476), .A2(new_n472), .A3(KEYINPUT83), .A4(new_n462), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n255), .A2(G45), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT82), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(new_n480), .A3(G250), .ZN(new_n481));
  AOI21_X1  g0281(.A(G274), .B1(KEYINPUT82), .B2(G250), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n481), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n275), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n251), .A2(new_n216), .ZN(new_n485));
  NOR2_X1   g0285(.A1(G238), .A2(G1698), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n486), .B1(new_n215), .B2(G1698), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n485), .B1(new_n388), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n484), .B1(new_n488), .B2(new_n275), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G169), .ZN(new_n490));
  OAI211_X1 g0290(.A(G179), .B(new_n484), .C1(new_n488), .C2(new_n275), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g0292(.A(G190), .B(new_n484), .C1(new_n488), .C2(new_n275), .ZN(new_n493));
  XNOR2_X1  g0293(.A(new_n493), .B(KEYINPUT84), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n489), .A2(G200), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n254), .A2(new_n471), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G87), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n495), .A2(new_n470), .A3(new_n497), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n478), .A2(new_n492), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT81), .ZN(new_n500));
  INV_X1    g0300(.A(G283), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n251), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n355), .A2(new_n357), .A3(G250), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT4), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n502), .B1(new_n504), .B2(G1698), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n406), .A2(G244), .A3(new_n355), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT4), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n358), .A2(new_n215), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n507), .A2(G1698), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n505), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(G45), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n513), .A2(G1), .ZN(new_n514));
  AND2_X1   g0314(.A1(KEYINPUT5), .A2(G41), .ZN(new_n515));
  NOR2_X1   g0315(.A1(KEYINPUT5), .A2(G41), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n517), .A2(G257), .A3(new_n275), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n514), .B(G274), .C1(new_n516), .C2(new_n515), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT80), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n518), .A2(KEYINPUT80), .A3(new_n519), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n512), .A2(new_n276), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n500), .B1(new_n524), .B2(new_n290), .ZN(new_n525));
  XNOR2_X1  g0325(.A(G97), .B(G107), .ZN(new_n526));
  NOR2_X1   g0326(.A1(KEYINPUT79), .A2(KEYINPUT6), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(KEYINPUT6), .A2(G107), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(KEYINPUT79), .B2(KEYINPUT6), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n528), .B1(new_n526), .B2(new_n530), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n531), .A2(G20), .B1(G77), .B2(new_n259), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n399), .A2(new_n400), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(G107), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n475), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  OR2_X1    g0335(.A1(new_n254), .A2(new_n471), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n536), .A2(new_n206), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n265), .A2(G97), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n535), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n524), .A2(G190), .ZN(new_n540));
  INV_X1    g0340(.A(new_n523), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT80), .B1(new_n518), .B2(new_n519), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n506), .A2(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n275), .B1(new_n544), .B2(new_n505), .ZN(new_n545));
  OAI211_X1 g0345(.A(KEYINPUT81), .B(G200), .C1(new_n543), .C2(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n525), .A2(new_n539), .A3(new_n540), .A4(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n496), .A2(G107), .ZN(new_n548));
  INV_X1    g0348(.A(new_n336), .ZN(new_n549));
  INV_X1    g0349(.A(G107), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G20), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g0352(.A(new_n552), .B(KEYINPUT25), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT22), .ZN(new_n554));
  NOR3_X1   g0354(.A1(new_n554), .A2(new_n204), .A3(G20), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n406), .A2(new_n355), .A3(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n355), .A2(new_n357), .A3(new_n226), .A4(G87), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n554), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT23), .ZN(new_n559));
  XNOR2_X1  g0359(.A(new_n551), .B(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n485), .A2(new_n226), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n556), .A2(new_n558), .A3(new_n560), .A4(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT90), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n563), .A2(KEYINPUT24), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n388), .A2(new_n555), .B1(new_n557), .B2(new_n554), .ZN(new_n566));
  INV_X1    g0366(.A(new_n564), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n566), .A2(new_n567), .A3(new_n560), .A4(new_n561), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n565), .A2(new_n568), .B1(new_n563), .B2(KEYINPUT24), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n548), .B(new_n553), .C1(new_n569), .C2(new_n475), .ZN(new_n570));
  AND3_X1   g0370(.A1(new_n517), .A2(G264), .A3(new_n275), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n205), .A2(new_n270), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n207), .A2(G1698), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n388), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(G33), .A2(G294), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n571), .B1(new_n576), .B2(new_n276), .ZN(new_n577));
  AOI21_X1  g0377(.A(G169), .B1(new_n577), .B2(new_n519), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n275), .B1(new_n574), .B2(new_n575), .ZN(new_n579));
  INV_X1    g0379(.A(new_n519), .ZN(new_n580));
  NOR4_X1   g0380(.A1(new_n579), .A2(G179), .A3(new_n580), .A4(new_n571), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n570), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n537), .ZN(new_n584));
  INV_X1    g0384(.A(new_n538), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n531), .A2(G20), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n259), .A2(G77), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n534), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n584), .B(new_n585), .C1(new_n588), .C2(new_n475), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n524), .A2(new_n298), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n300), .B1(new_n543), .B2(new_n545), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n499), .A2(new_n547), .A3(new_n583), .A4(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n570), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n577), .A2(new_n519), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(G200), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n577), .A2(G190), .A3(new_n519), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n594), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(KEYINPUT86), .A2(KEYINPUT20), .ZN(new_n600));
  AOI21_X1  g0400(.A(G20), .B1(G33), .B2(G283), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n251), .A2(G97), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n601), .A2(new_n602), .B1(G20), .B2(new_n216), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n254), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(KEYINPUT86), .A2(KEYINPUT20), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n254), .A2(new_n605), .A3(new_n603), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n600), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n315), .A2(G116), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n610), .B1(new_n536), .B2(G116), .ZN(new_n611));
  OAI21_X1  g0411(.A(G169), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n517), .A2(new_n275), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n519), .B1(new_n613), .B2(new_n217), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n207), .A2(G1698), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n355), .B(new_n615), .C1(new_n380), .C2(new_n381), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT85), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n388), .A2(KEYINPUT85), .A3(new_n615), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n388), .A2(G264), .A3(G1698), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n358), .A2(G303), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n618), .A2(new_n619), .A3(new_n620), .A4(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n614), .B1(new_n622), .B2(new_n276), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n612), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(KEYINPUT21), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT87), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n254), .A2(new_n605), .A3(new_n603), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n605), .B1(new_n254), .B2(new_n603), .ZN(new_n628));
  OAI22_X1  g0428(.A1(new_n627), .A2(new_n628), .B1(KEYINPUT86), .B2(KEYINPUT20), .ZN(new_n629));
  INV_X1    g0429(.A(new_n610), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n496), .B2(new_n216), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n298), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n626), .B1(new_n632), .B2(new_n623), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n632), .A2(new_n626), .A3(new_n623), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n625), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT88), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n636), .B1(new_n612), .B2(new_n623), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n622), .A2(new_n276), .ZN(new_n638));
  INV_X1    g0438(.A(new_n614), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n300), .B1(new_n629), .B2(new_n631), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(new_n641), .A3(KEYINPUT88), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT21), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n637), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT89), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n637), .A2(new_n642), .A3(KEYINPUT89), .A4(new_n643), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n635), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n623), .A2(new_n444), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n609), .A2(new_n611), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n649), .B(new_n650), .C1(new_n290), .C2(new_n623), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n599), .A2(new_n648), .A3(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n459), .A2(new_n652), .ZN(G372));
  INV_X1    g0453(.A(new_n302), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n427), .A2(new_n416), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n405), .A2(new_n655), .A3(KEYINPUT18), .ZN(new_n656));
  AOI21_X1  g0456(.A(KEYINPUT18), .B1(new_n405), .B2(new_n655), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n376), .A2(new_n377), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n369), .B2(new_n320), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n450), .A2(new_n454), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n654), .B1(new_n663), .B2(new_n297), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n470), .A2(new_n473), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n498), .A2(new_n493), .B1(new_n492), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n594), .A2(new_n596), .A3(new_n597), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n668), .A2(new_n592), .A3(new_n547), .ZN(new_n669));
  AOI211_X1 g0469(.A(new_n667), .B(new_n669), .C1(new_n648), .C2(new_n583), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n494), .A2(new_n498), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n665), .A2(KEYINPUT83), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n470), .A2(new_n460), .A3(new_n473), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(new_n492), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(KEYINPUT26), .B1(new_n675), .B2(new_n592), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n492), .A2(new_n665), .ZN(new_n677));
  XOR2_X1   g0477(.A(new_n677), .B(KEYINPUT91), .Z(new_n678));
  AND3_X1   g0478(.A1(new_n589), .A2(new_n591), .A3(new_n590), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT26), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(new_n680), .A3(new_n666), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n676), .A2(new_n678), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT92), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n676), .A2(new_n678), .A3(new_n681), .A4(KEYINPUT92), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n670), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n664), .B1(new_n459), .B2(new_n687), .ZN(G369));
  OR3_X1    g0488(.A1(new_n549), .A2(KEYINPUT27), .A3(G20), .ZN(new_n689));
  OAI21_X1  g0489(.A(KEYINPUT27), .B1(new_n549), .B2(G20), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G213), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(G343), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n650), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n648), .A2(new_n651), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n648), .B2(new_n696), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G330), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n583), .A2(new_n693), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n668), .B1(new_n594), .B2(new_n694), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n700), .B1(new_n701), .B2(new_n583), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n648), .A2(new_n693), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n700), .B1(new_n706), .B2(new_n702), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n705), .A2(new_n707), .ZN(G399));
  INV_X1    g0508(.A(new_n222), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G41), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n466), .A2(new_n204), .A3(new_n216), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n711), .A2(G1), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n231), .B2(new_n711), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT28), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n648), .A2(new_n583), .ZN(new_n717));
  INV_X1    g0517(.A(new_n669), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(new_n718), .A3(new_n666), .ZN(new_n719));
  OAI21_X1  g0519(.A(KEYINPUT26), .B1(new_n667), .B2(new_n592), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n499), .A2(new_n679), .A3(new_n680), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n720), .A2(new_n721), .A3(new_n678), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n693), .B1(new_n719), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT29), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n491), .A2(new_n579), .A3(new_n571), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n726), .A2(new_n524), .A3(new_n623), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT30), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n726), .A2(new_n524), .A3(KEYINPUT30), .A4(new_n623), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n640), .A2(KEYINPUT93), .A3(new_n298), .A4(new_n489), .ZN(new_n732));
  INV_X1    g0532(.A(new_n524), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n732), .A2(new_n595), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n640), .A2(new_n298), .A3(new_n489), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT93), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n731), .B1(new_n734), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(KEYINPUT31), .B1(new_n738), .B2(new_n694), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n737), .A2(new_n595), .A3(new_n733), .A4(new_n732), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(new_n729), .A3(new_n730), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT31), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n741), .A2(new_n742), .A3(new_n693), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n599), .A2(new_n648), .A3(new_n651), .A4(new_n694), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G330), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n724), .B(new_n694), .C1(new_n670), .C2(new_n686), .ZN(new_n748));
  AND3_X1   g0548(.A1(new_n725), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n716), .B1(new_n749), .B2(G1), .ZN(G364));
  AOI21_X1  g0550(.A(new_n225), .B1(G20), .B2(new_n300), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G179), .A2(G200), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n752), .A2(G20), .A3(new_n268), .ZN(new_n753));
  OR2_X1    g0553(.A1(new_n753), .A2(KEYINPUT95), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(KEYINPUT95), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AND2_X1   g0557(.A1(new_n757), .A2(KEYINPUT96), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(KEYINPUT96), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n226), .A2(new_n298), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G200), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n443), .A2(new_n763), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n761), .A2(G329), .B1(G326), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n762), .A2(new_n290), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G190), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n269), .B1(new_n767), .B2(G311), .ZN(new_n768));
  INV_X1    g0568(.A(G303), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n226), .A2(G179), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(G190), .A3(G200), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n763), .A2(G190), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  XOR2_X1   g0573(.A(KEYINPUT33), .B(G317), .Z(new_n774));
  OAI221_X1 g0574(.A(new_n768), .B1(new_n769), .B2(new_n771), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n443), .A2(new_n766), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n775), .B1(G322), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n770), .A2(new_n268), .A3(G200), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n765), .B(new_n777), .C1(new_n501), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n752), .A2(G190), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n779), .B1(G294), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G159), .ZN(new_n783));
  OR3_X1    g0583(.A1(new_n756), .A2(KEYINPUT32), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n781), .A2(G97), .ZN(new_n785));
  OAI21_X1  g0585(.A(KEYINPUT32), .B1(new_n756), .B2(new_n783), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n771), .A2(new_n204), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n784), .A2(new_n785), .A3(new_n786), .A4(new_n788), .ZN(new_n789));
  AOI22_X1  g0589(.A1(G68), .A2(new_n772), .B1(new_n767), .B2(G77), .ZN(new_n790));
  INV_X1    g0590(.A(new_n764), .ZN(new_n791));
  INV_X1    g0591(.A(new_n776), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n790), .B1(new_n330), .B2(new_n791), .C1(new_n391), .C2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n778), .A2(new_n550), .ZN(new_n794));
  NOR4_X1   g0594(.A1(new_n789), .A2(new_n793), .A3(new_n358), .A4(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n751), .B1(new_n782), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n335), .A2(G20), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(G45), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n711), .A2(G1), .A3(new_n798), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT94), .Z(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n388), .A2(new_n709), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n802), .B1(new_n231), .B2(new_n282), .C1(new_n245), .C2(new_n513), .ZN(new_n803));
  INV_X1    g0603(.A(G355), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n269), .A2(new_n222), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n803), .B1(G116), .B2(new_n222), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(G13), .A2(G33), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(G20), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n751), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n801), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n809), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n796), .B(new_n811), .C1(new_n698), .C2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n699), .A2(new_n801), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n698), .A2(G330), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(G396));
  XNOR2_X1  g0616(.A(new_n320), .B(KEYINPUT99), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n318), .A2(new_n693), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n817), .A2(new_n458), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(KEYINPUT100), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT100), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n817), .A2(new_n821), .A3(new_n458), .A4(new_n818), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n820), .A2(new_n822), .B1(new_n321), .B2(new_n693), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n687), .B2(new_n693), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n820), .A2(new_n822), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n694), .B(new_n826), .C1(new_n670), .C2(new_n686), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(new_n747), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n829), .A2(new_n801), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n761), .A2(G311), .B1(G116), .B2(new_n767), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n785), .B1(new_n791), .B2(new_n769), .ZN(new_n832));
  XNOR2_X1  g0632(.A(KEYINPUT97), .B(G283), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n773), .A2(new_n834), .B1(new_n204), .B2(new_n778), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(G294), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n831), .B(new_n836), .C1(new_n837), .C2(new_n792), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n358), .B1(new_n771), .B2(new_n550), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(KEYINPUT98), .Z(new_n840));
  AOI21_X1  g0640(.A(new_n382), .B1(new_n761), .B2(G132), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n778), .A2(new_n324), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(G58), .B2(new_n781), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n841), .B(new_n843), .C1(new_n330), .C2(new_n771), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n776), .A2(G143), .B1(new_n767), .B2(G159), .ZN(new_n845));
  INV_X1    g0645(.A(G137), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n845), .B1(new_n846), .B2(new_n791), .C1(new_n258), .C2(new_n773), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT34), .Z(new_n848));
  OAI22_X1  g0648(.A1(new_n838), .A2(new_n840), .B1(new_n844), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n801), .B1(new_n849), .B2(new_n751), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n751), .A2(new_n807), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n823), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n850), .B1(G77), .B2(new_n852), .C1(new_n853), .C2(new_n808), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT101), .Z(new_n855));
  NOR2_X1   g0655(.A1(new_n830), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(G384));
  INV_X1    g0657(.A(KEYINPUT37), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n397), .A2(new_n254), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT16), .B1(new_n390), .B2(new_n396), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n404), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n691), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n451), .A2(new_n440), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n861), .A2(new_n655), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n858), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n405), .A2(new_n862), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT102), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n405), .A2(KEYINPUT102), .A3(new_n862), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n871), .A2(new_n858), .A3(new_n446), .A4(new_n429), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n866), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n861), .A2(new_n862), .ZN(new_n874));
  OAI211_X1 g0674(.A(KEYINPUT38), .B(new_n873), .C1(new_n455), .C2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n405), .A2(new_n655), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT102), .B1(new_n405), .B2(new_n862), .ZN(new_n877));
  AOI211_X1 g0677(.A(new_n868), .B(new_n691), .C1(new_n403), .C2(new_n404), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n446), .B(new_n876), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT37), .ZN(new_n880));
  INV_X1    g0680(.A(new_n871), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n452), .B(new_n453), .C1(new_n656), .C2(new_n657), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n872), .A2(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT103), .B1(new_n883), .B2(KEYINPUT38), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT38), .ZN(new_n885));
  AOI221_X4 g0685(.A(KEYINPUT18), .B1(new_n403), .B2(new_n404), .C1(new_n434), .C2(new_n424), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n436), .B1(new_n435), .B2(new_n405), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n874), .B1(new_n661), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n446), .B1(new_n877), .B2(new_n878), .ZN(new_n890));
  INV_X1    g0690(.A(new_n429), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n865), .B1(new_n892), .B2(new_n858), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n885), .B1(new_n889), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n875), .A2(new_n884), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT39), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n872), .A2(new_n880), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n881), .A2(new_n882), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n885), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT103), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT39), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n875), .A2(new_n899), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n896), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n659), .A2(new_n693), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n817), .A2(new_n693), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n827), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n875), .A2(new_n894), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n377), .B(new_n693), .C1(new_n376), .C2(new_n369), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n377), .A2(new_n693), .ZN(new_n911));
  AOI211_X1 g0711(.A(KEYINPUT14), .B(new_n300), .C1(new_n362), .C2(new_n364), .ZN(new_n912));
  NOR3_X1   g0712(.A1(new_n371), .A2(new_n912), .A3(new_n373), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n368), .B(new_n911), .C1(new_n913), .C2(new_n347), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n908), .A2(new_n909), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n658), .A2(new_n691), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n905), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n725), .A2(new_n748), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n664), .B1(new_n920), .B2(new_n459), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n919), .B(new_n921), .ZN(new_n922));
  AND3_X1   g0722(.A1(new_n746), .A2(new_n853), .A3(new_n916), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n909), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT40), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(new_n875), .B2(new_n899), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n924), .A2(new_n925), .B1(new_n923), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n459), .B1(new_n745), .B2(new_n744), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n927), .B(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(G330), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n922), .B(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n255), .B2(new_n797), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n216), .B1(new_n531), .B2(KEYINPUT35), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n934), .B(new_n227), .C1(KEYINPUT35), .C2(new_n531), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT36), .ZN(new_n936));
  OAI21_X1  g0736(.A(G77), .B1(new_n391), .B2(new_n324), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n231), .A2(new_n937), .B1(G50), .B2(new_n324), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n938), .A2(G1), .A3(new_n335), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n933), .A2(new_n936), .A3(new_n939), .ZN(G367));
  AND2_X1   g0740(.A1(new_n237), .A2(new_n802), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n810), .B1(new_n222), .B2(new_n312), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n800), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n771), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT46), .B1(new_n944), .B2(G116), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n388), .B1(new_n767), .B2(new_n833), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n944), .A2(KEYINPUT46), .A3(G116), .ZN(new_n947));
  INV_X1    g0747(.A(G317), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n946), .B(new_n947), .C1(new_n948), .C2(new_n756), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n945), .B(new_n949), .C1(G107), .C2(new_n781), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n778), .A2(new_n206), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(new_n764), .B2(G311), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n953), .B1(new_n837), .B2(new_n773), .C1(new_n769), .C2(new_n792), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n269), .B1(new_n778), .B2(new_n214), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n764), .A2(G143), .B1(new_n772), .B2(G159), .ZN(new_n956));
  INV_X1    g0756(.A(new_n767), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n956), .B1(new_n330), .B2(new_n957), .C1(new_n391), .C2(new_n771), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n955), .B(new_n958), .C1(G68), .C2(new_n781), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n959), .B1(new_n846), .B2(new_n756), .C1(new_n258), .C2(new_n792), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n954), .A2(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n962));
  XNOR2_X1  g0762(.A(new_n961), .B(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n943), .B1(new_n963), .B2(new_n751), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT109), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n470), .A2(new_n497), .ZN(new_n966));
  OR3_X1    g0766(.A1(new_n678), .A2(new_n966), .A3(new_n694), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n666), .B1(new_n966), .B2(new_n694), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n965), .B1(new_n809), .B2(new_n970), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n547), .B(new_n592), .C1(new_n539), .C2(new_n694), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n679), .A2(new_n693), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n704), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT105), .ZN(new_n976));
  XNOR2_X1  g0776(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n970), .A2(new_n977), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n976), .A2(new_n978), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n706), .A2(new_n702), .A3(new_n974), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT42), .Z(new_n983));
  OAI21_X1  g0783(.A(new_n592), .B1(new_n972), .B2(new_n583), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n694), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n981), .B(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n710), .B(KEYINPUT41), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n707), .A2(new_n974), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT45), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(KEYINPUT45), .B1(new_n707), .B2(new_n974), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OR3_X1    g0795(.A1(new_n707), .A2(KEYINPUT44), .A3(new_n974), .ZN(new_n996));
  OAI21_X1  g0796(.A(KEYINPUT44), .B1(new_n707), .B2(new_n974), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n705), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n704), .B1(new_n995), .B2(new_n998), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n706), .ZN(new_n1003));
  AOI21_X1  g0803(.A(KEYINPUT106), .B1(new_n1003), .B2(new_n703), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n706), .A2(new_n702), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n698), .A2(G330), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1006), .B1(new_n698), .B2(G330), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1005), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1009), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1011), .A2(new_n1004), .A3(new_n1007), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  AND3_X1   g0813(.A1(new_n749), .A2(new_n1013), .A3(KEYINPUT107), .ZN(new_n1014));
  AOI21_X1  g0814(.A(KEYINPUT107), .B1(new_n749), .B2(new_n1013), .ZN(new_n1015));
  NOR3_X1   g0815(.A1(new_n1002), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n749), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n990), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n798), .A2(G1), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n971), .B1(new_n989), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(G387));
  OAI221_X1 g0823(.A(new_n710), .B1(new_n749), .B2(new_n1013), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1013), .A2(new_n1019), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT110), .Z(new_n1026));
  INV_X1    g0826(.A(new_n282), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n802), .B1(new_n241), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n713), .B2(new_n805), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n324), .A2(new_n214), .ZN(new_n1030));
  OR3_X1    g0830(.A1(new_n262), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1031));
  OAI21_X1  g0831(.A(KEYINPUT50), .B1(new_n262), .B2(G50), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1031), .A2(new_n513), .A3(new_n713), .A4(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1029), .B1(new_n1030), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n709), .A2(new_n550), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n751), .B(new_n809), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n791), .A2(new_n783), .B1(new_n773), .B2(new_n262), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(G150), .B2(new_n757), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n330), .B2(new_n792), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n944), .A2(G77), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n781), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1040), .B1(new_n312), .B2(new_n1041), .ZN(new_n1042));
  NOR3_X1   g0842(.A1(new_n1039), .A2(new_n951), .A3(new_n1042), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1043), .B(new_n388), .C1(new_n324), .C2(new_n957), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n776), .A2(G317), .B1(new_n772), .B2(G311), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(KEYINPUT111), .B(G322), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1045), .B1(new_n769), .B2(new_n957), .C1(new_n791), .C2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT48), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n837), .B2(new_n771), .C1(new_n1041), .C2(new_n834), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT49), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n757), .A2(G326), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n778), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(G116), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1052), .A2(new_n382), .A3(new_n1053), .A4(new_n1055), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1044), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n801), .B(new_n1036), .C1(new_n1058), .C2(new_n751), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n702), .B2(new_n812), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1024), .A2(new_n1026), .A3(new_n1060), .ZN(G393));
  NOR2_X1   g0861(.A1(new_n957), .A2(new_n262), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G150), .A2(new_n764), .B1(new_n776), .B2(G159), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT51), .Z(new_n1064));
  AOI22_X1  g0864(.A1(new_n944), .A2(G68), .B1(new_n1054), .B2(G87), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n772), .A2(G50), .B1(G77), .B2(new_n781), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1064), .A2(new_n388), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n1062), .B(new_n1067), .C1(G143), .C2(new_n757), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G311), .A2(new_n776), .B1(new_n764), .B2(G317), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT52), .Z(new_n1070));
  OAI221_X1 g0870(.A(new_n1070), .B1(new_n216), .B2(new_n1041), .C1(new_n771), .C2(new_n834), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n756), .A2(new_n1047), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n794), .B1(G303), .B2(new_n772), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n837), .B2(new_n957), .ZN(new_n1074));
  NOR4_X1   g0874(.A1(new_n1071), .A2(new_n269), .A3(new_n1072), .A4(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n751), .B1(new_n1068), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n810), .B1(new_n206), .B2(new_n222), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(new_n248), .B2(new_n802), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT112), .Z(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n800), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT113), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1076), .B(new_n1081), .C1(new_n812), .C2(new_n974), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT115), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1002), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT114), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n710), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1002), .B(KEYINPUT114), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1084), .B1(new_n1088), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n711), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1095), .A2(KEYINPUT115), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1083), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1090), .A2(new_n1019), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(G390));
  OAI21_X1  g0899(.A(new_n915), .B1(new_n747), .B2(new_n823), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n930), .B1(new_n744), .B2(new_n745), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1101), .A2(new_n853), .A3(new_n916), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n908), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT116), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n746), .B2(G330), .ZN(new_n1106));
  AOI211_X1 g0906(.A(KEYINPUT116), .B(new_n930), .C1(new_n744), .C2(new_n745), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n916), .B1(new_n1108), .B2(new_n853), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n906), .B1(new_n723), .B2(new_n826), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n1102), .ZN(new_n1111));
  NOR3_X1   g0911(.A1(new_n1109), .A2(KEYINPUT117), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT117), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n747), .A2(KEYINPUT116), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1114), .A2(new_n853), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n915), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1111), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1113), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1104), .B1(new_n1112), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n928), .A2(G330), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1121), .B(new_n664), .C1(new_n459), .C2(new_n920), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n904), .B1(new_n875), .B2(new_n899), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n1110), .B2(new_n915), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n904), .B1(new_n908), .B2(new_n916), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1126), .B1(new_n903), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1102), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1126), .B(new_n1102), .C1(new_n903), .C2(new_n1127), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n711), .B1(new_n1124), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n1132), .B2(new_n1124), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n851), .A2(new_n262), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n800), .A2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n903), .A2(new_n808), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n216), .A2(new_n792), .B1(new_n791), .B2(new_n501), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n761), .B2(G294), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(G97), .A2(new_n767), .B1(new_n772), .B2(G107), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1140), .B(KEYINPUT118), .Z(new_n1141));
  AOI211_X1 g0941(.A(new_n269), .B(new_n842), .C1(G77), .C2(new_n781), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1139), .A2(new_n788), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT119), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n761), .A2(G125), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n764), .A2(G128), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n772), .A2(G137), .ZN(new_n1147));
  OR3_X1    g0947(.A1(new_n771), .A2(KEYINPUT53), .A3(new_n258), .ZN(new_n1148));
  OAI21_X1  g0948(.A(KEYINPUT53), .B1(new_n771), .B2(new_n258), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n358), .B1(new_n781), .B2(G159), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  XOR2_X1   g0951(.A(KEYINPUT54), .B(G143), .Z(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n957), .A2(new_n1153), .B1(new_n330), .B2(new_n778), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1151), .B(new_n1154), .C1(G132), .C2(new_n776), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .A4(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1144), .A2(new_n1156), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1136), .B(new_n1137), .C1(new_n751), .C2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1132), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1158), .B1(new_n1159), .B2(new_n1019), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1134), .A2(new_n1160), .ZN(G378));
  INV_X1    g0961(.A(new_n1104), .ZN(new_n1162));
  OAI21_X1  g0962(.A(KEYINPUT117), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1117), .A2(new_n1113), .A3(new_n1118), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1162), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1123), .B1(new_n1132), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n926), .A2(new_n923), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n746), .A2(new_n853), .A3(new_n916), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(new_n894), .B2(new_n875), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1167), .B(G330), .C1(new_n1169), .C2(KEYINPUT40), .ZN(new_n1170));
  XOR2_X1   g0970(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1171));
  NAND2_X1  g0971(.A1(new_n303), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1171), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n297), .A2(new_n302), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n266), .A2(new_n862), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1172), .A2(new_n266), .A3(new_n862), .A4(new_n1174), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(KEYINPUT121), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1170), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1180), .B1(new_n927), .B2(G330), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n919), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1170), .A2(new_n1181), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n927), .A2(G330), .A3(new_n1180), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n903), .A2(new_n904), .B1(new_n658), .B2(new_n691), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .A4(new_n917), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1184), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1166), .A2(KEYINPUT57), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n710), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT122), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  AND2_X1   g0993(.A1(new_n1166), .A2(new_n1189), .ZN(new_n1194));
  OAI21_X1  g0994(.A(KEYINPUT123), .B1(new_n1194), .B2(KEYINPUT57), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1190), .A2(KEYINPUT122), .A3(new_n710), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1166), .A2(new_n1189), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT123), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT57), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1193), .A2(new_n1195), .A3(new_n1196), .A4(new_n1200), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n274), .B(new_n382), .C1(new_n792), .C2(new_n550), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n778), .A2(new_n391), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n461), .B2(new_n767), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1204), .B(new_n1040), .C1(new_n324), .C2(new_n1041), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1202), .B(new_n1205), .C1(G97), .C2(new_n772), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n216), .B2(new_n791), .C1(new_n501), .C2(new_n760), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT58), .ZN(new_n1208));
  INV_X1    g1008(.A(G124), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n274), .B1(new_n756), .B2(new_n1209), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n764), .A2(G125), .B1(new_n772), .B2(G132), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n776), .A2(G128), .B1(G150), .B2(new_n781), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(new_n846), .C2(new_n957), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n944), .B2(new_n1152), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT59), .ZN(new_n1215));
  AOI211_X1 g1015(.A(G33), .B(new_n1210), .C1(new_n1214), .C2(new_n1215), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1216), .B1(new_n1215), .B2(new_n1214), .C1(new_n783), .C2(new_n778), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n251), .B1(new_n386), .B2(new_n387), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n330), .B1(new_n1218), .B2(G41), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1208), .A2(new_n1217), .A3(new_n1219), .ZN(new_n1220));
  XOR2_X1   g1020(.A(new_n1220), .B(KEYINPUT120), .Z(new_n1221));
  AOI21_X1  g1021(.A(new_n801), .B1(new_n1221), .B2(new_n751), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(G50), .B2(new_n852), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n808), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n1189), .B2(new_n1019), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1201), .A2(new_n1226), .ZN(G375));
  OAI211_X1 g1027(.A(new_n1122), .B(new_n1104), .C1(new_n1112), .C2(new_n1119), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1124), .A2(new_n990), .A3(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n915), .A2(new_n807), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n852), .A2(G68), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n767), .A2(G150), .B1(G50), .B2(new_n781), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(KEYINPUT124), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1203), .B(new_n1233), .C1(G137), .C2(new_n776), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n772), .A2(new_n1152), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n761), .A2(G128), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n382), .B1(new_n764), .B2(G132), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n771), .A2(new_n783), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n957), .A2(new_n550), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n761), .A2(G303), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n773), .A2(new_n216), .B1(new_n214), .B2(new_n778), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n269), .B(new_n1242), .C1(G294), .C2(new_n764), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n776), .A2(G283), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n944), .A2(G97), .B1(new_n461), .B2(new_n781), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1241), .A2(new_n1243), .A3(new_n1244), .A4(new_n1245), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n1238), .A2(new_n1239), .B1(new_n1240), .B2(new_n1246), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n801), .B(new_n1231), .C1(new_n1247), .C2(new_n751), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n1120), .A2(new_n1019), .B1(new_n1230), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1229), .A2(new_n1249), .ZN(G381));
  INV_X1    g1050(.A(new_n1226), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n1190), .A2(KEYINPUT122), .A3(new_n710), .ZN(new_n1252));
  AOI21_X1  g1052(.A(KEYINPUT122), .B1(new_n1190), .B2(new_n710), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1198), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1255));
  AOI211_X1 g1055(.A(KEYINPUT123), .B(KEYINPUT57), .C1(new_n1166), .C2(new_n1189), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1251), .B1(new_n1254), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(G378), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1097), .A2(new_n1022), .A3(new_n1098), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(G393), .A2(G396), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  OR4_X1    g1063(.A1(G384), .A2(new_n1260), .A3(new_n1263), .A4(G381), .ZN(G407));
  OAI211_X1 g1064(.A(G407), .B(G213), .C1(G343), .C2(new_n1260), .ZN(G409));
  INV_X1    g1065(.A(KEYINPUT62), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1266), .A2(KEYINPUT127), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n692), .A2(G213), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1251), .B1(new_n990), .B2(new_n1194), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1259), .A2(new_n1269), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1268), .B(new_n1270), .C1(new_n1258), .C2(new_n1259), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT125), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT60), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1228), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1165), .A2(KEYINPUT60), .A3(new_n1122), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1274), .A2(new_n1275), .A3(new_n1124), .A4(new_n710), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(G384), .A3(new_n1249), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(G384), .B1(new_n1276), .B2(new_n1249), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1272), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1279), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1281), .A2(KEYINPUT125), .A3(new_n1277), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1280), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1267), .B1(new_n1271), .B2(new_n1284), .ZN(new_n1285));
  XOR2_X1   g1085(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1286));
  NAND3_X1  g1086(.A1(new_n692), .A2(G213), .A3(G2897), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(new_n1281), .B2(new_n1277), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1288), .B1(new_n1283), .B2(new_n1287), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1286), .B1(new_n1271), .B2(new_n1289), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(G375), .A2(G378), .B1(G213), .B2(new_n692), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1291), .A2(new_n1270), .A3(new_n1283), .A4(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1285), .A2(new_n1290), .A3(new_n1293), .ZN(new_n1294));
  XOR2_X1   g1094(.A(G393), .B(G396), .Z(new_n1295));
  AOI21_X1  g1095(.A(new_n1022), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1295), .B1(new_n1261), .B2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(G390), .A2(G387), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1097), .A2(new_n1022), .A3(new_n1098), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1295), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1298), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1297), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1294), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(G375), .A2(G378), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1304), .A2(new_n1268), .A3(new_n1270), .A4(new_n1283), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT63), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1302), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT61), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1271), .A2(new_n1289), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1291), .A2(KEYINPUT63), .A3(new_n1270), .A4(new_n1283), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1307), .A2(new_n1308), .A3(new_n1309), .A4(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1303), .A2(new_n1311), .ZN(G405));
  NAND2_X1  g1112(.A1(new_n1260), .A2(new_n1304), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1281), .A2(new_n1277), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1260), .A2(new_n1304), .A3(new_n1283), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(new_n1317), .B(new_n1302), .ZN(G402));
endmodule


