//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 1 0 1 1 0 0 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 0 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 0 1 0 1 1 0 1 1 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967;
  NAND2_X1  g000(.A1(G234), .A2(G237), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  AND3_X1   g002(.A1(new_n187), .A2(G952), .A3(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT21), .B(G898), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(KEYINPUT95), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n187), .A2(G902), .A3(G953), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n192), .B(KEYINPUT94), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n189), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  OAI21_X1  g008(.A(G210), .B1(G237), .B2(G902), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G143), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(KEYINPUT0), .A2(G128), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  NOR3_X1   g019(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n206));
  INV_X1    g020(.A(new_n202), .ZN(new_n207));
  NOR3_X1   g021(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n203), .B1(new_n201), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G125), .ZN(new_n210));
  OR2_X1    g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G128), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(KEYINPUT1), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(new_n198), .A3(new_n200), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n199), .B(G146), .C1(new_n212), .C2(KEYINPUT1), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n212), .A2(new_n197), .A3(G143), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n215), .A2(KEYINPUT66), .A3(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(KEYINPUT66), .B1(new_n215), .B2(new_n216), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n214), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(new_n210), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n211), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n188), .A2(G224), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n222), .B(new_n223), .ZN(new_n224));
  XOR2_X1   g038(.A(G110), .B(G122), .Z(new_n225));
  INV_X1    g039(.A(G104), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT3), .B1(new_n226), .B2(G107), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT76), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n226), .A2(G107), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n231));
  INV_X1    g045(.A(G107), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n232), .A3(G104), .ZN(new_n233));
  OAI211_X1 g047(.A(KEYINPUT76), .B(KEYINPUT3), .C1(new_n226), .C2(G107), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n229), .A2(new_n230), .A3(new_n233), .A4(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G101), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n233), .A2(new_n230), .ZN(new_n237));
  INV_X1    g051(.A(G101), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n237), .A2(new_n238), .A3(new_n229), .A4(new_n234), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n236), .A2(KEYINPUT4), .A3(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(G116), .B(G119), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT2), .B(G113), .ZN(new_n243));
  NOR3_X1   g057(.A1(new_n242), .A2(KEYINPUT67), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT67), .ZN(new_n245));
  XOR2_X1   g059(.A(KEYINPUT2), .B(G113), .Z(new_n246));
  AOI21_X1  g060(.A(new_n245), .B1(new_n246), .B2(new_n241), .ZN(new_n247));
  OAI22_X1  g061(.A1(new_n244), .A2(new_n247), .B1(new_n241), .B2(new_n246), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n235), .A2(new_n249), .A3(G101), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n240), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT82), .ZN(new_n252));
  INV_X1    g066(.A(new_n230), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n226), .A2(G107), .ZN(new_n254));
  OAI21_X1  g068(.A(G101), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n239), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT67), .B1(new_n242), .B2(new_n243), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n246), .A2(new_n245), .A3(new_n241), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n260));
  INV_X1    g074(.A(G119), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n261), .A3(G116), .ZN(new_n262));
  OAI211_X1 g076(.A(G113), .B(new_n262), .C1(new_n242), .C2(new_n260), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n256), .A2(new_n259), .A3(new_n263), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n251), .A2(new_n252), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n252), .B1(new_n251), .B2(new_n264), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n225), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n225), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n251), .A2(new_n264), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT6), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  OAI211_X1 g085(.A(KEYINPUT6), .B(new_n225), .C1(new_n265), .C2(new_n266), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n224), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G902), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT84), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n239), .A2(new_n255), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT83), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(new_n259), .A3(new_n263), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n256), .A2(KEYINPUT84), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n259), .A2(new_n263), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n281), .B(new_n275), .C1(new_n277), .C2(new_n276), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n279), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  XOR2_X1   g097(.A(new_n225), .B(KEYINPUT8), .Z(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT85), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n220), .A2(new_n286), .A3(new_n210), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n223), .A2(KEYINPUT7), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n287), .B(new_n288), .C1(new_n222), .C2(new_n286), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  OR2_X1    g104(.A1(new_n222), .A2(new_n288), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n269), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n274), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n196), .B1(new_n273), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n251), .A2(new_n264), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT82), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n251), .A2(new_n264), .A3(new_n252), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n268), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n270), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n272), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n224), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n287), .A2(new_n288), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n211), .A2(new_n221), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n303), .B1(new_n304), .B2(KEYINPUT85), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n305), .B1(new_n284), .B2(new_n283), .ZN(new_n306));
  INV_X1    g120(.A(new_n292), .ZN(new_n307));
  AOI21_X1  g121(.A(G902), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n302), .A2(new_n195), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n294), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(G214), .B1(G237), .B2(G902), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n311), .B(KEYINPUT81), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT86), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT86), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n310), .A2(new_n315), .A3(new_n312), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n194), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT11), .ZN(new_n318));
  INV_X1    g132(.A(G134), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n318), .B1(new_n319), .B2(G137), .ZN(new_n320));
  INV_X1    g134(.A(G137), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(KEYINPUT11), .A3(G134), .ZN(new_n322));
  INV_X1    g136(.A(G131), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n319), .A2(G137), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n320), .A2(new_n322), .A3(new_n323), .A4(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n321), .A2(G134), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n319), .A2(G137), .ZN(new_n327));
  OAI21_X1  g141(.A(G131), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT65), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT65), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n325), .A2(new_n328), .A3(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n330), .A2(new_n219), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT30), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n320), .A2(new_n324), .A3(new_n322), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G131), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n325), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n209), .A2(new_n337), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n333), .A2(new_n334), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n329), .A2(KEYINPUT68), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT68), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n325), .A2(new_n328), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(new_n219), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n334), .B1(new_n343), .B2(new_n338), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n248), .B1(new_n339), .B2(new_n344), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n257), .A2(new_n258), .B1(new_n242), .B2(new_n243), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n343), .A2(new_n346), .A3(new_n338), .ZN(new_n347));
  XOR2_X1   g161(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n348));
  NOR2_X1   g162(.A1(G237), .A2(G953), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G210), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n348), .B(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(KEYINPUT26), .B(G101), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n351), .B(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n345), .A2(new_n347), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT31), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n347), .A2(KEYINPUT28), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT28), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n343), .A2(new_n338), .A3(new_n346), .A4(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n333), .A2(new_n338), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n248), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n353), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT31), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n345), .A2(new_n365), .A3(new_n347), .A4(new_n353), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n355), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G472), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n368), .A3(new_n274), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT32), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n367), .A2(KEYINPUT32), .A3(new_n368), .A4(new_n274), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n343), .A2(new_n338), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n373), .A2(new_n346), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n374), .B1(new_n356), .B2(new_n358), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT29), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n363), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(G902), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n376), .B1(new_n362), .B2(new_n363), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n353), .B1(new_n345), .B2(new_n347), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G472), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n371), .A2(new_n372), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(KEYINPUT22), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n385), .B(new_n321), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n212), .A2(G119), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n261), .A2(G128), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(KEYINPUT24), .B(G110), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT73), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n389), .A2(new_n390), .A3(KEYINPUT73), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT23), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n387), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n212), .A2(KEYINPUT23), .A3(G119), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n388), .A3(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(KEYINPUT72), .B(G110), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n393), .B(new_n394), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(G140), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n210), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(G125), .A2(G140), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT16), .ZN(new_n405));
  NOR3_X1   g219(.A1(new_n210), .A2(KEYINPUT16), .A3(G140), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n405), .A2(G146), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n404), .A2(new_n197), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n400), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT16), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n411), .B1(new_n402), .B2(new_n403), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n197), .B1(new_n412), .B2(new_n406), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n398), .A2(G110), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT71), .ZN(new_n416));
  OR2_X1    g230(.A1(new_n389), .A2(new_n390), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT71), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n398), .A2(new_n418), .A3(G110), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n414), .A2(new_n416), .A3(new_n417), .A4(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n410), .A2(new_n420), .A3(KEYINPUT74), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(KEYINPUT74), .B1(new_n410), .B2(new_n420), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n386), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n386), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(new_n410), .A3(new_n420), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n424), .A2(new_n274), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT25), .ZN(new_n428));
  XOR2_X1   g242(.A(KEYINPUT70), .B(G217), .Z(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n430), .B1(G234), .B2(new_n274), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT25), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n424), .A2(new_n426), .A3(new_n432), .A4(new_n274), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n428), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n431), .A2(G902), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n424), .A2(new_n426), .A3(new_n435), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n383), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G221), .ZN(new_n439));
  XOR2_X1   g253(.A(KEYINPUT9), .B(G234), .Z(new_n440));
  AOI21_X1  g254(.A(new_n439), .B1(new_n440), .B2(new_n274), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n239), .A2(new_n255), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT77), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n239), .A2(KEYINPUT77), .A3(new_n255), .A4(new_n443), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  XOR2_X1   g262(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n256), .A2(KEYINPUT10), .A3(new_n219), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n240), .A2(new_n209), .A3(new_n250), .ZN(new_n453));
  XOR2_X1   g267(.A(new_n337), .B(KEYINPUT79), .Z(new_n454));
  NAND4_X1  g268(.A1(new_n451), .A2(new_n452), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n449), .B1(new_n446), .B2(new_n447), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n240), .A2(new_n209), .A3(new_n250), .ZN(new_n457));
  INV_X1    g271(.A(new_n452), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n337), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n455), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(G110), .B(G140), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(KEYINPUT75), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n188), .A2(G227), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n463), .B(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n220), .A2(new_n276), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n448), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT80), .ZN(new_n469));
  AOI21_X1  g283(.A(KEYINPUT12), .B1(new_n337), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n468), .A2(new_n337), .A3(new_n471), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n446), .A2(new_n447), .B1(new_n220), .B2(new_n276), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n470), .B1(new_n473), .B2(new_n460), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n465), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(new_n455), .A3(new_n476), .ZN(new_n477));
  AOI211_X1 g291(.A(G469), .B(G902), .C1(new_n466), .C2(new_n477), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n455), .B(new_n476), .C1(new_n459), .C2(new_n460), .ZN(new_n479));
  AOI22_X1  g293(.A1(new_n459), .A2(new_n454), .B1(new_n472), .B2(new_n474), .ZN(new_n480));
  OAI211_X1 g294(.A(G469), .B(new_n479), .C1(new_n480), .C2(new_n476), .ZN(new_n481));
  NAND2_X1  g295(.A1(G469), .A2(G902), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n442), .B1(new_n478), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(G475), .A2(G902), .ZN(new_n485));
  XNOR2_X1  g299(.A(G113), .B(G122), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(new_n226), .ZN(new_n487));
  INV_X1    g301(.A(new_n404), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(G146), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(KEYINPUT87), .A3(new_n409), .ZN(new_n490));
  INV_X1    g304(.A(G237), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(new_n188), .A3(G214), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n199), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n349), .A2(G143), .A3(G214), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n323), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(KEYINPUT18), .ZN(new_n496));
  NAND2_X1  g310(.A1(KEYINPUT18), .A2(G131), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n493), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  OR3_X1    g312(.A1(new_n404), .A2(KEYINPUT87), .A3(new_n197), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n490), .A2(new_n496), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n495), .A2(KEYINPUT17), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n408), .A2(new_n413), .A3(KEYINPUT89), .ZN(new_n502));
  AOI21_X1  g316(.A(KEYINPUT89), .B1(new_n408), .B2(new_n413), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n494), .ZN(new_n505));
  AOI21_X1  g319(.A(G143), .B1(new_n349), .B2(G214), .ZN(new_n506));
  OAI21_X1  g320(.A(G131), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT17), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n493), .A2(new_n323), .A3(new_n494), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT90), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT90), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n507), .A2(new_n512), .A3(new_n508), .A4(new_n509), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n487), .B(new_n500), .C1(new_n504), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n507), .A2(new_n509), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n408), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT88), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT19), .ZN(new_n519));
  OR2_X1    g333(.A1(new_n518), .A2(KEYINPUT19), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n488), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n404), .A2(new_n518), .A3(KEYINPUT19), .ZN(new_n522));
  AOI21_X1  g336(.A(G146), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n500), .B1(new_n517), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n487), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n515), .A2(KEYINPUT91), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(KEYINPUT91), .B1(new_n515), .B2(new_n526), .ZN(new_n528));
  OAI211_X1 g342(.A(KEYINPUT20), .B(new_n485), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT89), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n414), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n408), .A2(new_n413), .A3(KEYINPUT89), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n533), .A2(new_n501), .A3(new_n511), .A4(new_n513), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n487), .B1(new_n534), .B2(new_n500), .ZN(new_n535));
  INV_X1    g349(.A(new_n515), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n274), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(G475), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n515), .A2(new_n526), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n485), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT20), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n529), .A2(new_n538), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(G116), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(G122), .ZN(new_n546));
  INV_X1    g360(.A(G122), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(G116), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT92), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(G116), .B(G122), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(KEYINPUT92), .ZN(new_n553));
  OAI21_X1  g367(.A(G107), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n549), .A2(new_n550), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n552), .A2(KEYINPUT92), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(new_n556), .A3(new_n232), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n212), .A2(G143), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n199), .A2(G128), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n560), .A3(new_n319), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT13), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n562), .A2(new_n199), .A3(G128), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n559), .A2(new_n560), .ZN(new_n564));
  OAI211_X1 g378(.A(G134), .B(new_n563), .C1(new_n564), .C2(new_n562), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT93), .ZN(new_n566));
  OR2_X1    g380(.A1(new_n565), .A2(KEYINPUT93), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n558), .A2(new_n561), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n429), .A2(new_n440), .A3(new_n188), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n564), .A2(G134), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n561), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n545), .A2(KEYINPUT14), .A3(G122), .ZN(new_n573));
  OAI211_X1 g387(.A(G107), .B(new_n573), .C1(new_n549), .C2(KEYINPUT14), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n557), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n568), .A2(new_n570), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n570), .B1(new_n568), .B2(new_n575), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n274), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(G478), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(KEYINPUT15), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n568), .A2(new_n575), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n569), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n576), .ZN(new_n585));
  INV_X1    g399(.A(new_n581), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n274), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n582), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n544), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n484), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n317), .A2(new_n438), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(G101), .ZN(G3));
  NAND2_X1  g407(.A1(new_n367), .A2(new_n274), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(G472), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n369), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n475), .A2(new_n455), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n465), .B1(new_n459), .B2(new_n454), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n337), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n598), .A2(new_n465), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(G469), .B1(new_n602), .B2(G902), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n466), .A2(new_n477), .ZN(new_n604));
  INV_X1    g418(.A(G469), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(new_n605), .A3(new_n274), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n441), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n597), .A2(new_n437), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT96), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT96), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n597), .A2(new_n607), .A3(new_n610), .A4(new_n437), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n311), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n613), .B1(new_n294), .B2(new_n309), .ZN(new_n614));
  INV_X1    g428(.A(new_n194), .ZN(new_n615));
  NAND2_X1  g429(.A1(KEYINPUT97), .A2(KEYINPUT33), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n585), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n616), .ZN(new_n618));
  NOR2_X1   g432(.A1(KEYINPUT97), .A2(KEYINPUT33), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n584), .B(new_n576), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n617), .A2(G478), .A3(new_n620), .A4(new_n274), .ZN(new_n621));
  INV_X1    g435(.A(new_n579), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT98), .B(G478), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n614), .A2(new_n543), .A3(new_n615), .A4(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n612), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT34), .B(G104), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G6));
  OAI21_X1  g442(.A(new_n485), .B1(new_n527), .B2(new_n528), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n541), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n310), .A2(new_n615), .A3(new_n311), .A4(new_n630), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n529), .A2(new_n538), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n588), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n609), .A2(new_n611), .A3(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT35), .B(G107), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G9));
  OR2_X1    g451(.A1(new_n422), .A2(new_n423), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n386), .A2(KEYINPUT36), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n435), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n434), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n317), .A2(new_n591), .A3(new_n597), .A4(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT99), .B(KEYINPUT37), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G110), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n644), .B(new_n646), .ZN(G12));
  AOI221_X4 g461(.A(new_n613), .B1(new_n434), .B2(new_n642), .C1(new_n294), .C2(new_n309), .ZN(new_n648));
  INV_X1    g462(.A(G900), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n189), .B1(new_n193), .B2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n630), .A2(new_n538), .A3(new_n529), .A4(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n652), .A2(new_n589), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n648), .A2(new_n383), .A3(new_n607), .A4(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G128), .ZN(G30));
  NOR2_X1   g469(.A1(new_n544), .A2(new_n589), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n310), .B(KEYINPUT38), .Z(new_n657));
  INV_X1    g471(.A(new_n374), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n347), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n659), .A2(KEYINPUT100), .A3(new_n363), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n354), .ZN(new_n661));
  AOI21_X1  g475(.A(KEYINPUT100), .B1(new_n659), .B2(new_n363), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n274), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(G472), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n664), .A2(new_n371), .A3(new_n372), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NOR4_X1   g480(.A1(new_n657), .A2(new_n613), .A3(new_n643), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n650), .B(KEYINPUT39), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n484), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT101), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n670), .A2(KEYINPUT40), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n670), .A2(KEYINPUT40), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n656), .B(new_n667), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G143), .ZN(G45));
  NAND3_X1  g488(.A1(new_n543), .A2(new_n624), .A3(new_n651), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n648), .A2(new_n383), .A3(new_n607), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G146), .ZN(G48));
  AOI22_X1  g492(.A1(new_n461), .A2(new_n465), .B1(new_n599), .B2(new_n475), .ZN(new_n679));
  OAI21_X1  g493(.A(G469), .B1(new_n679), .B2(G902), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n680), .A2(new_n442), .A3(new_n606), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n681), .A2(new_n383), .A3(new_n437), .ZN(new_n682));
  INV_X1    g496(.A(new_n625), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT41), .B(G113), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G15));
  NAND2_X1  g500(.A1(new_n682), .A2(new_n634), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G116), .ZN(G18));
  NAND3_X1  g502(.A1(new_n310), .A2(new_n311), .A3(new_n643), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n680), .A2(new_n442), .A3(new_n606), .ZN(new_n690));
  NOR4_X1   g504(.A1(new_n689), .A2(new_n690), .A3(new_n590), .A4(new_n194), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n383), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G119), .ZN(G21));
  NAND2_X1  g507(.A1(new_n658), .A2(new_n359), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n363), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n355), .A2(new_n695), .A3(new_n366), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n696), .A2(new_n368), .A3(new_n274), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n368), .B1(new_n367), .B2(new_n274), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n437), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n700), .A2(new_n690), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n614), .A2(new_n656), .A3(new_n615), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G122), .ZN(G24));
  NOR3_X1   g518(.A1(new_n675), .A2(new_n697), .A3(new_n698), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n648), .A2(new_n705), .A3(new_n681), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G125), .ZN(G27));
  NAND2_X1  g521(.A1(new_n371), .A2(KEYINPUT102), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n382), .A2(new_n372), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT102), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n369), .A2(new_n710), .A3(new_n370), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n708), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n294), .A2(new_n309), .A3(new_n311), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n484), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n712), .A2(new_n714), .A3(new_n437), .A4(new_n676), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n294), .A2(new_n309), .A3(new_n311), .ZN(new_n716));
  AND4_X1   g530(.A1(new_n383), .A2(new_n607), .A3(new_n716), .A4(new_n437), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n675), .A2(KEYINPUT42), .ZN(new_n718));
  AOI22_X1  g532(.A1(new_n715), .A2(KEYINPUT42), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G131), .ZN(G33));
  NAND2_X1  g534(.A1(new_n717), .A2(new_n653), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G134), .ZN(G36));
  NAND3_X1  g536(.A1(new_n632), .A2(new_n542), .A3(new_n624), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT43), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(new_n596), .A3(new_n643), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT105), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n602), .A2(KEYINPUT45), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n602), .A2(KEYINPUT45), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n731), .A2(G469), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n482), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT46), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(KEYINPUT103), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n733), .A2(KEYINPUT46), .A3(new_n482), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT103), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n734), .A2(new_n739), .A3(new_n735), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n737), .A2(new_n606), .A3(new_n738), .A4(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT104), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n742), .B1(new_n726), .B2(new_n727), .ZN(new_n743));
  INV_X1    g557(.A(new_n668), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n741), .A2(new_n743), .A3(new_n442), .A4(new_n744), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n726), .A2(new_n742), .A3(new_n727), .ZN(new_n746));
  NOR4_X1   g560(.A1(new_n730), .A2(new_n745), .A3(new_n746), .A4(new_n713), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n321), .ZN(G39));
  NAND2_X1  g562(.A1(new_n741), .A2(new_n442), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT47), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n383), .A2(new_n437), .A3(new_n675), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n751), .A2(KEYINPUT106), .A3(new_n716), .A4(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n749), .A2(new_n750), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT47), .B1(new_n741), .B2(new_n442), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n716), .B(new_n752), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT106), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n753), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(KEYINPUT107), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G140), .ZN(G42));
  AND2_X1   g575(.A1(new_n680), .A2(new_n606), .ZN(new_n762));
  XOR2_X1   g576(.A(new_n762), .B(KEYINPUT49), .Z(new_n763));
  NOR3_X1   g577(.A1(new_n763), .A2(new_n665), .A3(new_n723), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n657), .A2(new_n437), .A3(new_n442), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n312), .A3(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n543), .A2(new_n624), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT108), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n588), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n582), .A2(new_n587), .A3(KEYINPUT108), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n768), .B1(new_n772), .B2(new_n543), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n317), .A2(new_n609), .A3(new_n611), .A4(new_n773), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n774), .A2(new_n644), .A3(new_n592), .ZN(new_n775));
  INV_X1    g589(.A(new_n643), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n529), .A2(new_n538), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT91), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n539), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n515), .A2(new_n526), .A3(KEYINPUT91), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT20), .B1(new_n781), .B2(new_n485), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n777), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n783), .A2(KEYINPUT109), .A3(new_n772), .A4(new_n651), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT109), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n582), .A2(new_n587), .A3(KEYINPUT108), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT108), .B1(new_n582), .B2(new_n587), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n785), .B1(new_n652), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n784), .A2(new_n383), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n699), .A2(new_n676), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n776), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  AOI22_X1  g606(.A1(new_n792), .A2(new_n714), .B1(new_n653), .B2(new_n717), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n654), .A2(new_n677), .A3(new_n706), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n665), .A2(new_n776), .A3(new_n651), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n607), .A2(new_n614), .A3(new_n656), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g611(.A(KEYINPUT52), .B1(new_n794), .B2(new_n797), .ZN(new_n798));
  AND4_X1   g612(.A1(new_n383), .A2(new_n607), .A3(new_n614), .A4(new_n643), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n689), .A2(new_n690), .ZN(new_n800));
  AOI22_X1  g614(.A1(new_n799), .A2(new_n653), .B1(new_n800), .B2(new_n705), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n795), .A2(new_n796), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n801), .A2(new_n802), .A3(new_n677), .A4(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n775), .A2(new_n793), .A3(new_n798), .A4(new_n804), .ZN(new_n805));
  AOI22_X1  g619(.A1(new_n691), .A2(new_n383), .B1(new_n682), .B2(new_n634), .ZN(new_n806));
  AOI22_X1  g620(.A1(new_n683), .A2(new_n682), .B1(new_n701), .B2(new_n702), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n719), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n767), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT110), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n804), .A2(new_n798), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n793), .A2(new_n592), .A3(new_n644), .A4(new_n774), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n719), .A2(new_n806), .A3(KEYINPUT53), .A4(new_n807), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n810), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  NOR4_X1   g630(.A1(new_n811), .A2(new_n812), .A3(new_n814), .A4(KEYINPUT110), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n809), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OR2_X1    g632(.A1(new_n818), .A2(KEYINPUT54), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n725), .A2(new_n189), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n690), .A2(new_n713), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(KEYINPUT112), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n712), .A2(new_n437), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n825), .B(KEYINPUT48), .Z(new_n826));
  NAND4_X1  g640(.A1(new_n666), .A2(new_n821), .A3(new_n437), .A4(new_n189), .ZN(new_n827));
  OAI211_X1 g641(.A(G952), .B(new_n188), .C1(new_n827), .C2(new_n768), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n820), .A2(new_n614), .A3(new_n701), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n813), .A2(new_n815), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n809), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT54), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n819), .A2(new_n829), .A3(new_n830), .A4(new_n833), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n820), .A2(new_n437), .A3(new_n699), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n716), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n754), .A2(new_n755), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n762), .A2(new_n441), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT113), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n836), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n841), .B1(new_n840), .B2(new_n839), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n681), .A2(KEYINPUT111), .A3(new_n613), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT111), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n844), .B1(new_n690), .B2(new_n311), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n835), .A2(new_n657), .A3(new_n843), .A4(new_n845), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT50), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n823), .A2(new_n643), .A3(new_n699), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n827), .A2(new_n543), .A3(new_n624), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n842), .A2(KEYINPUT51), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n839), .A2(new_n716), .A3(new_n835), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT51), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n834), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(G952), .A2(G953), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n766), .B1(new_n854), .B2(new_n855), .ZN(G75));
  NAND3_X1  g670(.A1(new_n818), .A2(G210), .A3(G902), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT115), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT56), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n818), .A2(KEYINPUT115), .A3(G210), .A4(G902), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n300), .B(new_n224), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(KEYINPUT114), .ZN(new_n864));
  XOR2_X1   g678(.A(new_n864), .B(KEYINPUT55), .Z(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n862), .A2(KEYINPUT116), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT116), .B1(new_n862), .B2(new_n866), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n857), .A2(new_n860), .A3(new_n865), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n188), .A2(G952), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n867), .A2(new_n868), .A3(new_n872), .ZN(G51));
  INV_X1    g687(.A(KEYINPUT117), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n818), .A2(KEYINPUT54), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n819), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n818), .A2(KEYINPUT117), .A3(KEYINPUT54), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n482), .B(KEYINPUT57), .Z(new_n878));
  NAND3_X1  g692(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n604), .ZN(new_n880));
  INV_X1    g694(.A(new_n808), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT53), .B1(new_n813), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n831), .A2(KEYINPUT110), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n813), .A2(new_n810), .A3(new_n815), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OR3_X1    g699(.A1(new_n885), .A2(new_n274), .A3(new_n733), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n870), .B1(new_n880), .B2(new_n886), .ZN(G54));
  NAND4_X1  g701(.A1(new_n818), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT118), .ZN(new_n889));
  INV_X1    g703(.A(new_n781), .ZN(new_n890));
  OR3_X1    g704(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n870), .B1(new_n888), .B2(new_n890), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n889), .B1(new_n888), .B2(new_n890), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(G60));
  XNOR2_X1  g708(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n580), .A2(new_n274), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n895), .B(new_n896), .Z(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n898), .B1(new_n819), .B2(new_n833), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n617), .A2(new_n620), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n871), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n876), .A2(new_n877), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n900), .A2(new_n897), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(G63));
  NAND2_X1  g718(.A1(G217), .A2(G902), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT60), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n640), .A2(new_n641), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT120), .ZN(new_n908));
  OR3_X1    g722(.A1(new_n885), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n424), .A2(new_n426), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n910), .B1(new_n885), .B2(new_n906), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n909), .A2(new_n871), .A3(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n912), .B(new_n913), .ZN(G66));
  INV_X1    g728(.A(G224), .ZN(new_n915));
  OAI21_X1  g729(.A(G953), .B1(new_n191), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n775), .A2(new_n807), .A3(new_n806), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n916), .B1(new_n918), .B2(G953), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n271), .B(new_n272), .C1(G898), .C2(new_n188), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n919), .B(new_n920), .ZN(G69));
  NOR2_X1   g735(.A1(new_n339), .A2(new_n344), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n521), .A2(new_n522), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT121), .Z(new_n924));
  XNOR2_X1  g738(.A(new_n922), .B(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(G900), .A2(G953), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n719), .A2(new_n721), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n927), .A2(KEYINPUT124), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n927), .A2(KEYINPUT124), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n747), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n794), .B(KEYINPUT123), .Z(new_n931));
  NOR2_X1   g745(.A1(new_n749), .A2(new_n668), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n932), .A2(new_n614), .A3(new_n656), .A4(new_n824), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n759), .A2(new_n930), .A3(new_n931), .A4(new_n933), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n925), .B(new_n926), .C1(new_n934), .C2(G953), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n673), .A2(new_n931), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT62), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n673), .A2(new_n931), .A3(KEYINPUT62), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n747), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n670), .A2(new_n438), .A3(new_n716), .A4(new_n773), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n759), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n942), .A2(new_n188), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n925), .B(KEYINPUT122), .Z(new_n944));
  OAI21_X1  g758(.A(new_n935), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n946), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n935), .B(new_n948), .C1(new_n943), .C2(new_n944), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n947), .A2(new_n949), .ZN(G72));
  NAND4_X1  g764(.A1(new_n759), .A2(new_n940), .A3(new_n918), .A4(new_n941), .ZN(new_n951));
  XOR2_X1   g765(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n952));
  NOR2_X1   g766(.A1(new_n368), .A2(new_n274), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT126), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n951), .A2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT127), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n345), .A2(new_n347), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n951), .A2(KEYINPUT127), .A3(new_n955), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n958), .A2(new_n353), .A3(new_n959), .A4(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n955), .B1(new_n934), .B2(new_n917), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n959), .A2(new_n353), .ZN(new_n963));
  INV_X1    g777(.A(new_n380), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n354), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n954), .B1(new_n809), .B2(new_n831), .ZN(new_n966));
  AOI22_X1  g780(.A1(new_n962), .A2(new_n963), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n961), .A2(new_n967), .A3(new_n871), .ZN(G57));
endmodule


