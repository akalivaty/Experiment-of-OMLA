//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 1 1 0 0 0 0 1 1 1 1 0 1 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 0 1 0 0 0 1 0 1 0 1 0 0 1 0 0 0 0 0 0 1 0 0 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n450, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n605, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1207, new_n1208;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  INV_X1    g024(.A(G2106), .ZN(new_n450));
  NOR2_X1   g025(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT66), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT67), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT68), .Z(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI22_X1  g035(.A1(new_n454), .A2(new_n450), .B1(new_n460), .B2(new_n456), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT69), .Z(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT70), .Z(G319));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT71), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT71), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(new_n467), .A3(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n469), .A2(G137), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G101), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(G2105), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n467), .A2(G2104), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n470), .A2(new_n476), .A3(G125), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n474), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n467), .A2(G2104), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n485), .B1(new_n465), .B2(new_n468), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G124), .ZN(new_n488));
  INV_X1    g063(.A(G136), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n486), .A2(new_n475), .ZN(new_n490));
  OAI221_X1 g065(.A(new_n484), .B1(new_n487), .B2(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT72), .ZN(new_n492));
  XNOR2_X1  g067(.A(new_n492), .B(KEYINPUT73), .ZN(G162));
  AND2_X1   g068(.A1(KEYINPUT4), .A2(G138), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n469), .A2(new_n475), .A3(new_n470), .A4(new_n494), .ZN(new_n495));
  AND3_X1   g070(.A1(new_n475), .A2(G102), .A3(G2104), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n470), .A2(new_n476), .A3(G138), .A4(new_n475), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(G114), .A2(G2104), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n501), .B1(new_n486), .B2(G126), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n495), .B(new_n499), .C1(new_n502), .C2(new_n475), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(KEYINPUT74), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT74), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT5), .A3(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT75), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n510), .A2(KEYINPUT75), .A3(new_n511), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G88), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  OAI21_X1  g094(.A(KEYINPUT76), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n511), .A2(G543), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G50), .ZN(new_n523));
  OR3_X1    g098(.A1(new_n518), .A2(KEYINPUT76), .A3(new_n519), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n517), .A2(new_n520), .A3(new_n523), .A4(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  NAND3_X1  g101(.A1(new_n510), .A2(G63), .A3(G651), .ZN(new_n527));
  INV_X1    g102(.A(G51), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n528), .B2(new_n521), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT77), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n529), .B(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n516), .A2(G89), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n507), .A2(new_n509), .ZN(new_n538));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g115(.A(KEYINPUT78), .B(G52), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n540), .A2(G651), .B1(new_n522), .B2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n514), .A2(new_n515), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  AOI22_X1  g121(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n519), .ZN(new_n548));
  INV_X1    g123(.A(G43), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n549), .B2(new_n521), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n550), .B1(new_n516), .B2(G81), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND3_X1  g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(KEYINPUT8), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n555), .A2(KEYINPUT8), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n554), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  XOR2_X1   g133(.A(new_n558), .B(KEYINPUT79), .Z(G188));
  NAND3_X1  g134(.A1(new_n511), .A2(G53), .A3(G543), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT9), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n514), .A2(G91), .A3(new_n515), .ZN(new_n562));
  AND2_X1   g137(.A1(new_n510), .A2(G65), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  XOR2_X1   g139(.A(new_n564), .B(KEYINPUT80), .Z(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n561), .A2(new_n562), .A3(new_n566), .ZN(G299));
  INV_X1    g142(.A(KEYINPUT81), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n516), .A2(new_n568), .A3(G87), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n510), .A2(G74), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n570), .A2(G651), .B1(new_n522), .B2(G49), .ZN(new_n571));
  INV_X1    g146(.A(G87), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT81), .B1(new_n544), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n569), .A2(new_n571), .A3(new_n573), .ZN(G288));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n538), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n577), .A2(G651), .B1(G48), .B2(new_n522), .ZN(new_n578));
  INV_X1    g153(.A(G86), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n579), .B2(new_n544), .ZN(G305));
  NAND2_X1  g155(.A1(new_n522), .A2(G47), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G85), .ZN(new_n583));
  OAI221_X1 g158(.A(new_n581), .B1(new_n519), .B2(new_n582), .C1(new_n544), .C2(new_n583), .ZN(new_n584));
  XOR2_X1   g159(.A(new_n584), .B(KEYINPUT82), .Z(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G290));
  NAND2_X1  g161(.A1(G301), .A2(G868), .ZN(new_n587));
  INV_X1    g162(.A(G92), .ZN(new_n588));
  OAI21_X1  g163(.A(KEYINPUT10), .B1(new_n544), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(G79), .A2(G543), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT83), .ZN(new_n591));
  INV_X1    g166(.A(G66), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n538), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n593), .A2(G651), .B1(G54), .B2(new_n522), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n514), .A2(new_n595), .A3(G92), .A4(new_n515), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n589), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n587), .B1(new_n598), .B2(G868), .ZN(G284));
  OAI21_X1  g174(.A(new_n587), .B1(new_n598), .B2(G868), .ZN(G321));
  NAND2_X1  g175(.A1(G286), .A2(G868), .ZN(new_n601));
  INV_X1    g176(.A(G299), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(G868), .B2(new_n602), .ZN(G297));
  OAI21_X1  g178(.A(new_n601), .B1(G868), .B2(new_n602), .ZN(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n598), .B1(new_n605), .B2(G860), .ZN(G148));
  OAI21_X1  g181(.A(KEYINPUT84), .B1(new_n551), .B2(G868), .ZN(new_n607));
  OAI21_X1  g182(.A(G868), .B1(new_n597), .B2(G559), .ZN(new_n608));
  MUX2_X1   g183(.A(KEYINPUT84), .B(new_n607), .S(new_n608), .Z(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g185(.A(new_n487), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G123), .ZN(new_n612));
  INV_X1    g187(.A(new_n490), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G135), .ZN(new_n614));
  NOR2_X1   g189(.A1(G99), .A2(G2105), .ZN(new_n615));
  OAI21_X1  g190(.A(G2104), .B1(new_n475), .B2(G111), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n612), .B(new_n614), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(G2096), .Z(new_n618));
  NAND3_X1  g193(.A1(new_n475), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT85), .B(G2100), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n618), .A2(new_n623), .ZN(G156));
  XNOR2_X1  g199(.A(G2443), .B(G2446), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2435), .ZN(new_n628));
  XOR2_X1   g203(.A(G2427), .B(G2438), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(KEYINPUT14), .ZN(new_n631));
  XOR2_X1   g206(.A(G2451), .B(G2454), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n631), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G1341), .B(G1348), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n634), .A2(new_n635), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n626), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n634), .A2(new_n635), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n640), .A2(new_n636), .A3(new_n625), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n639), .A2(new_n641), .A3(G14), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(G401));
  XOR2_X1   g218(.A(G2067), .B(G2678), .Z(new_n644));
  XNOR2_X1  g219(.A(G2084), .B(G2090), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(new_n647), .A3(KEYINPUT17), .ZN(new_n648));
  INV_X1    g223(.A(KEYINPUT18), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G2072), .B(G2078), .Z(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(new_n646), .B2(KEYINPUT18), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n650), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2096), .B(G2100), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT86), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n653), .B(new_n655), .ZN(G227));
  XNOR2_X1  g231(.A(G1991), .B(G1996), .ZN(new_n657));
  INV_X1    g232(.A(G1981), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1956), .B(G2474), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT87), .ZN(new_n662));
  XOR2_X1   g237(.A(G1961), .B(G1966), .Z(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT88), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1971), .B(G1976), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT20), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n662), .A2(new_n663), .ZN(new_n672));
  AOI22_X1  g247(.A1(new_n670), .A2(new_n671), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n666), .A2(KEYINPUT20), .A3(new_n669), .ZN(new_n674));
  INV_X1    g249(.A(new_n672), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n675), .A2(new_n668), .A3(new_n664), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n673), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g255(.A1(new_n673), .A2(new_n678), .A3(new_n674), .A4(new_n676), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n660), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT89), .B(G1986), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n680), .A2(new_n660), .A3(new_n681), .ZN(new_n685));
  AND3_X1   g260(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n684), .B1(new_n683), .B2(new_n685), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(G229));
  NAND2_X1  g264(.A1(KEYINPUT93), .A2(KEYINPUT36), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT34), .ZN(new_n691));
  INV_X1    g266(.A(G288), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G16), .ZN(new_n693));
  OR2_X1    g268(.A1(G16), .A2(G23), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT33), .B(G1976), .Z(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(G303), .A2(G16), .ZN(new_n699));
  INV_X1    g274(.A(G22), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(G16), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G1971), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n693), .A2(new_n694), .A3(new_n696), .ZN(new_n703));
  INV_X1    g278(.A(G1971), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n699), .B(new_n704), .C1(G16), .C2(new_n700), .ZN(new_n705));
  NAND4_X1  g280(.A1(new_n698), .A2(new_n702), .A3(new_n703), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT32), .B(G1981), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT92), .ZN(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n516), .A2(G86), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(new_n578), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n709), .A2(G6), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n708), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n712), .B1(G305), .B2(G16), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(KEYINPUT92), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n707), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n713), .A2(new_n715), .A3(new_n707), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n691), .B1(new_n706), .B2(new_n719), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n702), .A2(new_n705), .ZN(new_n721));
  INV_X1    g296(.A(new_n718), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n722), .A2(new_n716), .ZN(new_n723));
  AND3_X1   g298(.A1(new_n693), .A2(new_n694), .A3(new_n696), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n696), .B1(new_n693), .B2(new_n694), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n721), .A2(new_n723), .A3(new_n726), .A4(KEYINPUT34), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n720), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n611), .A2(G119), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n613), .A2(G131), .ZN(new_n730));
  NOR2_X1   g305(.A1(G95), .A2(G2105), .ZN(new_n731));
  OAI21_X1  g306(.A(G2104), .B1(new_n475), .B2(G107), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n729), .B(new_n730), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G29), .ZN(new_n734));
  INV_X1    g309(.A(G25), .ZN(new_n735));
  OAI21_X1  g310(.A(KEYINPUT90), .B1(new_n735), .B2(G29), .ZN(new_n736));
  OR3_X1    g311(.A1(new_n735), .A2(KEYINPUT90), .A3(G29), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n734), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT35), .B(G1991), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n709), .A2(G24), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n585), .B2(new_n709), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT91), .B(G1986), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n728), .A2(new_n741), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n746), .A2(KEYINPUT94), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT94), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n740), .B1(new_n720), .B2(new_n727), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(new_n745), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n690), .B1(new_n747), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n746), .A2(KEYINPUT94), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n749), .A2(new_n748), .A3(new_n745), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n752), .A2(KEYINPUT93), .A3(KEYINPUT36), .A4(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT29), .ZN(new_n755));
  NAND2_X1  g330(.A1(G162), .A2(G29), .ZN(new_n756));
  NOR2_X1   g331(.A1(G29), .A2(G35), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n755), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  AOI211_X1 g335(.A(KEYINPUT29), .B(new_n757), .C1(G162), .C2(G29), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n760), .A2(new_n762), .A3(G2090), .ZN(new_n763));
  INV_X1    g338(.A(G2090), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n759), .B2(new_n761), .ZN(new_n765));
  INV_X1    g340(.A(G29), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G33), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT25), .Z(new_n769));
  INV_X1    g344(.A(G139), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n470), .A2(new_n476), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n771), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n772));
  OAI221_X1 g347(.A(new_n769), .B1(new_n490), .B2(new_n770), .C1(new_n475), .C2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT96), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n767), .B1(new_n775), .B2(new_n766), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(G2072), .Z(new_n777));
  NAND3_X1  g352(.A1(new_n763), .A2(new_n765), .A3(new_n777), .ZN(new_n778));
  AND2_X1   g353(.A1(KEYINPUT24), .A2(G34), .ZN(new_n779));
  NOR2_X1   g354(.A1(KEYINPUT24), .A2(G34), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n766), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n481), .B2(new_n766), .ZN(new_n782));
  INV_X1    g357(.A(G2084), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT31), .ZN(new_n784));
  OAI22_X1  g359(.A1(new_n782), .A2(new_n783), .B1(new_n784), .B2(G11), .ZN(new_n785));
  NOR2_X1   g360(.A1(G5), .A2(G16), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G171), .B2(G16), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n787), .A2(G1961), .ZN(new_n788));
  AOI211_X1 g363(.A(new_n785), .B(new_n788), .C1(new_n784), .C2(G11), .ZN(new_n789));
  INV_X1    g364(.A(G27), .ZN(new_n790));
  OAI21_X1  g365(.A(KEYINPUT100), .B1(new_n790), .B2(G29), .ZN(new_n791));
  OR3_X1    g366(.A1(new_n790), .A2(KEYINPUT100), .A3(G29), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n791), .B(new_n792), .C1(G164), .C2(new_n766), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n793), .A2(G2078), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n617), .A2(new_n766), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT30), .B(G28), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n787), .A2(G1961), .B1(new_n766), .B2(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n789), .A2(new_n794), .A3(new_n795), .A4(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(G286), .A2(new_n709), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT99), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(KEYINPUT99), .B1(G16), .B2(G21), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n803), .A2(G1966), .B1(new_n783), .B2(new_n782), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n709), .A2(G4), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n598), .B2(new_n709), .ZN(new_n806));
  INV_X1    g381(.A(G1348), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n804), .B(new_n808), .C1(G1966), .C2(new_n803), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n709), .A2(G19), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n551), .B2(new_n709), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(G1341), .Z(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G2078), .B2(new_n793), .ZN(new_n813));
  NOR4_X1   g388(.A1(new_n778), .A2(new_n798), .A3(new_n809), .A4(new_n813), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n709), .A2(KEYINPUT23), .A3(G20), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT23), .ZN(new_n816));
  INV_X1    g391(.A(G20), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(G16), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n815), .B(new_n818), .C1(new_n602), .C2(new_n709), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT101), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G1956), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n751), .A2(new_n754), .A3(new_n814), .A4(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n766), .A2(G26), .ZN(new_n823));
  OR2_X1    g398(.A1(G104), .A2(G2105), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n824), .B(G2104), .C1(G116), .C2(new_n475), .ZN(new_n825));
  INV_X1    g400(.A(G128), .ZN(new_n826));
  INV_X1    g401(.A(G140), .ZN(new_n827));
  OAI221_X1 g402(.A(new_n825), .B1(new_n487), .B2(new_n826), .C1(new_n827), .C2(new_n490), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT95), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n829), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n823), .B1(new_n833), .B2(new_n766), .ZN(new_n834));
  MUX2_X1   g409(.A(new_n823), .B(new_n834), .S(KEYINPUT28), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(G2067), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n613), .A2(G141), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT97), .ZN(new_n838));
  NAND3_X1  g413(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT26), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n475), .A2(G105), .A3(G2104), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT98), .ZN(new_n842));
  AOI211_X1 g417(.A(new_n840), .B(new_n842), .C1(new_n611), .C2(G129), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n838), .A2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(G29), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(G29), .B2(G32), .ZN(new_n847));
  XNOR2_X1  g422(.A(KEYINPUT27), .B(G1996), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  NOR3_X1   g424(.A1(new_n822), .A2(new_n836), .A3(new_n849), .ZN(G311));
  AND3_X1   g425(.A1(new_n751), .A2(new_n754), .A3(new_n814), .ZN(new_n851));
  INV_X1    g426(.A(new_n836), .ZN(new_n852));
  INV_X1    g427(.A(new_n849), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .A4(new_n821), .ZN(G150));
  AOI22_X1  g429(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n855), .A2(new_n519), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n514), .A2(G93), .A3(new_n515), .ZN(new_n857));
  XOR2_X1   g432(.A(KEYINPUT102), .B(G55), .Z(new_n858));
  NAND2_X1  g433(.A1(new_n522), .A2(new_n858), .ZN(new_n859));
  AND3_X1   g434(.A1(new_n857), .A2(KEYINPUT103), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(KEYINPUT103), .B1(new_n857), .B2(new_n859), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n856), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(G860), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT37), .Z(new_n864));
  NOR2_X1   g439(.A1(new_n597), .A2(new_n605), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT38), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT39), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n862), .A2(KEYINPUT104), .ZN(new_n868));
  INV_X1    g443(.A(new_n551), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT104), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n870), .B(new_n856), .C1(new_n860), .C2(new_n861), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n868), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n862), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n873), .A2(new_n870), .A3(new_n551), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n867), .B(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n864), .B1(new_n876), .B2(G860), .ZN(G145));
  XNOR2_X1  g452(.A(new_n617), .B(new_n481), .ZN(new_n878));
  XNOR2_X1  g453(.A(KEYINPUT105), .B(KEYINPUT106), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(G162), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n832), .B(G164), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n775), .B(new_n844), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n883), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(G142), .ZN(new_n887));
  NOR2_X1   g462(.A1(G106), .A2(G2105), .ZN(new_n888));
  OAI21_X1  g463(.A(G2104), .B1(new_n475), .B2(G118), .ZN(new_n889));
  OAI22_X1  g464(.A1(new_n490), .A2(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n890), .B1(G130), .B2(new_n611), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(new_n620), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n892), .A2(new_n733), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n733), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(KEYINPUT107), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT107), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(new_n893), .B2(new_n894), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n886), .A2(new_n899), .ZN(new_n900));
  AOI22_X1  g475(.A1(new_n884), .A2(new_n885), .B1(new_n896), .B2(new_n898), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n881), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n886), .A2(new_n895), .ZN(new_n903));
  INV_X1    g478(.A(new_n881), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n903), .B(new_n904), .C1(new_n899), .C2(new_n886), .ZN(new_n905));
  INV_X1    g480(.A(G37), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n902), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g483(.A1(new_n597), .A2(G559), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n875), .B(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT108), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n597), .A2(new_n911), .A3(new_n602), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n911), .B1(new_n597), .B2(new_n602), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n597), .A2(new_n602), .ZN(new_n915));
  NOR3_X1   g490(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n910), .A2(new_n917), .ZN(new_n918));
  NOR3_X1   g493(.A1(new_n913), .A2(KEYINPUT109), .A3(new_n914), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT109), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n597), .A2(new_n602), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT108), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n920), .B1(new_n922), .B2(new_n912), .ZN(new_n923));
  OAI22_X1  g498(.A1(new_n919), .A2(new_n923), .B1(new_n602), .B2(new_n597), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT41), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n924), .A2(KEYINPUT110), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT110), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT109), .B1(new_n913), .B2(new_n914), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n922), .A2(new_n920), .A3(new_n912), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n915), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n927), .B1(new_n930), .B2(KEYINPUT41), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n916), .A2(KEYINPUT41), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n910), .A2(new_n926), .A3(new_n931), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n918), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT42), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT111), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n692), .A2(G303), .ZN(new_n937));
  NAND2_X1  g512(.A1(G166), .A2(G288), .ZN(new_n938));
  AOI21_X1  g513(.A(G305), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n937), .A2(new_n938), .A3(G305), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(new_n585), .A3(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n941), .ZN(new_n943));
  OAI21_X1  g518(.A(G290), .B1(new_n943), .B2(new_n939), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n934), .A2(new_n936), .A3(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n935), .A2(KEYINPUT111), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n945), .A2(new_n936), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n918), .A2(new_n933), .A3(new_n949), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n946), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n948), .B1(new_n946), .B2(new_n950), .ZN(new_n952));
  OAI21_X1  g527(.A(G868), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n953), .B1(G868), .B2(new_n873), .ZN(G295));
  OAI21_X1  g529(.A(new_n953), .B1(G868), .B2(new_n873), .ZN(G331));
  XNOR2_X1  g530(.A(G286), .B(G301), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n956), .A2(new_n872), .A3(new_n874), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n956), .B1(new_n874), .B2(new_n872), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n926), .A2(new_n960), .A3(new_n931), .A4(new_n932), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n916), .B1(new_n958), .B2(new_n959), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(G37), .B1(new_n963), .B2(new_n945), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n942), .A2(new_n944), .ZN(new_n965));
  XNOR2_X1  g540(.A(G286), .B(G171), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n875), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n967), .A2(KEYINPUT41), .A3(new_n957), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n916), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n924), .A2(new_n967), .A3(KEYINPUT41), .A4(new_n957), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n965), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n965), .A2(new_n969), .A3(KEYINPUT112), .A4(new_n970), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AND3_X1   g550(.A1(new_n964), .A2(new_n975), .A3(KEYINPUT43), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n961), .A2(new_n962), .A3(new_n965), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT43), .B1(new_n964), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT44), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT43), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n964), .A2(new_n975), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n981), .B1(new_n964), .B2(new_n977), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n979), .A2(new_n984), .ZN(G397));
  XNOR2_X1  g560(.A(G305), .B(G1981), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT49), .ZN(new_n987));
  OR2_X1    g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n987), .ZN(new_n989));
  INV_X1    g564(.A(G40), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n473), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n480), .ZN(new_n992));
  INV_X1    g567(.A(G1384), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n469), .A2(G126), .A3(new_n470), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n475), .B1(new_n994), .B2(new_n500), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n499), .A2(new_n495), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n993), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT115), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT115), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n999), .B(new_n993), .C1(new_n995), .C2(new_n996), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n992), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G8), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n988), .A2(new_n989), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1976), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1004), .A2(new_n1005), .A3(new_n692), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1006), .B1(G1981), .B2(G305), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n1003), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1000), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n999), .B1(new_n503), .B2(new_n993), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n992), .B1(KEYINPUT50), .B2(new_n997), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1012), .A2(new_n764), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT116), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT116), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1012), .A2(new_n1013), .A3(new_n1016), .A4(new_n764), .ZN(new_n1017));
  OAI211_X1 g592(.A(KEYINPUT45), .B(new_n993), .C1(new_n995), .C2(new_n996), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n473), .A2(new_n990), .A3(new_n479), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT45), .B1(new_n503), .B2(new_n993), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1022), .A2(G1971), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1015), .A2(new_n1017), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(G303), .A2(G8), .ZN(new_n1026));
  XOR2_X1   g601(.A(new_n1026), .B(KEYINPUT55), .Z(new_n1027));
  NAND3_X1  g602(.A1(new_n1025), .A2(G8), .A3(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n1028), .B(KEYINPUT117), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT52), .B1(G288), .B2(new_n1005), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n1030), .A2(KEYINPUT119), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n692), .A2(G1976), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1030), .A2(KEYINPUT119), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1031), .A2(new_n1003), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1019), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1035), .B(G8), .C1(new_n1005), .C2(G288), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n1036), .A2(KEYINPUT118), .A3(KEYINPUT52), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT118), .B1(new_n1036), .B2(KEYINPUT52), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1034), .B(new_n1004), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1008), .B1(new_n1029), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT62), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT45), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n998), .A2(new_n1042), .A3(new_n1000), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1020), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G1966), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT120), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT120), .ZN(new_n1048));
  AOI211_X1 g623(.A(new_n1048), .B(G1966), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT50), .B1(new_n998), .B2(new_n1000), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n997), .A2(KEYINPUT50), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n1019), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n1050), .A2(new_n1052), .A3(G2084), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n1047), .A2(new_n1049), .A3(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT51), .B1(new_n1054), .B2(G168), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1002), .B1(new_n1054), .B2(G168), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT51), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n1048), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1053), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1045), .A2(KEYINPUT120), .A3(new_n1046), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1060), .A2(new_n1061), .A3(G168), .A4(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1058), .B1(new_n1063), .B2(G8), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1041), .B1(new_n1057), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1039), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1027), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n998), .A2(KEYINPUT50), .A3(new_n1000), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n503), .A2(new_n1009), .A3(new_n993), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(new_n1019), .A3(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1071), .A2(G2090), .ZN(new_n1072));
  OAI21_X1  g647(.A(G8), .B1(new_n1072), .B2(new_n1023), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1068), .A2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1028), .A2(KEYINPUT117), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1023), .B1(new_n1014), .B2(KEYINPUT116), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1002), .B1(new_n1077), .B2(new_n1017), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1076), .B1(new_n1078), .B2(new_n1027), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1067), .B(new_n1074), .C1(new_n1075), .C2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1066), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(G2078), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1022), .A2(new_n1082), .ZN(new_n1083));
  XNOR2_X1  g658(.A(KEYINPUT123), .B(KEYINPUT53), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1082), .A2(KEYINPUT53), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1043), .A2(new_n1044), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G1961), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1088), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1085), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(G171), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1064), .B1(new_n1056), .B2(new_n1055), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1091), .B1(new_n1092), .B2(new_n1041), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1040), .B1(new_n1081), .B2(new_n1093), .ZN(new_n1094));
  XOR2_X1   g669(.A(KEYINPUT121), .B(G1956), .Z(new_n1095));
  NAND2_X1  g670(.A1(new_n1071), .A2(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT56), .B(G2072), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n1020), .A2(new_n1021), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1096), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT57), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n561), .A2(new_n562), .A3(new_n1103), .A4(new_n566), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1105), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1096), .A2(new_n1100), .A3(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1106), .A2(KEYINPUT61), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT61), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1107), .B1(new_n1096), .B2(new_n1100), .ZN(new_n1111));
  AOI211_X1 g686(.A(new_n1105), .B(new_n1099), .C1(new_n1071), .C2(new_n1095), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1110), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT58), .B(G1341), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1001), .A2(new_n1114), .ZN(new_n1115));
  NOR3_X1   g690(.A1(new_n1020), .A2(new_n1021), .A3(G1996), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n551), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT59), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1119), .B(new_n551), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1109), .A2(new_n1113), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1109), .A2(new_n1113), .A3(new_n1121), .A4(KEYINPUT122), .ZN(new_n1125));
  AOI21_X1  g700(.A(G1348), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1126));
  INV_X1    g701(.A(G2067), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1126), .B1(new_n1127), .B2(new_n1001), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1128), .A2(KEYINPUT60), .A3(new_n597), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n597), .B1(new_n1128), .B2(KEYINPUT60), .ZN(new_n1130));
  OAI22_X1  g705(.A1(new_n1129), .A2(new_n1130), .B1(KEYINPUT60), .B2(new_n1128), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1124), .A2(new_n1125), .A3(new_n1131), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1112), .A2(new_n1128), .A3(new_n597), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1133), .A2(new_n1111), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT54), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1091), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n997), .A2(new_n1042), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1138), .A2(new_n1018), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n477), .A2(new_n478), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n475), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n1141), .B2(new_n1140), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1139), .A2(new_n991), .A3(new_n1086), .A4(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1085), .A2(new_n1089), .A3(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1145), .A2(G171), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1136), .B1(new_n1137), .B2(new_n1146), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1085), .A2(new_n1089), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1148), .A2(KEYINPUT125), .A3(G301), .A4(new_n1087), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1136), .B1(new_n1145), .B2(G171), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT125), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1151), .B1(new_n1090), .B2(G171), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1149), .A2(new_n1150), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1147), .A2(new_n1153), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1080), .A2(new_n1154), .A3(new_n1092), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1135), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT63), .ZN(new_n1157));
  NOR3_X1   g732(.A1(new_n1054), .A2(new_n1002), .A3(G286), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1157), .B1(new_n1080), .B2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1078), .A2(new_n1027), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1161), .A2(new_n1157), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1029), .A2(new_n1158), .A3(new_n1067), .A4(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1094), .A2(new_n1156), .A3(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1138), .A2(new_n992), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n832), .B(new_n1127), .ZN(new_n1168));
  INV_X1    g743(.A(G1996), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n844), .B(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1167), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT114), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n733), .A2(new_n739), .ZN(new_n1173));
  AND2_X1   g748(.A1(new_n733), .A2(new_n739), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1166), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  AND2_X1   g750(.A1(new_n1172), .A2(new_n1175), .ZN(new_n1176));
  OR3_X1    g751(.A1(G290), .A2(G1986), .A3(new_n1167), .ZN(new_n1177));
  NAND3_X1  g752(.A1(G290), .A2(G1986), .A3(new_n1166), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1179), .B(KEYINPUT113), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n1176), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1165), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1167), .B1(new_n1168), .B2(new_n845), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1184));
  XOR2_X1   g759(.A(new_n1184), .B(KEYINPUT46), .Z(new_n1185));
  NOR2_X1   g760(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(KEYINPUT47), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n833), .A2(new_n1127), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1167), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1177), .B(KEYINPUT48), .ZN(new_n1191));
  AOI211_X1 g766(.A(new_n1187), .B(new_n1190), .C1(new_n1176), .C2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1182), .A2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g768(.A1(new_n462), .A2(G227), .ZN(new_n1195));
  NAND2_X1  g769(.A1(new_n642), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g770(.A(KEYINPUT126), .ZN(new_n1197));
  NAND2_X1  g771(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g772(.A1(new_n642), .A2(KEYINPUT126), .A3(new_n1195), .ZN(new_n1199));
  OAI211_X1 g773(.A(new_n1198), .B(new_n1199), .C1(new_n686), .C2(new_n687), .ZN(new_n1200));
  AND2_X1   g774(.A1(new_n1200), .A2(KEYINPUT127), .ZN(new_n1201));
  OAI21_X1  g775(.A(new_n907), .B1(new_n1200), .B2(KEYINPUT127), .ZN(new_n1202));
  NAND2_X1  g776(.A1(new_n964), .A2(new_n977), .ZN(new_n1203));
  NAND2_X1  g777(.A1(new_n1203), .A2(KEYINPUT43), .ZN(new_n1204));
  NAND3_X1  g778(.A1(new_n964), .A2(new_n975), .A3(new_n981), .ZN(new_n1205));
  AOI211_X1 g779(.A(new_n1201), .B(new_n1202), .C1(new_n1204), .C2(new_n1205), .ZN(G308));
  AOI21_X1  g780(.A(new_n1201), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1207));
  INV_X1    g781(.A(new_n1202), .ZN(new_n1208));
  NAND2_X1  g782(.A1(new_n1207), .A2(new_n1208), .ZN(G225));
endmodule


