

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594;

  XNOR2_X1 U320 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U321 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U322 ( .A(n327), .B(n326), .ZN(n375) );
  OR2_X1 U323 ( .A1(n572), .A2(n580), .ZN(n349) );
  OR2_X1 U324 ( .A1(n369), .A2(n368), .ZN(n370) );
  INV_X1 U325 ( .A(KEYINPUT71), .ZN(n315) );
  XNOR2_X1 U326 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U327 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U328 ( .A(n391), .B(n390), .ZN(n455) );
  XNOR2_X1 U329 ( .A(n318), .B(n317), .ZN(n319) );
  NAND2_X1 U330 ( .A1(n486), .A2(n485), .ZN(n496) );
  XNOR2_X1 U331 ( .A(n397), .B(n396), .ZN(n398) );
  INV_X1 U332 ( .A(KEYINPUT64), .ZN(n426) );
  XNOR2_X1 U333 ( .A(n427), .B(n426), .ZN(n579) );
  INV_X1 U334 ( .A(G36GAT), .ZN(n492) );
  XNOR2_X1 U335 ( .A(n463), .B(G190GAT), .ZN(n464) );
  XNOR2_X1 U336 ( .A(n492), .B(KEYINPUT108), .ZN(n493) );
  XNOR2_X1 U337 ( .A(n465), .B(n464), .ZN(G1351GAT) );
  XNOR2_X1 U338 ( .A(n494), .B(n493), .ZN(G1329GAT) );
  XOR2_X1 U339 ( .A(G50GAT), .B(G162GAT), .Z(n440) );
  XOR2_X1 U340 ( .A(G106GAT), .B(KEYINPUT76), .Z(n289) );
  XNOR2_X1 U341 ( .A(KEYINPUT10), .B(KEYINPUT77), .ZN(n288) );
  XNOR2_X1 U342 ( .A(n289), .B(n288), .ZN(n290) );
  XOR2_X1 U343 ( .A(n440), .B(n290), .Z(n294) );
  XOR2_X1 U344 ( .A(G29GAT), .B(G36GAT), .Z(n292) );
  XNOR2_X1 U345 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n291) );
  XNOR2_X1 U346 ( .A(n292), .B(n291), .ZN(n329) );
  XOR2_X1 U347 ( .A(G43GAT), .B(G134GAT), .Z(n447) );
  XNOR2_X1 U348 ( .A(n329), .B(n447), .ZN(n293) );
  XNOR2_X1 U349 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U350 ( .A(G85GAT), .B(G92GAT), .Z(n321) );
  XOR2_X1 U351 ( .A(n295), .B(n321), .Z(n297) );
  XNOR2_X1 U352 ( .A(G218GAT), .B(KEYINPUT9), .ZN(n296) );
  XNOR2_X1 U353 ( .A(n297), .B(n296), .ZN(n302) );
  XOR2_X1 U354 ( .A(G99GAT), .B(KEYINPUT11), .Z(n299) );
  NAND2_X1 U355 ( .A1(G232GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U356 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U357 ( .A(G190GAT), .B(n300), .Z(n301) );
  XNOR2_X1 U358 ( .A(n302), .B(n301), .ZN(n569) );
  INV_X1 U359 ( .A(n569), .ZN(n462) );
  INV_X1 U360 ( .A(KEYINPUT41), .ZN(n328) );
  INV_X1 U361 ( .A(KEYINPUT72), .ZN(n303) );
  NAND2_X1 U362 ( .A1(n303), .A2(G78GAT), .ZN(n306) );
  INV_X1 U363 ( .A(G78GAT), .ZN(n304) );
  NAND2_X1 U364 ( .A1(n304), .A2(KEYINPUT72), .ZN(n305) );
  NAND2_X1 U365 ( .A1(n306), .A2(n305), .ZN(n308) );
  XNOR2_X1 U366 ( .A(G148GAT), .B(G106GAT), .ZN(n307) );
  XNOR2_X1 U367 ( .A(n308), .B(n307), .ZN(n433) );
  XNOR2_X1 U368 ( .A(n433), .B(KEYINPUT32), .ZN(n309) );
  AND2_X1 U369 ( .A1(G230GAT), .A2(G233GAT), .ZN(n310) );
  NAND2_X1 U370 ( .A1(n309), .A2(n310), .ZN(n314) );
  INV_X1 U371 ( .A(n309), .ZN(n312) );
  INV_X1 U372 ( .A(n310), .ZN(n311) );
  NAND2_X1 U373 ( .A1(n312), .A2(n311), .ZN(n313) );
  NAND2_X1 U374 ( .A1(n314), .A2(n313), .ZN(n318) );
  XOR2_X1 U375 ( .A(G204GAT), .B(G64GAT), .Z(n399) );
  XNOR2_X1 U376 ( .A(n399), .B(KEYINPUT73), .ZN(n316) );
  XOR2_X1 U377 ( .A(G57GAT), .B(KEYINPUT13), .Z(n350) );
  XNOR2_X1 U378 ( .A(n319), .B(n350), .ZN(n327) );
  XNOR2_X1 U379 ( .A(G99GAT), .B(G120GAT), .ZN(n320) );
  XNOR2_X1 U380 ( .A(n320), .B(G71GAT), .ZN(n446) );
  XOR2_X1 U381 ( .A(n446), .B(n321), .Z(n325) );
  XOR2_X1 U382 ( .A(KEYINPUT74), .B(KEYINPUT31), .Z(n323) );
  XNOR2_X1 U383 ( .A(G176GAT), .B(KEYINPUT33), .ZN(n322) );
  XOR2_X1 U384 ( .A(n323), .B(n322), .Z(n324) );
  XNOR2_X1 U385 ( .A(n328), .B(n375), .ZN(n572) );
  XOR2_X1 U386 ( .A(n329), .B(G15GAT), .Z(n331) );
  NAND2_X1 U387 ( .A1(G229GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U388 ( .A(n331), .B(n330), .ZN(n347) );
  XOR2_X1 U389 ( .A(KEYINPUT66), .B(KEYINPUT30), .Z(n333) );
  XNOR2_X1 U390 ( .A(G169GAT), .B(KEYINPUT68), .ZN(n332) );
  XNOR2_X1 U391 ( .A(n333), .B(n332), .ZN(n345) );
  XOR2_X1 U392 ( .A(G113GAT), .B(G141GAT), .Z(n335) );
  XNOR2_X1 U393 ( .A(G50GAT), .B(G43GAT), .ZN(n334) );
  XNOR2_X1 U394 ( .A(n335), .B(n334), .ZN(n343) );
  XOR2_X1 U395 ( .A(G197GAT), .B(KEYINPUT70), .Z(n337) );
  XNOR2_X1 U396 ( .A(KEYINPUT67), .B(KEYINPUT29), .ZN(n336) );
  XNOR2_X1 U397 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U398 ( .A(KEYINPUT69), .B(G22GAT), .Z(n339) );
  XNOR2_X1 U399 ( .A(G1GAT), .B(G8GAT), .ZN(n338) );
  XNOR2_X1 U400 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U401 ( .A(n341), .B(n340), .Z(n342) );
  XNOR2_X1 U402 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U403 ( .A(n345), .B(n344), .Z(n346) );
  XNOR2_X1 U404 ( .A(n347), .B(n346), .ZN(n580) );
  XOR2_X1 U405 ( .A(KEYINPUT46), .B(KEYINPUT114), .Z(n348) );
  XNOR2_X1 U406 ( .A(n349), .B(n348), .ZN(n369) );
  XOR2_X1 U407 ( .A(G15GAT), .B(G127GAT), .Z(n448) );
  XOR2_X1 U408 ( .A(n350), .B(n448), .Z(n352) );
  NAND2_X1 U409 ( .A1(G231GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U410 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U411 ( .A(G211GAT), .B(KEYINPUT81), .Z(n354) );
  XNOR2_X1 U412 ( .A(KEYINPUT12), .B(KEYINPUT82), .ZN(n353) );
  XNOR2_X1 U413 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U414 ( .A(n356), .B(n355), .Z(n361) );
  XOR2_X1 U415 ( .A(KEYINPUT80), .B(KEYINPUT14), .Z(n358) );
  XNOR2_X1 U416 ( .A(KEYINPUT15), .B(KEYINPUT79), .ZN(n357) );
  XNOR2_X1 U417 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U418 ( .A(G183GAT), .B(n359), .ZN(n360) );
  XNOR2_X1 U419 ( .A(n361), .B(n360), .ZN(n365) );
  XOR2_X1 U420 ( .A(G8GAT), .B(KEYINPUT78), .Z(n395) );
  XOR2_X1 U421 ( .A(G22GAT), .B(G155GAT), .Z(n439) );
  XOR2_X1 U422 ( .A(n395), .B(n439), .Z(n363) );
  XNOR2_X1 U423 ( .A(G71GAT), .B(G64GAT), .ZN(n362) );
  XNOR2_X1 U424 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U425 ( .A(n365), .B(n364), .Z(n367) );
  XNOR2_X1 U426 ( .A(G1GAT), .B(G78GAT), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n367), .B(n366), .ZN(n588) );
  NAND2_X1 U428 ( .A1(n588), .A2(n462), .ZN(n368) );
  XNOR2_X1 U429 ( .A(n370), .B(KEYINPUT47), .ZN(n371) );
  XNOR2_X1 U430 ( .A(n371), .B(KEYINPUT115), .ZN(n379) );
  XNOR2_X1 U431 ( .A(KEYINPUT45), .B(KEYINPUT116), .ZN(n374) );
  XNOR2_X1 U432 ( .A(KEYINPUT36), .B(KEYINPUT104), .ZN(n372) );
  XNOR2_X1 U433 ( .A(n462), .B(n372), .ZN(n591) );
  NOR2_X1 U434 ( .A1(n588), .A2(n591), .ZN(n373) );
  XNOR2_X1 U435 ( .A(n374), .B(n373), .ZN(n377) );
  INV_X1 U436 ( .A(n580), .ZN(n558) );
  INV_X1 U437 ( .A(n375), .ZN(n469) );
  NOR2_X1 U438 ( .A1(n558), .A2(n469), .ZN(n376) );
  NAND2_X1 U439 ( .A1(n377), .A2(n376), .ZN(n378) );
  NAND2_X1 U440 ( .A1(n379), .A2(n378), .ZN(n381) );
  XOR2_X1 U441 ( .A(KEYINPUT48), .B(KEYINPUT117), .Z(n380) );
  XNOR2_X1 U442 ( .A(n381), .B(n380), .ZN(n543) );
  XOR2_X1 U443 ( .A(KEYINPUT21), .B(G211GAT), .Z(n383) );
  XNOR2_X1 U444 ( .A(G197GAT), .B(G218GAT), .ZN(n382) );
  XNOR2_X1 U445 ( .A(n383), .B(n382), .ZN(n437) );
  XOR2_X1 U446 ( .A(n437), .B(KEYINPUT96), .Z(n393) );
  XOR2_X1 U447 ( .A(KEYINPUT87), .B(KEYINPUT17), .Z(n385) );
  XNOR2_X1 U448 ( .A(KEYINPUT88), .B(KEYINPUT19), .ZN(n384) );
  XNOR2_X1 U449 ( .A(n385), .B(n384), .ZN(n387) );
  INV_X1 U450 ( .A(KEYINPUT18), .ZN(n386) );
  XNOR2_X1 U451 ( .A(n387), .B(n386), .ZN(n391) );
  XNOR2_X1 U452 ( .A(G169GAT), .B(G183GAT), .ZN(n389) );
  XNOR2_X1 U453 ( .A(G190GAT), .B(G176GAT), .ZN(n388) );
  XNOR2_X1 U454 ( .A(n455), .B(KEYINPUT97), .ZN(n392) );
  XNOR2_X1 U455 ( .A(n393), .B(n392), .ZN(n397) );
  XNOR2_X1 U456 ( .A(G36GAT), .B(G92GAT), .ZN(n394) );
  XNOR2_X1 U457 ( .A(n399), .B(n398), .ZN(n401) );
  NAND2_X1 U458 ( .A1(G226GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U459 ( .A(n401), .B(n400), .ZN(n476) );
  NAND2_X1 U460 ( .A1(n543), .A2(n476), .ZN(n403) );
  XOR2_X1 U461 ( .A(KEYINPUT54), .B(KEYINPUT122), .Z(n402) );
  XNOR2_X1 U462 ( .A(n403), .B(n402), .ZN(n425) );
  XOR2_X1 U463 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n405) );
  XNOR2_X1 U464 ( .A(KEYINPUT93), .B(KEYINPUT1), .ZN(n404) );
  XNOR2_X1 U465 ( .A(n405), .B(n404), .ZN(n409) );
  XOR2_X1 U466 ( .A(G155GAT), .B(KEYINPUT95), .Z(n407) );
  XNOR2_X1 U467 ( .A(G120GAT), .B(KEYINPUT94), .ZN(n406) );
  XNOR2_X1 U468 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U469 ( .A(n409), .B(n408), .ZN(n424) );
  XOR2_X1 U470 ( .A(G162GAT), .B(G85GAT), .Z(n411) );
  XNOR2_X1 U471 ( .A(G29GAT), .B(G134GAT), .ZN(n410) );
  XNOR2_X1 U472 ( .A(n411), .B(n410), .ZN(n416) );
  XNOR2_X1 U473 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n412) );
  XNOR2_X1 U474 ( .A(n412), .B(KEYINPUT2), .ZN(n434) );
  XOR2_X1 U475 ( .A(G57GAT), .B(n434), .Z(n414) );
  NAND2_X1 U476 ( .A1(G225GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U477 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U478 ( .A(n416), .B(n415), .Z(n422) );
  XNOR2_X1 U479 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n417), .B(KEYINPUT83), .ZN(n450) );
  XOR2_X1 U481 ( .A(G148GAT), .B(KEYINPUT4), .Z(n419) );
  XNOR2_X1 U482 ( .A(G1GAT), .B(G127GAT), .ZN(n418) );
  XNOR2_X1 U483 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U484 ( .A(n450), .B(n420), .ZN(n421) );
  XNOR2_X1 U485 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U486 ( .A(n424), .B(n423), .ZN(n533) );
  NAND2_X1 U487 ( .A1(n425), .A2(n533), .ZN(n427) );
  XOR2_X1 U488 ( .A(KEYINPUT90), .B(KEYINPUT92), .Z(n429) );
  XNOR2_X1 U489 ( .A(G204GAT), .B(KEYINPUT24), .ZN(n428) );
  XNOR2_X1 U490 ( .A(n429), .B(n428), .ZN(n444) );
  XOR2_X1 U491 ( .A(KEYINPUT23), .B(KEYINPUT91), .Z(n431) );
  NAND2_X1 U492 ( .A1(G228GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U493 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U494 ( .A(n432), .B(KEYINPUT22), .Z(n436) );
  XNOR2_X1 U495 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U496 ( .A(n436), .B(n435), .ZN(n438) );
  XOR2_X1 U497 ( .A(n438), .B(n437), .Z(n442) );
  XNOR2_X1 U498 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U499 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U500 ( .A(n444), .B(n443), .ZN(n482) );
  NAND2_X1 U501 ( .A1(n579), .A2(n482), .ZN(n445) );
  XNOR2_X1 U502 ( .A(n445), .B(KEYINPUT55), .ZN(n461) );
  XNOR2_X1 U503 ( .A(n447), .B(n446), .ZN(n449) );
  XNOR2_X1 U504 ( .A(n449), .B(n448), .ZN(n454) );
  XOR2_X1 U505 ( .A(n450), .B(KEYINPUT85), .Z(n452) );
  NAND2_X1 U506 ( .A1(G227GAT), .A2(G233GAT), .ZN(n451) );
  XNOR2_X1 U507 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U508 ( .A(n454), .B(n453), .Z(n460) );
  XOR2_X1 U509 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n457) );
  XNOR2_X1 U510 ( .A(KEYINPUT86), .B(KEYINPUT65), .ZN(n456) );
  XNOR2_X1 U511 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U512 ( .A(n455), .B(n458), .ZN(n459) );
  XNOR2_X1 U513 ( .A(n460), .B(n459), .ZN(n504) );
  NAND2_X1 U514 ( .A1(n461), .A2(n504), .ZN(n573) );
  NOR2_X1 U515 ( .A1(n462), .A2(n573), .ZN(n465) );
  INV_X1 U516 ( .A(KEYINPUT58), .ZN(n463) );
  NOR2_X1 U517 ( .A1(n588), .A2(n573), .ZN(n468) );
  INV_X1 U518 ( .A(G183GAT), .ZN(n466) );
  XNOR2_X1 U519 ( .A(n466), .B(KEYINPUT124), .ZN(n467) );
  XNOR2_X1 U520 ( .A(n468), .B(n467), .ZN(G1350GAT) );
  INV_X1 U521 ( .A(n476), .ZN(n535) );
  NOR2_X1 U522 ( .A1(n469), .A2(n580), .ZN(n470) );
  XNOR2_X1 U523 ( .A(n470), .B(KEYINPUT75), .ZN(n499) );
  NAND2_X1 U524 ( .A1(n504), .A2(n476), .ZN(n471) );
  XNOR2_X1 U525 ( .A(n471), .B(KEYINPUT98), .ZN(n472) );
  NAND2_X1 U526 ( .A1(n472), .A2(n482), .ZN(n474) );
  XNOR2_X1 U527 ( .A(KEYINPUT25), .B(KEYINPUT99), .ZN(n473) );
  XNOR2_X1 U528 ( .A(n474), .B(n473), .ZN(n479) );
  NOR2_X1 U529 ( .A1(n482), .A2(n504), .ZN(n475) );
  XNOR2_X1 U530 ( .A(n475), .B(KEYINPUT26), .ZN(n578) );
  XOR2_X1 U531 ( .A(n476), .B(KEYINPUT27), .Z(n481) );
  INV_X1 U532 ( .A(n481), .ZN(n477) );
  NAND2_X1 U533 ( .A1(n578), .A2(n477), .ZN(n478) );
  NAND2_X1 U534 ( .A1(n479), .A2(n478), .ZN(n480) );
  NAND2_X1 U535 ( .A1(n480), .A2(n533), .ZN(n486) );
  NOR2_X1 U536 ( .A1(n533), .A2(n481), .ZN(n542) );
  XOR2_X1 U537 ( .A(KEYINPUT28), .B(n482), .Z(n507) );
  XOR2_X1 U538 ( .A(n504), .B(KEYINPUT89), .Z(n483) );
  NOR2_X1 U539 ( .A1(n507), .A2(n483), .ZN(n484) );
  NAND2_X1 U540 ( .A1(n542), .A2(n484), .ZN(n485) );
  NAND2_X1 U541 ( .A1(n588), .A2(n496), .ZN(n487) );
  NOR2_X1 U542 ( .A1(n487), .A2(n591), .ZN(n488) );
  XNOR2_X1 U543 ( .A(n488), .B(KEYINPUT37), .ZN(n530) );
  NOR2_X1 U544 ( .A1(n499), .A2(n530), .ZN(n490) );
  XNOR2_X1 U545 ( .A(KEYINPUT106), .B(KEYINPUT38), .ZN(n489) );
  XNOR2_X1 U546 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U547 ( .A(KEYINPUT105), .B(n491), .ZN(n518) );
  NOR2_X1 U548 ( .A1(n535), .A2(n518), .ZN(n494) );
  NOR2_X1 U549 ( .A1(n588), .A2(n569), .ZN(n495) );
  XNOR2_X1 U550 ( .A(KEYINPUT16), .B(n495), .ZN(n497) );
  NAND2_X1 U551 ( .A1(n497), .A2(n496), .ZN(n498) );
  XNOR2_X1 U552 ( .A(n498), .B(KEYINPUT100), .ZN(n521) );
  NOR2_X1 U553 ( .A1(n521), .A2(n499), .ZN(n500) );
  XNOR2_X1 U554 ( .A(KEYINPUT101), .B(n500), .ZN(n508) );
  NOR2_X1 U555 ( .A1(n533), .A2(n508), .ZN(n501) );
  XOR2_X1 U556 ( .A(KEYINPUT34), .B(n501), .Z(n502) );
  XNOR2_X1 U557 ( .A(G1GAT), .B(n502), .ZN(G1324GAT) );
  NOR2_X1 U558 ( .A1(n535), .A2(n508), .ZN(n503) );
  XOR2_X1 U559 ( .A(G8GAT), .B(n503), .Z(G1325GAT) );
  INV_X1 U560 ( .A(n504), .ZN(n546) );
  NOR2_X1 U561 ( .A1(n546), .A2(n508), .ZN(n506) );
  XNOR2_X1 U562 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n505) );
  XNOR2_X1 U563 ( .A(n506), .B(n505), .ZN(G1326GAT) );
  INV_X1 U564 ( .A(n507), .ZN(n544) );
  NOR2_X1 U565 ( .A1(n544), .A2(n508), .ZN(n509) );
  XOR2_X1 U566 ( .A(G22GAT), .B(n509), .Z(n510) );
  XNOR2_X1 U567 ( .A(KEYINPUT102), .B(n510), .ZN(G1327GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT107), .B(KEYINPUT39), .Z(n512) );
  XNOR2_X1 U569 ( .A(G29GAT), .B(KEYINPUT103), .ZN(n511) );
  XNOR2_X1 U570 ( .A(n512), .B(n511), .ZN(n514) );
  NOR2_X1 U571 ( .A1(n533), .A2(n518), .ZN(n513) );
  XOR2_X1 U572 ( .A(n514), .B(n513), .Z(G1328GAT) );
  NOR2_X1 U573 ( .A1(n546), .A2(n518), .ZN(n516) );
  XNOR2_X1 U574 ( .A(KEYINPUT109), .B(KEYINPUT40), .ZN(n515) );
  XNOR2_X1 U575 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U576 ( .A(G43GAT), .B(n517), .ZN(G1330GAT) );
  NOR2_X1 U577 ( .A1(n544), .A2(n518), .ZN(n519) );
  XOR2_X1 U578 ( .A(G50GAT), .B(n519), .Z(G1331GAT) );
  INV_X1 U579 ( .A(n572), .ZN(n560) );
  NAND2_X1 U580 ( .A1(n560), .A2(n580), .ZN(n520) );
  XNOR2_X1 U581 ( .A(n520), .B(KEYINPUT110), .ZN(n531) );
  OR2_X1 U582 ( .A1(n521), .A2(n531), .ZN(n527) );
  NOR2_X1 U583 ( .A1(n533), .A2(n527), .ZN(n522) );
  XOR2_X1 U584 ( .A(n522), .B(KEYINPUT42), .Z(n523) );
  XNOR2_X1 U585 ( .A(G57GAT), .B(n523), .ZN(G1332GAT) );
  NOR2_X1 U586 ( .A1(n535), .A2(n527), .ZN(n524) );
  XOR2_X1 U587 ( .A(G64GAT), .B(n524), .Z(G1333GAT) );
  NOR2_X1 U588 ( .A1(n546), .A2(n527), .ZN(n526) );
  XNOR2_X1 U589 ( .A(G71GAT), .B(KEYINPUT111), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n526), .B(n525), .ZN(G1334GAT) );
  NOR2_X1 U591 ( .A1(n544), .A2(n527), .ZN(n529) );
  XNOR2_X1 U592 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n529), .B(n528), .ZN(G1335GAT) );
  NOR2_X1 U594 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U595 ( .A(KEYINPUT112), .B(n532), .Z(n539) );
  NOR2_X1 U596 ( .A1(n533), .A2(n539), .ZN(n534) );
  XOR2_X1 U597 ( .A(G85GAT), .B(n534), .Z(G1336GAT) );
  NOR2_X1 U598 ( .A1(n539), .A2(n535), .ZN(n537) );
  XNOR2_X1 U599 ( .A(G92GAT), .B(KEYINPUT113), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n537), .B(n536), .ZN(G1337GAT) );
  NOR2_X1 U601 ( .A1(n539), .A2(n546), .ZN(n538) );
  XOR2_X1 U602 ( .A(G99GAT), .B(n538), .Z(G1338GAT) );
  NOR2_X1 U603 ( .A1(n544), .A2(n539), .ZN(n540) );
  XOR2_X1 U604 ( .A(KEYINPUT44), .B(n540), .Z(n541) );
  XNOR2_X1 U605 ( .A(G106GAT), .B(n541), .ZN(G1339GAT) );
  AND2_X1 U606 ( .A1(n543), .A2(n542), .ZN(n556) );
  NAND2_X1 U607 ( .A1(n544), .A2(n556), .ZN(n545) );
  NOR2_X1 U608 ( .A1(n546), .A2(n545), .ZN(n553) );
  NAND2_X1 U609 ( .A1(n558), .A2(n553), .ZN(n547) );
  XNOR2_X1 U610 ( .A(n547), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U611 ( .A(G120GAT), .B(KEYINPUT49), .Z(n549) );
  NAND2_X1 U612 ( .A1(n553), .A2(n560), .ZN(n548) );
  XNOR2_X1 U613 ( .A(n549), .B(n548), .ZN(G1341GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n551) );
  INV_X1 U615 ( .A(n588), .ZN(n565) );
  NAND2_X1 U616 ( .A1(n553), .A2(n565), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U618 ( .A(G127GAT), .B(n552), .Z(G1342GAT) );
  XOR2_X1 U619 ( .A(G134GAT), .B(KEYINPUT51), .Z(n555) );
  NAND2_X1 U620 ( .A1(n553), .A2(n569), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(G1343GAT) );
  NAND2_X1 U622 ( .A1(n556), .A2(n578), .ZN(n557) );
  XNOR2_X1 U623 ( .A(KEYINPUT119), .B(n557), .ZN(n568) );
  NAND2_X1 U624 ( .A1(n558), .A2(n568), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(G141GAT), .ZN(G1344GAT) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n564) );
  XOR2_X1 U627 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n562) );
  NAND2_X1 U628 ( .A1(n568), .A2(n560), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1345GAT) );
  XOR2_X1 U631 ( .A(G155GAT), .B(KEYINPUT121), .Z(n567) );
  NAND2_X1 U632 ( .A1(n568), .A2(n565), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1346GAT) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n570), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U636 ( .A1(n580), .A2(n573), .ZN(n571) );
  XOR2_X1 U637 ( .A(G169GAT), .B(n571), .Z(G1348GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n577) );
  XOR2_X1 U639 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n575) );
  XNOR2_X1 U640 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1349GAT) );
  NAND2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n590) );
  NOR2_X1 U644 ( .A1(n590), .A2(n580), .ZN(n584) );
  XOR2_X1 U645 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n582) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(G1352GAT) );
  NOR2_X1 U649 ( .A1(n375), .A2(n590), .ZN(n586) );
  XNOR2_X1 U650 ( .A(KEYINPUT126), .B(KEYINPUT61), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(G204GAT), .B(n587), .ZN(G1353GAT) );
  NOR2_X1 U653 ( .A1(n588), .A2(n590), .ZN(n589) );
  XOR2_X1 U654 ( .A(G211GAT), .B(n589), .Z(G1354GAT) );
  NOR2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n593) );
  XNOR2_X1 U656 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U658 ( .A(G218GAT), .B(n594), .ZN(G1355GAT) );
endmodule

