//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 0 0 1 0 0 0 0 0 1 0 1 1 1 1 1 0 1 0 1 0 0 1 0 0 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n450, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n545, new_n546, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n586, new_n587, new_n588,
    new_n591, new_n593, new_n594, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1126, new_n1127, new_n1128, new_n1129;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT66), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(G125), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g040(.A(KEYINPUT68), .B(G125), .C1(new_n461), .C2(new_n462), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  OAI211_X1 g047(.A(G137), .B(new_n470), .C1(new_n461), .C2(new_n462), .ZN(new_n473));
  AND3_X1   g048(.A1(new_n469), .A2(new_n472), .A3(new_n473), .ZN(G160));
  INV_X1    g049(.A(new_n462), .ZN(new_n475));
  NAND2_X1  g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(G2105), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  XOR2_X1   g053(.A(new_n478), .B(KEYINPUT69), .Z(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(G112), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(new_n481), .B2(G2105), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT70), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n470), .B1(new_n475), .B2(new_n476), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(G124), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n479), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT71), .ZN(G162));
  OAI211_X1 g062(.A(G126), .B(G2105), .C1(new_n461), .C2(new_n462), .ZN(new_n488));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n489), .A2(new_n491), .A3(G2104), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(new_n461), .B2(new_n462), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n495), .B(new_n498), .C1(new_n462), .C2(new_n461), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n493), .B1(new_n497), .B2(new_n499), .ZN(G164));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  OR2_X1    g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G50), .ZN(new_n505));
  XNOR2_X1  g080(.A(new_n505), .B(KEYINPUT72), .ZN(new_n506));
  OR2_X1    g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n502), .A2(new_n503), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(new_n509), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n510), .A2(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n506), .A2(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  XOR2_X1   g092(.A(KEYINPUT73), .B(KEYINPUT7), .Z(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n518), .B(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n504), .A2(G51), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n523));
  INV_X1    g098(.A(G89), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n513), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n522), .A2(new_n525), .ZN(G168));
  AOI22_X1  g101(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n527), .A2(new_n511), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n504), .A2(G52), .ZN(new_n529));
  INV_X1    g104(.A(G90), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n513), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n528), .A2(new_n531), .ZN(G171));
  AND2_X1   g107(.A1(new_n509), .A2(G56), .ZN(new_n533));
  AND2_X1   g108(.A1(G68), .A2(G543), .ZN(new_n534));
  OAI21_X1  g109(.A(G651), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT74), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n512), .A2(new_n509), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n538), .A2(G81), .B1(G43), .B2(new_n504), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n535), .A2(new_n536), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  NAND4_X1  g118(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(G188));
  NAND2_X1  g122(.A1(new_n504), .A2(G53), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT9), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n538), .A2(G91), .ZN(new_n550));
  XNOR2_X1  g125(.A(KEYINPUT75), .B(G65), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n509), .A2(new_n551), .B1(G78), .B2(G543), .ZN(new_n552));
  OAI211_X1 g127(.A(new_n549), .B(new_n550), .C1(new_n511), .C2(new_n552), .ZN(G299));
  XNOR2_X1  g128(.A(G171), .B(KEYINPUT76), .ZN(G301));
  INV_X1    g129(.A(G168), .ZN(G286));
  OAI21_X1  g130(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT77), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n512), .A2(new_n509), .A3(G87), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT77), .ZN(new_n559));
  OAI211_X1 g134(.A(new_n559), .B(G651), .C1(new_n509), .C2(G74), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n504), .A2(G49), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n557), .A2(new_n558), .A3(new_n560), .A4(new_n561), .ZN(G288));
  INV_X1    g137(.A(G61), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n563), .B1(new_n507), .B2(new_n508), .ZN(new_n564));
  AND2_X1   g139(.A1(G73), .A2(G543), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n504), .A2(G48), .ZN(new_n567));
  AND2_X1   g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n538), .A2(G86), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT78), .ZN(G305));
  AOI22_X1  g146(.A1(new_n538), .A2(G85), .B1(G47), .B2(new_n504), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT79), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n511), .B2(new_n574), .ZN(G290));
  INV_X1    g150(.A(G868), .ZN(new_n576));
  NOR2_X1   g151(.A1(G301), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n504), .A2(G54), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n509), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n579));
  AND3_X1   g154(.A1(new_n538), .A2(KEYINPUT10), .A3(G92), .ZN(new_n580));
  AOI21_X1  g155(.A(KEYINPUT10), .B1(new_n538), .B2(G92), .ZN(new_n581));
  OAI221_X1 g156(.A(new_n578), .B1(new_n511), .B2(new_n579), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT80), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n577), .B1(new_n583), .B2(new_n576), .ZN(G321));
  XOR2_X1   g159(.A(G321), .B(KEYINPUT81), .Z(G284));
  INV_X1    g160(.A(KEYINPUT82), .ZN(new_n586));
  NOR2_X1   g161(.A1(G168), .A2(new_n576), .ZN(new_n587));
  AOI211_X1 g162(.A(new_n586), .B(new_n587), .C1(new_n576), .C2(G299), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(new_n586), .B2(new_n587), .ZN(G297));
  AOI21_X1  g164(.A(new_n588), .B1(new_n586), .B2(new_n587), .ZN(G280));
  INV_X1    g165(.A(G559), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n583), .B1(new_n591), .B2(G860), .ZN(G148));
  NAND2_X1  g167(.A1(new_n583), .A2(new_n591), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(G868), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(G868), .B2(new_n542), .ZN(G323));
  XNOR2_X1  g170(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g171(.A1(new_n477), .A2(G135), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n470), .A2(G111), .ZN(new_n598));
  OAI21_X1  g173(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n599));
  AND3_X1   g174(.A1(new_n484), .A2(KEYINPUT83), .A3(G123), .ZN(new_n600));
  AOI21_X1  g175(.A(KEYINPUT83), .B1(new_n484), .B2(G123), .ZN(new_n601));
  OAI221_X1 g176(.A(new_n597), .B1(new_n598), .B2(new_n599), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(G2096), .ZN(new_n603));
  INV_X1    g178(.A(G2100), .ZN(new_n604));
  XNOR2_X1  g179(.A(KEYINPUT3), .B(G2104), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(new_n471), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT12), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT13), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n603), .B1(new_n604), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n602), .A2(G2096), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n609), .B(new_n610), .C1(new_n604), .C2(new_n608), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(KEYINPUT84), .Z(G156));
  XOR2_X1   g187(.A(KEYINPUT15), .B(G2435), .Z(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(G2438), .ZN(new_n614));
  XNOR2_X1  g189(.A(G2427), .B(G2430), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT86), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n614), .A2(new_n616), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n617), .A2(KEYINPUT14), .A3(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(G1341), .B(G1348), .Z(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n619), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(G2451), .B(G2454), .Z(new_n624));
  XNOR2_X1  g199(.A(G2443), .B(G2446), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n623), .A2(new_n626), .ZN(new_n628));
  AND3_X1   g203(.A1(new_n627), .A2(G14), .A3(new_n628), .ZN(G401));
  INV_X1    g204(.A(KEYINPUT18), .ZN(new_n630));
  XOR2_X1   g205(.A(G2084), .B(G2090), .Z(new_n631));
  XNOR2_X1  g206(.A(G2067), .B(G2678), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(KEYINPUT17), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n631), .A2(new_n632), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n630), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(new_n604), .ZN(new_n637));
  XOR2_X1   g212(.A(G2072), .B(G2078), .Z(new_n638));
  AOI21_X1  g213(.A(new_n638), .B1(new_n633), .B2(KEYINPUT18), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2096), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n637), .B(new_n640), .ZN(G227));
  XOR2_X1   g216(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n642));
  XNOR2_X1  g217(.A(G1971), .B(G1976), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G1956), .B(G2474), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1961), .B(G1966), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT20), .ZN(new_n649));
  AND2_X1   g224(.A1(new_n645), .A2(new_n646), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n644), .A2(new_n650), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n647), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n649), .B(new_n651), .C1(new_n644), .C2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT88), .ZN(new_n654));
  XOR2_X1   g229(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1991), .B(G1996), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G1981), .B(G1986), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(G229));
  INV_X1    g235(.A(G16), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n542), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n662), .B1(new_n661), .B2(G19), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  AND2_X1   g239(.A1(new_n664), .A2(G1341), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(G1341), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n661), .A2(G20), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT23), .Z(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(G299), .B2(G16), .ZN(new_n669));
  INV_X1    g244(.A(G1956), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n665), .A2(new_n666), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n661), .A2(G4), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n673), .B1(new_n583), .B2(new_n661), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT90), .B(G1348), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n677));
  INV_X1    g252(.A(G29), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(G26), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n677), .B(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n477), .A2(G140), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n484), .A2(G128), .ZN(new_n682));
  OR2_X1    g257(.A1(G104), .A2(G2105), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n683), .B(G2104), .C1(G116), .C2(new_n470), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n681), .A2(new_n682), .A3(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n680), .B1(new_n686), .B2(new_n678), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT92), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G2067), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n672), .A2(new_n676), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n678), .A2(G35), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT100), .Z(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G162), .B2(new_n678), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT29), .ZN(new_n694));
  INV_X1    g269(.A(G2090), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(G27), .A2(G29), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(G164), .B2(G29), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n698), .A2(G2078), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n661), .A2(G5), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G171), .B2(new_n661), .ZN(new_n701));
  OAI22_X1  g276(.A1(new_n701), .A2(G1961), .B1(G2078), .B2(new_n698), .ZN(new_n702));
  AOI22_X1  g277(.A1(new_n477), .A2(G141), .B1(G105), .B2(new_n471), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n484), .A2(G129), .ZN(new_n704));
  NAND3_X1  g279(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT26), .Z(new_n706));
  NAND3_X1  g281(.A1(new_n703), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  MUX2_X1   g282(.A(G32), .B(new_n707), .S(G29), .Z(new_n708));
  XOR2_X1   g283(.A(KEYINPUT27), .B(G1996), .Z(new_n709));
  AOI211_X1 g284(.A(new_n699), .B(new_n702), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n661), .A2(G21), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G168), .B2(new_n661), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT96), .B(G1966), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n708), .A2(new_n709), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT31), .B(G11), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT97), .B(G28), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n717), .A2(KEYINPUT30), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(KEYINPUT30), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(new_n678), .ZN(new_n720));
  OAI221_X1 g295(.A(new_n716), .B1(new_n718), .B2(new_n720), .C1(new_n602), .C2(new_n678), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n715), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n710), .A2(new_n714), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n701), .A2(G1961), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT98), .Z(new_n725));
  XOR2_X1   g300(.A(KEYINPUT94), .B(KEYINPUT25), .Z(new_n726));
  NAND3_X1  g301(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n477), .A2(G139), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n605), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n730), .A2(new_n470), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT95), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n728), .B(new_n729), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n732), .B2(new_n731), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G29), .ZN(new_n735));
  NOR2_X1   g310(.A1(G29), .A2(G33), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT93), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G2072), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT24), .ZN(new_n741));
  INV_X1    g316(.A(G34), .ZN(new_n742));
  AOI21_X1  g317(.A(G29), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n741), .B2(new_n742), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G160), .B2(new_n678), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n745), .A2(G2084), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(G2084), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n740), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n738), .A2(new_n739), .ZN(new_n749));
  NOR4_X1   g324(.A1(new_n723), .A2(new_n725), .A3(new_n748), .A4(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n696), .B1(KEYINPUT99), .B2(new_n750), .ZN(new_n751));
  AOI211_X1 g326(.A(new_n690), .B(new_n751), .C1(KEYINPUT99), .C2(new_n750), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n678), .A2(G25), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n477), .A2(G131), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n484), .A2(G119), .ZN(new_n755));
  OR2_X1    g330(.A1(G95), .A2(G2105), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n756), .B(G2104), .C1(G107), .C2(new_n470), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n754), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n753), .B1(new_n759), .B2(new_n678), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT35), .B(G1991), .Z(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n661), .A2(G24), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G290), .B2(G16), .ZN(new_n764));
  INV_X1    g339(.A(G1986), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n762), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n765), .B2(new_n764), .ZN(new_n767));
  MUX2_X1   g342(.A(G6), .B(G305), .S(G16), .Z(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT32), .B(G1981), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT89), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n768), .A2(new_n770), .ZN(new_n772));
  MUX2_X1   g347(.A(G23), .B(G288), .S(G16), .Z(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT33), .B(G1976), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n661), .A2(G22), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G166), .B2(new_n661), .ZN(new_n777));
  INV_X1    g352(.A(G1971), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n771), .A2(new_n772), .A3(new_n775), .A4(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n767), .B1(new_n780), .B2(KEYINPUT34), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(KEYINPUT34), .B2(new_n780), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT36), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n752), .A2(new_n783), .ZN(G150));
  INV_X1    g359(.A(G150), .ZN(G311));
  AOI22_X1  g360(.A1(new_n538), .A2(G93), .B1(G55), .B2(new_n504), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT101), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n509), .A2(G67), .ZN(new_n788));
  NAND2_X1  g363(.A1(G80), .A2(G543), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n511), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n786), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n790), .A2(new_n787), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n793), .A2(G860), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT37), .Z(new_n795));
  AOI21_X1  g370(.A(new_n793), .B1(KEYINPUT102), .B2(new_n542), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(KEYINPUT102), .B2(new_n542), .ZN(new_n797));
  INV_X1    g372(.A(new_n793), .ZN(new_n798));
  OR3_X1    g373(.A1(new_n798), .A2(KEYINPUT102), .A3(new_n542), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT38), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n583), .A2(G559), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n802), .B(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT39), .ZN(new_n806));
  AOI21_X1  g381(.A(G860), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n802), .B(new_n803), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(KEYINPUT39), .ZN(new_n809));
  AND3_X1   g384(.A1(new_n807), .A2(KEYINPUT103), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(KEYINPUT103), .B1(new_n807), .B2(new_n809), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n795), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(KEYINPUT104), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT104), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n814), .B(new_n795), .C1(new_n810), .C2(new_n811), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(new_n815), .ZN(G145));
  XNOR2_X1  g391(.A(new_n734), .B(new_n707), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n758), .B(KEYINPUT105), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(new_n607), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n817), .B(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(G164), .B(new_n685), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n484), .A2(G130), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n470), .A2(G118), .ZN(new_n823));
  OAI21_X1  g398(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(G142), .B2(new_n477), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n821), .B(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n820), .B(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(G160), .B(new_n602), .ZN(new_n830));
  XNOR2_X1  g405(.A(G162), .B(new_n830), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT107), .Z(new_n832));
  NAND2_X1  g407(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n833), .A2(KEYINPUT108), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(KEYINPUT108), .ZN(new_n835));
  AOI21_X1  g410(.A(G37), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n828), .A2(new_n831), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT106), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n836), .A2(KEYINPUT40), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(KEYINPUT40), .B1(new_n836), .B2(new_n838), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n839), .A2(new_n840), .ZN(G395));
  XNOR2_X1  g416(.A(new_n800), .B(new_n593), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n582), .B(G299), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT41), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(new_n843), .B2(new_n842), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT42), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n847), .ZN(new_n849));
  XNOR2_X1  g424(.A(G290), .B(G305), .ZN(new_n850));
  XNOR2_X1  g425(.A(G303), .B(G288), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n853), .A2(KEYINPUT109), .ZN(new_n854));
  AND3_X1   g429(.A1(new_n848), .A2(new_n849), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n854), .B1(new_n848), .B2(new_n849), .ZN(new_n856));
  OAI21_X1  g431(.A(G868), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(G868), .B2(new_n798), .ZN(G295));
  OAI21_X1  g433(.A(new_n857), .B1(G868), .B2(new_n798), .ZN(G331));
  NOR2_X1   g434(.A1(G168), .A2(G171), .ZN(new_n860));
  INV_X1    g435(.A(G301), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n860), .B1(new_n861), .B2(G168), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n800), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n862), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n797), .A2(new_n799), .A3(new_n864), .ZN(new_n865));
  AND3_X1   g440(.A1(new_n863), .A2(new_n865), .A3(new_n844), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n843), .B1(new_n863), .B2(new_n865), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n853), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(G37), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n866), .ZN(new_n871));
  INV_X1    g446(.A(new_n867), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n871), .A2(new_n852), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT110), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT110), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n871), .A2(new_n872), .A3(new_n875), .A4(new_n852), .ZN(new_n876));
  AOI211_X1 g451(.A(KEYINPUT43), .B(new_n870), .C1(new_n874), .C2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT111), .ZN(new_n878));
  OAI21_X1  g453(.A(KEYINPUT44), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n870), .B1(new_n874), .B2(new_n876), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT43), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n879), .B1(new_n882), .B2(new_n877), .ZN(new_n883));
  INV_X1    g458(.A(new_n882), .ZN(new_n884));
  INV_X1    g459(.A(new_n877), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n884), .A2(new_n885), .A3(new_n878), .A4(KEYINPUT44), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n883), .A2(new_n886), .ZN(G397));
  AOI22_X1  g462(.A1(new_n463), .A2(new_n464), .B1(G113), .B2(G2104), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n470), .B1(new_n888), .B2(new_n466), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n473), .A2(new_n472), .A3(G40), .ZN(new_n890));
  OAI21_X1  g465(.A(KEYINPUT112), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT112), .ZN(new_n892));
  INV_X1    g467(.A(new_n890), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n469), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT45), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n896), .B1(G164), .B2(G1384), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  OR3_X1    g474(.A1(new_n899), .A2(G1986), .A3(G290), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(G1996), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n707), .B(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(G2067), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n685), .B(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n759), .A2(new_n761), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n759), .A2(new_n761), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n903), .A2(new_n905), .A3(new_n906), .A4(new_n907), .ZN(new_n908));
  AOI22_X1  g483(.A1(new_n901), .A2(KEYINPUT48), .B1(new_n898), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(KEYINPUT48), .B2(new_n901), .ZN(new_n910));
  INV_X1    g485(.A(new_n905), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n898), .B1(new_n707), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n898), .A2(new_n902), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n913), .A2(KEYINPUT46), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(KEYINPUT46), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n912), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT47), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n903), .A2(new_n905), .ZN(new_n918));
  OAI22_X1  g493(.A1(new_n918), .A2(new_n906), .B1(G2067), .B2(new_n685), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(new_n898), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n910), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT127), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n896), .A2(G1384), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT113), .B1(G164), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n499), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n498), .B1(new_n605), .B2(new_n495), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n488), .B(new_n492), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT113), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n928), .A2(new_n929), .A3(new_n923), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n897), .A2(new_n925), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n892), .B1(new_n469), .B2(new_n893), .ZN(new_n932));
  AOI211_X1 g507(.A(KEYINPUT112), .B(new_n890), .C1(new_n468), .C2(G2105), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(G1971), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT50), .ZN(new_n937));
  INV_X1    g512(.A(G1384), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n926), .A2(new_n927), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n937), .B(new_n938), .C1(new_n939), .C2(new_n493), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n891), .A2(new_n936), .A3(new_n894), .A4(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n941), .A2(G2090), .ZN(new_n942));
  OAI21_X1  g517(.A(G8), .B1(new_n935), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(G303), .A2(G8), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT55), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n943), .A2(new_n949), .A3(KEYINPUT116), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT116), .ZN(new_n951));
  INV_X1    g526(.A(G8), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n934), .A2(new_n695), .A3(new_n936), .A4(new_n940), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n897), .A2(new_n925), .A3(new_n930), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n778), .B1(new_n954), .B2(new_n895), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n952), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n951), .B1(new_n956), .B2(new_n948), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n950), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT125), .ZN(new_n959));
  NOR2_X1   g534(.A1(G164), .A2(G1384), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n891), .A2(new_n894), .A3(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(G1976), .ZN(new_n962));
  OR2_X1    g537(.A1(G288), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n961), .A2(G8), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT52), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT52), .B1(G288), .B2(new_n962), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n961), .A2(G8), .A3(new_n963), .A4(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT49), .ZN(new_n968));
  INV_X1    g543(.A(G1981), .ZN(new_n969));
  AND4_X1   g544(.A1(new_n969), .A2(new_n569), .A3(new_n566), .A4(new_n567), .ZN(new_n970));
  XOR2_X1   g545(.A(KEYINPUT115), .B(G86), .Z(new_n971));
  NAND3_X1  g546(.A1(new_n971), .A2(new_n512), .A3(new_n509), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n566), .A2(new_n567), .A3(new_n972), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n973), .A2(G1981), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n968), .B1(new_n970), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n568), .A2(new_n969), .A3(new_n569), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n973), .A2(G1981), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n976), .A2(KEYINPUT49), .A3(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n975), .A2(new_n961), .A3(new_n978), .A4(G8), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n965), .A2(new_n967), .A3(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n936), .A2(KEYINPUT114), .A3(new_n940), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n928), .A2(new_n938), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT114), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n982), .A2(new_n983), .A3(KEYINPUT50), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n985), .A2(new_n695), .A3(new_n934), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n952), .B1(new_n986), .B2(new_n955), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n980), .B1(new_n948), .B2(new_n987), .ZN(new_n988));
  AND3_X1   g563(.A1(new_n958), .A2(new_n959), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n959), .B1(new_n958), .B2(new_n988), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT62), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT51), .ZN(new_n993));
  XOR2_X1   g568(.A(KEYINPUT117), .B(G2084), .Z(new_n994));
  AND3_X1   g569(.A1(new_n891), .A2(new_n894), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n928), .A2(new_n923), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n891), .A2(new_n897), .A3(new_n894), .A4(new_n996), .ZN(new_n997));
  AOI22_X1  g572(.A1(new_n985), .A2(new_n995), .B1(new_n997), .B2(new_n713), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n952), .B1(new_n998), .B2(G168), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n891), .A2(new_n894), .A3(new_n994), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n1000), .B1(new_n984), .B2(new_n981), .ZN(new_n1001));
  INV_X1    g576(.A(new_n713), .ZN(new_n1002));
  AOI22_X1  g577(.A1(new_n982), .A2(new_n896), .B1(new_n928), .B2(new_n923), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1002), .B1(new_n934), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(G286), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n993), .B1(new_n999), .B2(new_n1005), .ZN(new_n1006));
  AOI211_X1 g581(.A(KEYINPUT51), .B(new_n952), .C1(new_n998), .C2(G168), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n1006), .A2(KEYINPUT123), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT123), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n985), .A2(new_n995), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n997), .A2(new_n713), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(G168), .A3(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1005), .A2(G8), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT51), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n999), .A2(new_n993), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1009), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n992), .B1(new_n1008), .B2(new_n1016), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n954), .A2(new_n895), .A3(G2078), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n895), .B1(new_n981), .B2(new_n984), .ZN(new_n1019));
  OAI22_X1  g594(.A1(new_n1018), .A2(KEYINPUT53), .B1(new_n1019), .B2(G1961), .ZN(new_n1020));
  INV_X1    g595(.A(G2078), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT53), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n997), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n861), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT123), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1014), .A2(new_n1009), .A3(new_n1015), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1026), .A2(new_n1027), .A3(KEYINPUT62), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n991), .A2(new_n1017), .A3(new_n1025), .A4(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT63), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT116), .B1(new_n943), .B2(new_n949), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n956), .A2(new_n951), .A3(new_n948), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n988), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI211_X1 g608(.A(G8), .B(G168), .C1(new_n1001), .C2(new_n1004), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1030), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT118), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1037), .B(new_n1030), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1034), .A2(new_n1030), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n988), .B(new_n1039), .C1(new_n948), .C2(new_n987), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1036), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(G288), .A2(G1976), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n970), .B1(new_n979), .B2(new_n1042), .ZN(new_n1043));
  AOI211_X1 g618(.A(new_n952), .B(new_n1043), .C1(new_n960), .C2(new_n934), .ZN(new_n1044));
  INV_X1    g619(.A(new_n987), .ZN(new_n1045));
  NOR3_X1   g620(.A1(new_n1045), .A2(new_n949), .A3(new_n980), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  AND3_X1   g622(.A1(new_n1029), .A2(new_n1041), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1033), .A2(KEYINPUT125), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n958), .A2(new_n959), .A3(new_n988), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n985), .A2(new_n934), .ZN(new_n1051));
  INV_X1    g626(.A(G1961), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n931), .A2(new_n1021), .A3(new_n934), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n469), .A2(new_n893), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n954), .A2(new_n1057), .A3(new_n1022), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1053), .A2(new_n1056), .A3(G301), .A4(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1024), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT124), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT124), .ZN(new_n1064));
  AOI211_X1 g639(.A(new_n1064), .B(KEYINPUT54), .C1(new_n1024), .C2(new_n1060), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1049), .B(new_n1050), .C1(new_n1063), .C2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1020), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1023), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1067), .A2(G301), .A3(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(G171), .B1(new_n1020), .B2(new_n1058), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(new_n1070), .A3(KEYINPUT54), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1026), .A2(new_n1027), .A3(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT126), .B1(new_n1066), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT54), .B1(new_n1024), .B2(new_n1060), .ZN(new_n1074));
  XNOR2_X1  g649(.A(new_n1074), .B(KEYINPUT124), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1026), .A2(new_n1027), .A3(new_n1071), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT126), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1075), .A2(new_n991), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n542), .A2(KEYINPUT122), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n954), .A2(new_n895), .ZN(new_n1080));
  XOR2_X1   g655(.A(KEYINPUT58), .B(G1341), .Z(new_n1081));
  AOI22_X1  g656(.A1(new_n1080), .A2(new_n902), .B1(new_n961), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT121), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT121), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n954), .A2(new_n895), .A3(G1996), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n961), .A2(new_n1081), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1084), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1079), .B1(new_n1083), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n961), .A2(G2067), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n1051), .B2(new_n675), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n1092), .B(new_n582), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1089), .A2(new_n1090), .B1(new_n1093), .B2(KEYINPUT60), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n582), .A2(KEYINPUT60), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n1088), .A2(KEYINPUT59), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT56), .B(G2072), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1080), .A2(new_n1097), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n941), .A2(KEYINPUT119), .A3(new_n670), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT119), .B1(new_n941), .B2(new_n670), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  XOR2_X1   g676(.A(G299), .B(KEYINPUT57), .Z(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1102), .B(new_n1098), .C1(new_n1100), .C2(new_n1099), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT61), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1104), .A2(KEYINPUT61), .A3(new_n1105), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1094), .A2(new_n1096), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1092), .A2(new_n582), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n1105), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n1104), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1113), .B(KEYINPUT120), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1110), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1073), .A2(new_n1078), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1048), .A2(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g692(.A(G290), .B(new_n765), .ZN(new_n1118));
  INV_X1    g693(.A(new_n908), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n899), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n922), .B1(new_n1117), .B2(new_n1121), .ZN(new_n1122));
  AOI211_X1 g697(.A(KEYINPUT127), .B(new_n1120), .C1(new_n1048), .C2(new_n1116), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n921), .B1(new_n1122), .B2(new_n1123), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n1126));
  NAND2_X1  g700(.A1(new_n836), .A2(new_n838), .ZN(new_n1127));
  OR2_X1    g701(.A1(G227), .A2(new_n459), .ZN(new_n1128));
  NOR3_X1   g702(.A1(G229), .A2(G401), .A3(new_n1128), .ZN(new_n1129));
  AND3_X1   g703(.A1(new_n1126), .A2(new_n1127), .A3(new_n1129), .ZN(G308));
  NAND3_X1  g704(.A1(new_n1126), .A2(new_n1127), .A3(new_n1129), .ZN(G225));
endmodule


