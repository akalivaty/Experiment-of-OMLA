//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0 1 1 1 1 0 0 0 0 1 1 0 0 0 0 0 0 0 0 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n456, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n544, new_n545, new_n546, new_n547, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n558, new_n559,
    new_n560, new_n561, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n629, new_n630, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1230, new_n1231, new_n1232,
    new_n1233;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT65), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  AOI22_X1  g029(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n452), .ZN(G319));
  INV_X1    g030(.A(G2105), .ZN(new_n456));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n457));
  AND2_X1   g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n463), .A2(KEYINPUT66), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n460), .A2(new_n465), .A3(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n456), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n462), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n463), .A2(new_n464), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(new_n456), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n468), .A2(new_n474), .ZN(G160));
  NOR2_X1   g050(.A1(new_n458), .A2(new_n459), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n476), .A2(new_n456), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n456), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  INV_X1    g059(.A(G138), .ZN(new_n485));
  NOR3_X1   g060(.A1(new_n485), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n460), .A2(new_n465), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n460), .A2(new_n465), .A3(KEYINPUT69), .A4(new_n486), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n471), .A2(G138), .A3(new_n456), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n489), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n471), .A2(G126), .A3(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  AND2_X1   g070(.A1(KEYINPUT67), .A2(G114), .ZN(new_n496));
  NOR2_X1   g071(.A1(KEYINPUT67), .A2(G114), .ZN(new_n497));
  OAI21_X1  g072(.A(G2105), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT68), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT68), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n500), .B(G2105), .C1(new_n496), .C2(new_n497), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n495), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n493), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT70), .B1(new_n508), .B2(G651), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT6), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n509), .A2(new_n512), .B1(new_n508), .B2(G651), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(G50), .A3(G543), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n513), .A2(G88), .A3(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n519), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n521));
  OAI211_X1 g096(.A(new_n514), .B(new_n520), .C1(new_n511), .C2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT71), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n521), .A2(new_n511), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT71), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n524), .A2(new_n525), .A3(new_n514), .A4(new_n520), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n523), .A2(new_n526), .ZN(G166));
  NAND2_X1  g102(.A1(new_n513), .A2(G543), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G51), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n509), .A2(new_n512), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n508), .A2(G651), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n531), .A2(new_n532), .A3(new_n519), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  XNOR2_X1  g109(.A(KEYINPUT72), .B(G89), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n539));
  AND2_X1   g114(.A1(G63), .A2(G651), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n538), .A2(new_n539), .B1(new_n519), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n530), .A2(new_n536), .A3(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  NAND2_X1  g118(.A1(new_n529), .A2(G52), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n534), .A2(G90), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n511), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  AOI22_X1  g124(.A1(new_n519), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(new_n511), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n513), .A2(G81), .A3(new_n519), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n513), .A2(G43), .A3(G543), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT74), .ZN(new_n559));
  XOR2_X1   g134(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n560));
  XNOR2_X1  g135(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  INV_X1    g137(.A(KEYINPUT76), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n513), .A2(new_n563), .A3(G91), .A4(new_n519), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n531), .A2(G91), .A3(new_n532), .A4(new_n519), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(KEYINPUT76), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT77), .ZN(new_n567));
  AND2_X1   g142(.A1(KEYINPUT5), .A2(G543), .ZN(new_n568));
  NOR2_X1   g143(.A1(KEYINPUT5), .A2(G543), .ZN(new_n569));
  OAI21_X1  g144(.A(G65), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n567), .B1(new_n572), .B2(G651), .ZN(new_n573));
  AOI211_X1 g148(.A(KEYINPUT77), .B(new_n511), .C1(new_n570), .C2(new_n571), .ZN(new_n574));
  OAI211_X1 g149(.A(new_n564), .B(new_n566), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n531), .A2(G53), .A3(G543), .A4(new_n532), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT75), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n577), .A2(KEYINPUT9), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g154(.A(KEYINPUT75), .B(KEYINPUT9), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n513), .A2(G53), .A3(G543), .A4(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n575), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G299));
  INV_X1    g159(.A(G166), .ZN(G303));
  NAND3_X1  g160(.A1(new_n513), .A2(G49), .A3(G543), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n587));
  INV_X1    g162(.A(G87), .ZN(new_n588));
  OAI211_X1 g163(.A(new_n586), .B(new_n587), .C1(new_n533), .C2(new_n588), .ZN(G288));
  NAND3_X1  g164(.A1(new_n513), .A2(G86), .A3(new_n519), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n531), .A2(G48), .A3(G543), .A4(new_n532), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n517), .B2(new_n518), .ZN(new_n593));
  AND2_X1   g168(.A1(G73), .A2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n590), .A2(new_n591), .A3(new_n595), .ZN(G305));
  NAND2_X1  g171(.A1(new_n534), .A2(G85), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n598), .A2(new_n511), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n513), .A2(G47), .A3(G543), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n597), .A2(new_n599), .A3(new_n600), .ZN(G290));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NOR2_X1   g177(.A1(G301), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(G92), .ZN(new_n604));
  OR3_X1    g179(.A1(new_n533), .A2(KEYINPUT78), .A3(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(KEYINPUT78), .B1(new_n533), .B2(new_n604), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n605), .A2(KEYINPUT10), .A3(new_n606), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n519), .A2(G66), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT80), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n511), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n528), .A2(KEYINPUT79), .ZN(new_n615));
  INV_X1    g190(.A(G54), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(new_n528), .B2(KEYINPUT79), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n614), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n609), .A2(new_n610), .A3(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  OR2_X1    g195(.A1(new_n620), .A2(KEYINPUT81), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(KEYINPUT81), .ZN(new_n622));
  AND2_X1   g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n603), .B1(new_n623), .B2(new_n602), .ZN(G284));
  AOI21_X1  g199(.A(new_n603), .B1(new_n623), .B2(new_n602), .ZN(G321));
  NAND2_X1  g200(.A1(G286), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(new_n583), .B2(G868), .ZN(G297));
  OAI21_X1  g202(.A(new_n626), .B1(new_n583), .B2(G868), .ZN(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n623), .B1(new_n629), .B2(G860), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT82), .ZN(G148));
  NAND3_X1  g206(.A1(new_n621), .A2(new_n629), .A3(new_n622), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G868), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g210(.A1(new_n460), .A2(new_n465), .ZN(new_n636));
  NOR3_X1   g211(.A1(new_n636), .A2(new_n462), .A3(G2105), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT12), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT13), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n643), .A2(G2100), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT83), .Z(new_n645));
  NAND2_X1  g220(.A1(new_n477), .A2(G135), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n479), .A2(G123), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n456), .A2(G111), .ZN(new_n648));
  OAI21_X1  g223(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n649));
  OAI211_X1 g224(.A(new_n646), .B(new_n647), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2096), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(new_n643), .B2(G2100), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n645), .A2(new_n652), .ZN(G156));
  INV_X1    g228(.A(KEYINPUT14), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2427), .B(G2438), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2430), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT15), .B(G2435), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n654), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n658), .B1(new_n657), .B2(new_n656), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2451), .B(G2454), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1341), .B(G1348), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n659), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2443), .B(G2446), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(G14), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n664), .A2(new_n665), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(G401));
  XOR2_X1   g244(.A(G2072), .B(G2078), .Z(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT17), .Z(new_n671));
  XNOR2_X1  g246(.A(G2067), .B(G2678), .ZN(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n671), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT84), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n671), .A2(new_n672), .ZN(new_n677));
  INV_X1    g252(.A(new_n670), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n677), .B(new_n674), .C1(new_n678), .C2(new_n672), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n678), .A2(new_n672), .A3(new_n673), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT18), .Z(new_n681));
  NAND3_X1  g256(.A1(new_n676), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G2096), .B(G2100), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(G227));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1956), .B(G2474), .Z(new_n688));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n690), .A2(KEYINPUT85), .ZN(new_n691));
  XOR2_X1   g266(.A(G1971), .B(G1976), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT19), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(KEYINPUT85), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n691), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT20), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT86), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n688), .A2(new_n689), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(new_n690), .ZN(new_n699));
  MUX2_X1   g274(.A(new_n699), .B(new_n698), .S(new_n693), .Z(new_n700));
  NAND3_X1  g275(.A1(new_n696), .A2(new_n697), .A3(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n697), .B1(new_n696), .B2(new_n700), .ZN(new_n703));
  OAI21_X1  g278(.A(G1981), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n703), .ZN(new_n705));
  INV_X1    g280(.A(G1981), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n705), .A2(new_n706), .A3(new_n701), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n704), .A2(new_n707), .A3(G1986), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(G1986), .B1(new_n704), .B2(new_n707), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT87), .ZN(new_n712));
  NOR3_X1   g287(.A1(new_n709), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n712), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n704), .A2(new_n707), .ZN(new_n715));
  INV_X1    g290(.A(G1986), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n714), .B1(new_n717), .B2(new_n708), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n687), .B1(new_n713), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n712), .B1(new_n709), .B2(new_n710), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n717), .A2(new_n714), .A3(new_n708), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n720), .A2(new_n686), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n719), .A2(new_n722), .ZN(G229));
  NAND2_X1  g298(.A1(G303), .A2(G16), .ZN(new_n724));
  INV_X1    g299(.A(G22), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(G16), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G1971), .ZN(new_n727));
  INV_X1    g302(.A(G1971), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n724), .B(new_n728), .C1(G16), .C2(new_n725), .ZN(new_n729));
  INV_X1    g304(.A(G16), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G23), .ZN(new_n731));
  INV_X1    g306(.A(G288), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(new_n730), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT33), .B(G1976), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n727), .A2(new_n729), .A3(new_n735), .ZN(new_n736));
  MUX2_X1   g311(.A(G6), .B(G305), .S(G16), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT32), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G1981), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT90), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT34), .ZN(new_n743));
  NOR3_X1   g318(.A1(new_n736), .A2(new_n739), .A3(KEYINPUT90), .ZN(new_n744));
  OR3_X1    g319(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n743), .B1(new_n742), .B2(new_n744), .ZN(new_n746));
  NOR2_X1   g321(.A1(G16), .A2(G24), .ZN(new_n747));
  INV_X1    g322(.A(G290), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(G16), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT88), .B(G1986), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n751), .A2(KEYINPUT89), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n751), .A2(KEYINPUT89), .ZN(new_n753));
  INV_X1    g328(.A(G29), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G25), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n477), .A2(G131), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n479), .A2(G119), .ZN(new_n757));
  OR2_X1    g332(.A1(G95), .A2(G2105), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n758), .B(G2104), .C1(G107), .C2(new_n456), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n756), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n755), .B1(new_n761), .B2(new_n754), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT35), .B(G1991), .Z(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n762), .B(new_n764), .ZN(new_n765));
  NOR4_X1   g340(.A1(new_n752), .A2(new_n753), .A3(KEYINPUT91), .A4(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n745), .A2(new_n746), .A3(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT36), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n745), .A2(new_n746), .A3(KEYINPUT36), .A4(new_n766), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n456), .A2(G103), .A3(G2104), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT25), .Z(new_n772));
  INV_X1    g347(.A(G139), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n472), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT94), .ZN(new_n775));
  NAND2_X1  g350(.A1(G115), .A2(G2104), .ZN(new_n776));
  INV_X1    g351(.A(G127), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n636), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(G2105), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n780), .A2(new_n754), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n754), .B2(G33), .ZN(new_n782));
  INV_X1    g357(.A(G2072), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n477), .A2(G141), .B1(G105), .B2(new_n469), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n479), .A2(G129), .ZN(new_n786));
  NAND3_X1  g361(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT26), .Z(new_n788));
  NAND3_X1  g363(.A1(new_n785), .A2(new_n786), .A3(new_n788), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n789), .A2(KEYINPUT96), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(KEYINPUT96), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n793), .A2(new_n754), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n754), .B2(G32), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT27), .B(G1996), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT24), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(G34), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n754), .B1(new_n798), .B2(G34), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT95), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n801), .B2(new_n800), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G160), .B2(G29), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(G2084), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n754), .A2(G35), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G162), .B2(new_n754), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT29), .Z(new_n808));
  INV_X1    g383(.A(G2090), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n784), .A2(new_n797), .A3(new_n805), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n754), .A2(G27), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G164), .B2(new_n754), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G2078), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n555), .A2(G16), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G16), .B2(G19), .ZN(new_n816));
  INV_X1    g391(.A(G1341), .ZN(new_n817));
  OAI22_X1  g392(.A1(new_n816), .A2(new_n817), .B1(new_n804), .B2(G2084), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(new_n817), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(new_n795), .B2(new_n796), .ZN(new_n820));
  NOR4_X1   g395(.A1(new_n811), .A2(new_n814), .A3(new_n818), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n730), .A2(G4), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n623), .B2(new_n730), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT92), .B(G1348), .Z(new_n824));
  XOR2_X1   g399(.A(new_n823), .B(new_n824), .Z(new_n825));
  NAND2_X1  g400(.A1(new_n730), .A2(G20), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT23), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(new_n583), .B2(new_n730), .ZN(new_n828));
  INV_X1    g403(.A(G1956), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n808), .A2(new_n809), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT98), .ZN(new_n832));
  INV_X1    g407(.A(G1966), .ZN(new_n833));
  OAI21_X1  g408(.A(KEYINPUT97), .B1(G16), .B2(G21), .ZN(new_n834));
  NOR2_X1   g409(.A1(G286), .A2(new_n730), .ZN(new_n835));
  MUX2_X1   g410(.A(new_n834), .B(KEYINPUT97), .S(new_n835), .Z(new_n836));
  AOI22_X1  g411(.A1(new_n831), .A2(new_n832), .B1(new_n833), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n754), .A2(G26), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT28), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n477), .A2(G140), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n479), .A2(G128), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n456), .A2(G116), .ZN(new_n842));
  OAI21_X1  g417(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n840), .B(new_n841), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT93), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n839), .B1(new_n845), .B2(G29), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(G2067), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n837), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n730), .A2(G5), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(G171), .B2(new_n730), .ZN(new_n850));
  INV_X1    g425(.A(G1961), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  XOR2_X1   g427(.A(KEYINPUT31), .B(G11), .Z(new_n853));
  NOR2_X1   g428(.A1(new_n650), .A2(new_n754), .ZN(new_n854));
  INV_X1    g429(.A(G28), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n855), .A2(KEYINPUT30), .ZN(new_n856));
  AOI21_X1  g431(.A(G29), .B1(new_n855), .B2(KEYINPUT30), .ZN(new_n857));
  AOI211_X1 g432(.A(new_n853), .B(new_n854), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n852), .B(new_n858), .C1(new_n782), .C2(new_n783), .ZN(new_n859));
  OAI22_X1  g434(.A1(new_n831), .A2(new_n832), .B1(new_n833), .B2(new_n836), .ZN(new_n860));
  NOR3_X1   g435(.A1(new_n848), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  AND4_X1   g436(.A1(new_n821), .A2(new_n825), .A3(new_n830), .A4(new_n861), .ZN(new_n862));
  AND3_X1   g437(.A1(new_n769), .A2(new_n770), .A3(new_n862), .ZN(G311));
  NAND3_X1  g438(.A1(new_n769), .A2(new_n770), .A3(new_n862), .ZN(G150));
  NAND2_X1  g439(.A1(new_n623), .A2(G559), .ZN(new_n865));
  XOR2_X1   g440(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n866), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n623), .A2(G559), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  AOI22_X1  g445(.A1(new_n519), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n871), .A2(new_n511), .ZN(new_n872));
  XNOR2_X1  g447(.A(KEYINPUT100), .B(G55), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n513), .A2(G543), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n513), .A2(G93), .A3(new_n519), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n872), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n554), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n554), .A2(new_n876), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n870), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n867), .A2(new_n879), .A3(new_n869), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT39), .ZN(new_n884));
  AOI21_X1  g459(.A(G860), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(new_n884), .B2(new_n883), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n876), .A2(G860), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n887), .B(KEYINPUT37), .Z(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(G145));
  NAND3_X1  g464(.A1(new_n790), .A2(G164), .A3(new_n791), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(G164), .B1(new_n790), .B2(new_n791), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n780), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n792), .A2(new_n506), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n775), .A2(new_n779), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n894), .A2(new_n895), .A3(new_n890), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(new_n845), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n477), .A2(G142), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n479), .A2(G130), .ZN(new_n900));
  OR2_X1    g475(.A1(G106), .A2(G2105), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n901), .B(G2104), .C1(G118), .C2(new_n456), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n639), .A2(new_n640), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n903), .B1(new_n639), .B2(new_n640), .ZN(new_n905));
  OR3_X1    g480(.A1(new_n904), .A2(new_n905), .A3(new_n760), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n760), .B1(new_n904), .B2(new_n905), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n845), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n893), .A2(new_n910), .A3(new_n896), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n898), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n912), .A2(KEYINPUT102), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n898), .A2(new_n911), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT101), .B1(new_n914), .B2(new_n908), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT101), .ZN(new_n916));
  AOI211_X1 g491(.A(new_n916), .B(new_n909), .C1(new_n898), .C2(new_n911), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n913), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(G160), .B(new_n650), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(G162), .ZN(new_n920));
  AOI21_X1  g495(.A(G37), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n920), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n913), .B(new_n922), .C1(new_n915), .C2(new_n917), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n921), .A2(KEYINPUT40), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT40), .B1(new_n921), .B2(new_n923), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(G395));
  XNOR2_X1  g501(.A(new_n632), .B(new_n879), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n619), .A2(new_n583), .ZN(new_n928));
  NAND4_X1  g503(.A1(G299), .A2(new_n610), .A3(new_n609), .A4(new_n618), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OR2_X1    g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(new_n929), .A3(KEYINPUT41), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT41), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n927), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n590), .A2(new_n591), .A3(new_n595), .ZN(new_n936));
  XNOR2_X1  g511(.A(G290), .B(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n523), .A2(new_n526), .A3(G288), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(G288), .B1(new_n523), .B2(new_n526), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(G290), .B(G305), .ZN(new_n942));
  INV_X1    g517(.A(new_n940), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n942), .A2(new_n943), .A3(new_n938), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT103), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n941), .A2(new_n944), .A3(KEYINPUT103), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT42), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT42), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n945), .A2(new_n951), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n931), .A2(new_n935), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n953), .B1(new_n931), .B2(new_n935), .ZN(new_n955));
  OAI21_X1  g530(.A(G868), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n872), .A2(new_n874), .A3(new_n875), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n956), .B1(G868), .B2(new_n957), .ZN(G295));
  OAI21_X1  g533(.A(new_n956), .B1(G868), .B2(new_n957), .ZN(G331));
  XOR2_X1   g534(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT106), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n941), .A2(new_n944), .A3(KEYINPUT103), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT103), .B1(new_n941), .B2(new_n944), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n947), .A2(KEYINPUT106), .A3(new_n948), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(G171), .B1(new_n877), .B2(new_n878), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n555), .A2(new_n957), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n554), .A2(new_n876), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n969), .A2(G301), .A3(new_n970), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n968), .A2(new_n971), .A3(G168), .ZN(new_n972));
  AOI21_X1  g547(.A(G168), .B1(new_n968), .B2(new_n971), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n930), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n877), .A2(new_n878), .A3(G171), .ZN(new_n977));
  AOI21_X1  g552(.A(G301), .B1(new_n969), .B2(new_n970), .ZN(new_n978));
  OAI21_X1  g553(.A(G286), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n968), .A2(new_n971), .A3(G168), .ZN(new_n980));
  AOI22_X1  g555(.A1(new_n979), .A2(new_n980), .B1(new_n928), .B2(new_n929), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n934), .A2(new_n932), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n972), .A2(new_n973), .ZN(new_n983));
  AOI22_X1  g558(.A1(KEYINPUT105), .A2(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n967), .B1(new_n976), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n982), .A2(new_n983), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n930), .B(KEYINPUT105), .C1(new_n972), .C2(new_n973), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n986), .A2(new_n976), .A3(new_n949), .A4(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G37), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n961), .B1(new_n985), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n986), .A2(new_n974), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n993), .A2(new_n966), .A3(new_n965), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n994), .A2(new_n989), .A3(new_n988), .A4(new_n960), .ZN(new_n995));
  AND3_X1   g570(.A1(new_n991), .A2(new_n992), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n967), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT107), .B1(new_n990), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT107), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n994), .A2(new_n1000), .A3(new_n989), .A4(new_n988), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n999), .A2(KEYINPUT43), .A3(new_n1001), .ZN(new_n1002));
  OR3_X1    g577(.A1(new_n985), .A2(new_n990), .A3(new_n961), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n996), .B1(new_n1004), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g580(.A(G1384), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n506), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n1008));
  INV_X1    g583(.A(G40), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n468), .A2(new_n1009), .A3(new_n474), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1007), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  NOR3_X1   g586(.A1(new_n1011), .A2(new_n792), .A3(G1996), .ZN(new_n1012));
  OR2_X1    g587(.A1(new_n1012), .A2(KEYINPUT108), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(KEYINPUT108), .ZN(new_n1014));
  INV_X1    g589(.A(G2067), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n845), .B(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G1996), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1016), .B1(new_n1017), .B2(new_n793), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1011), .ZN(new_n1019));
  AOI22_X1  g594(.A1(new_n1013), .A2(new_n1014), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n761), .A2(new_n763), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n760), .A2(new_n764), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1019), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g599(.A(G290), .B(G1986), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1024), .B1(new_n1019), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT63), .ZN(new_n1027));
  AOI21_X1  g602(.A(G1384), .B1(new_n493), .B2(new_n505), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1010), .B1(new_n1028), .B2(KEYINPUT45), .ZN(new_n1029));
  AOI211_X1 g604(.A(new_n1008), .B(G1384), .C1(new_n493), .C2(new_n505), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n728), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT109), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1007), .A2(KEYINPUT50), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1028), .A2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1033), .A2(new_n809), .A3(new_n1010), .A4(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT110), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT109), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1039), .B(new_n728), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1010), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1041), .B1(new_n1007), .B2(KEYINPUT50), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1042), .A2(KEYINPUT110), .A3(new_n809), .A4(new_n1035), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1032), .A2(new_n1038), .A3(new_n1040), .A4(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(G8), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n523), .A2(new_n526), .A3(G8), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1046), .B(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1045), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n506), .A2(new_n1010), .A3(new_n1006), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n732), .A2(G1976), .ZN(new_n1052));
  XOR2_X1   g627(.A(KEYINPUT111), .B(G1976), .Z(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT52), .B1(G288), .B2(new_n1053), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1051), .A2(G8), .A3(new_n1052), .A4(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT112), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G8), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1058), .B1(new_n1028), .B2(new_n1010), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1059), .A2(KEYINPUT112), .A3(new_n1052), .A4(new_n1054), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1052), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT52), .ZN(new_n1063));
  NAND2_X1  g638(.A1(G305), .A2(G1981), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n590), .A2(new_n706), .A3(new_n595), .A4(new_n591), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT113), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT49), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT113), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1064), .A2(new_n1069), .A3(new_n1065), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1067), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  OR3_X1    g646(.A1(new_n1066), .A2(KEYINPUT114), .A3(new_n1068), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT114), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1071), .A2(new_n1072), .A3(new_n1059), .A4(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1061), .A2(new_n1063), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1041), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1028), .A2(KEYINPUT45), .ZN(new_n1077));
  AOI21_X1  g652(.A(G1966), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1010), .B1(new_n1028), .B2(new_n1034), .ZN(new_n1079));
  AOI211_X1 g654(.A(KEYINPUT50), .B(G1384), .C1(new_n493), .C2(new_n505), .ZN(new_n1080));
  NOR3_X1   g655(.A1(new_n1079), .A2(G2084), .A3(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(G8), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1075), .A2(G286), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1027), .B1(new_n1050), .B2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n833), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1085));
  INV_X1    g660(.A(G2084), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1033), .A2(new_n1086), .A3(new_n1010), .A4(new_n1035), .ZN(new_n1087));
  AOI211_X1 g662(.A(new_n1058), .B(G286), .C1(new_n1085), .C2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1058), .B1(new_n1031), .B2(new_n1036), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1088), .B(new_n1027), .C1(new_n1048), .C2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1044), .A2(G8), .A3(new_n1048), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1075), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(G288), .A2(G1976), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1074), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT116), .ZN(new_n1095));
  XOR2_X1   g670(.A(new_n1065), .B(KEYINPUT115), .Z(new_n1096));
  AND3_X1   g671(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1095), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1059), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n1084), .A2(new_n1092), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT51), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1058), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n1104));
  NAND3_X1  g679(.A1(G286), .A2(new_n1104), .A3(G8), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1104), .B1(G286), .B2(G8), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1102), .B1(new_n1103), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT122), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1107), .ZN(new_n1112));
  NAND2_X1  g687(.A1(KEYINPUT122), .A2(KEYINPUT51), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1112), .A2(new_n1105), .A3(new_n1113), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1082), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1108), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1110), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1031), .A2(new_n1036), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1048), .B1(new_n1120), .B2(G8), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1121), .A2(new_n1075), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1119), .A2(new_n1091), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT54), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n1029), .A2(G2078), .A3(new_n1030), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1033), .A2(new_n1010), .A3(new_n1035), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n1125), .A2(KEYINPUT53), .B1(new_n1126), .B2(new_n851), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1128));
  INV_X1    g703(.A(G2078), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1128), .A2(new_n1129), .A3(new_n1077), .A4(new_n1010), .ZN(new_n1130));
  XOR2_X1   g705(.A(KEYINPUT123), .B(KEYINPUT53), .Z(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(G301), .B1(new_n1127), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1126), .A2(new_n851), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1076), .A2(KEYINPUT53), .A3(new_n1129), .A4(new_n1077), .ZN(new_n1135));
  AND4_X1   g710(.A1(G301), .A2(new_n1132), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1124), .B1(new_n1133), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT124), .ZN(new_n1138));
  OR3_X1    g713(.A1(new_n1133), .A2(new_n1136), .A3(new_n1124), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT124), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1140), .B(new_n1124), .C1(new_n1133), .C2(new_n1136), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1123), .A2(new_n1138), .A3(new_n1139), .A4(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT117), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n582), .A2(new_n1143), .ZN(new_n1144));
  OR2_X1    g719(.A1(new_n573), .A2(new_n574), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n566), .A2(new_n564), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n579), .A2(KEYINPUT117), .A3(new_n581), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .A4(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT118), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT57), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n583), .A2(KEYINPUT57), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1149), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g730(.A(KEYINPUT56), .B(G2072), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1076), .A2(new_n1077), .A3(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n829), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(G1348), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1160), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1028), .A2(new_n1015), .A3(new_n1010), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  AOI22_X1  g738(.A1(new_n1155), .A2(new_n1159), .B1(new_n1163), .B2(new_n620), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1158), .B(new_n1157), .C1(new_n1153), .C2(new_n1154), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(KEYINPUT119), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(KEYINPUT117), .B1(new_n579), .B2(new_n581), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n575), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(KEYINPUT57), .B1(new_n1169), .B2(new_n1147), .ZN(new_n1170));
  AOI22_X1  g745(.A1(new_n1170), .A2(new_n1149), .B1(KEYINPUT57), .B2(new_n583), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1154), .ZN(new_n1172));
  AOI21_X1  g747(.A(G1956), .B1(new_n1042), .B2(new_n1035), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1156), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1029), .A2(new_n1030), .A3(new_n1174), .ZN(new_n1175));
  OAI211_X1 g750(.A(new_n1171), .B(new_n1172), .C1(new_n1173), .C2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1163), .A2(new_n620), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT119), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1178), .A2(new_n1179), .A3(new_n1165), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1167), .A2(new_n1180), .ZN(new_n1181));
  AND3_X1   g756(.A1(new_n1176), .A2(KEYINPUT61), .A3(new_n1165), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT60), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n620), .B1(new_n1163), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(KEYINPUT60), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(KEYINPUT61), .B1(new_n1176), .B2(new_n1165), .ZN(new_n1187));
  NOR3_X1   g762(.A1(new_n1182), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1076), .A2(new_n1017), .A3(new_n1077), .ZN(new_n1189));
  XOR2_X1   g764(.A(KEYINPUT58), .B(G1341), .Z(new_n1190));
  NAND2_X1  g765(.A1(new_n1051), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT120), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1051), .A2(KEYINPUT120), .A3(new_n1190), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1189), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  AND3_X1   g770(.A1(new_n1195), .A2(KEYINPUT59), .A3(new_n555), .ZN(new_n1196));
  AOI21_X1  g771(.A(KEYINPUT59), .B1(new_n1195), .B2(new_n555), .ZN(new_n1197));
  NOR3_X1   g772(.A1(new_n1163), .A2(new_n620), .A3(new_n1183), .ZN(new_n1198));
  NOR3_X1   g773(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1181), .B1(new_n1188), .B2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1101), .B1(new_n1142), .B2(new_n1200), .ZN(new_n1201));
  AND2_X1   g776(.A1(new_n1122), .A2(new_n1091), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1117), .B1(new_n1082), .B2(new_n1115), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT62), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1203), .A2(new_n1204), .A3(new_n1110), .ZN(new_n1205));
  NAND4_X1  g780(.A1(new_n1202), .A2(KEYINPUT125), .A3(new_n1205), .A4(new_n1133), .ZN(new_n1206));
  INV_X1    g781(.A(KEYINPUT125), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1122), .A2(new_n1091), .A3(new_n1133), .ZN(new_n1208));
  AND3_X1   g783(.A1(new_n1203), .A2(new_n1204), .A3(new_n1110), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1207), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1119), .A2(KEYINPUT62), .ZN(new_n1211));
  AND3_X1   g786(.A1(new_n1206), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1026), .B1(new_n1201), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1011), .B1(new_n1016), .B2(new_n793), .ZN(new_n1214));
  OAI21_X1  g789(.A(KEYINPUT46), .B1(new_n1011), .B2(G1996), .ZN(new_n1215));
  OR3_X1    g790(.A1(new_n1011), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1214), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  XOR2_X1   g792(.A(new_n1217), .B(KEYINPUT47), .Z(new_n1218));
  AOI22_X1  g793(.A1(new_n1020), .A2(new_n1022), .B1(new_n1015), .B2(new_n910), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1218), .B1(new_n1219), .B2(new_n1011), .ZN(new_n1220));
  NAND3_X1  g795(.A1(new_n1020), .A2(KEYINPUT126), .A3(new_n1023), .ZN(new_n1221));
  NOR3_X1   g796(.A1(new_n1011), .A2(G1986), .A3(G290), .ZN(new_n1222));
  XNOR2_X1  g797(.A(new_n1222), .B(KEYINPUT127), .ZN(new_n1223));
  XNOR2_X1  g798(.A(new_n1223), .B(KEYINPUT48), .ZN(new_n1224));
  AOI21_X1  g799(.A(KEYINPUT126), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1225));
  NOR2_X1   g800(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g801(.A(new_n1220), .B1(new_n1221), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1213), .A2(new_n1227), .ZN(G329));
  assign    G231 = 1'b0;
  OAI211_X1 g803(.A(new_n684), .B(G319), .C1(new_n668), .C2(new_n667), .ZN(new_n1230));
  NOR2_X1   g804(.A1(G229), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g805(.A1(new_n921), .A2(new_n923), .ZN(new_n1232));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n995), .ZN(new_n1233));
  AND3_X1   g807(.A1(new_n1231), .A2(new_n1232), .A3(new_n1233), .ZN(G308));
  NAND3_X1  g808(.A1(new_n1231), .A2(new_n1232), .A3(new_n1233), .ZN(G225));
endmodule


