//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 1 1 0 0 0 1 1 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1301, new_n1302, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1359,
    new_n1360, new_n1361;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  NOR3_X1   g0004(.A1(new_n202), .A2(G77), .A3(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT65), .Z(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND3_X1  g0015(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n204), .A2(G50), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT66), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G50), .A2(G226), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G116), .A2(G270), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(KEYINPUT66), .B1(new_n218), .B2(new_n219), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n212), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n226), .C2(KEYINPUT1), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G264), .B(G270), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT67), .Z(new_n232));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n232), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G87), .B(G97), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XOR2_X1   g0043(.A(G50), .B(G58), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  OR2_X1    g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  NAND4_X1  g0048(.A1(new_n247), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT77), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AND2_X1   g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND4_X1  g0054(.A1(new_n254), .A2(KEYINPUT77), .A3(KEYINPUT7), .A4(new_n210), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n247), .A2(new_n210), .A3(new_n248), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT7), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n251), .A2(new_n255), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G68), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n210), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G159), .ZN(new_n263));
  OAI21_X1  g0063(.A(KEYINPUT78), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT78), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(new_n266), .A3(G159), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G58), .ZN(new_n269));
  INV_X1    g0069(.A(G68), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(G20), .B1(new_n271), .B2(new_n203), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n260), .A2(KEYINPUT16), .A3(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT16), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n270), .B1(new_n258), .B2(new_n249), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n276), .B1(new_n277), .B2(new_n273), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G1), .A2(G13), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n275), .A2(new_n278), .A3(new_n281), .ZN(new_n282));
  OR2_X1    g0082(.A1(KEYINPUT70), .A2(G1), .ZN(new_n283));
  NAND2_X1  g0083(.A1(KEYINPUT70), .A2(G1), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n283), .A2(G13), .A3(G20), .A4(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT8), .B(G58), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AND2_X1   g0088(.A1(KEYINPUT70), .A2(G1), .ZN(new_n289));
  NOR2_X1   g0089(.A1(KEYINPUT70), .A2(G1), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n281), .ZN(new_n293));
  INV_X1    g0093(.A(new_n287), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n288), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n282), .A2(new_n297), .ZN(new_n298));
  OR2_X1    g0098(.A1(KEYINPUT69), .A2(G41), .ZN(new_n299));
  NAND2_X1  g0099(.A1(KEYINPUT69), .A2(G41), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n209), .B(G274), .C1(new_n301), .C2(G45), .ZN(new_n302));
  INV_X1    g0102(.A(G41), .ZN(new_n303));
  OAI211_X1 g0103(.A(G1), .B(G13), .C1(new_n261), .C2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n283), .A2(new_n284), .ZN(new_n305));
  NOR2_X1   g0105(.A1(G41), .A2(G45), .ZN(new_n306));
  OAI211_X1 g0106(.A(G232), .B(new_n304), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT80), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT80), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n302), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT71), .B(G179), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  OAI211_X1 g0115(.A(G226), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT79), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n247), .A2(new_n248), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n319), .A2(KEYINPUT79), .A3(G226), .A4(G1698), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G1698), .ZN(new_n322));
  OAI211_X1 g0122(.A(G223), .B(new_n322), .C1(new_n252), .C2(new_n253), .ZN(new_n323));
  NAND2_X1  g0123(.A1(G33), .A2(G87), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n321), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n280), .B1(G33), .B2(G41), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n315), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n323), .A2(new_n324), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n328), .B1(new_n318), .B2(new_n320), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n302), .B(new_n307), .C1(new_n329), .C2(new_n304), .ZN(new_n330));
  INV_X1    g0130(.A(G169), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n313), .A2(new_n327), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n298), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT18), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n333), .B(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n308), .B1(new_n325), .B2(new_n326), .ZN(new_n336));
  INV_X1    g0136(.A(G190), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(new_n329), .B2(new_n304), .ZN(new_n338));
  OAI22_X1  g0138(.A1(new_n336), .A2(G200), .B1(new_n312), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n339), .A2(new_n282), .A3(new_n297), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n340), .B(KEYINPUT17), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n335), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT72), .ZN(new_n343));
  INV_X1    g0143(.A(new_n306), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n326), .B1(new_n291), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G226), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n346), .A2(new_n302), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n319), .A2(G222), .A3(new_n322), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n319), .A2(G223), .A3(G1698), .ZN(new_n349));
  INV_X1    g0149(.A(G77), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n348), .B(new_n349), .C1(new_n350), .C2(new_n319), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n326), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n343), .B1(new_n353), .B2(new_n315), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n285), .A2(new_n293), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n356), .A2(G50), .A3(new_n292), .ZN(new_n357));
  INV_X1    g0157(.A(G50), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n286), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n210), .A2(G33), .ZN(new_n360));
  INV_X1    g0160(.A(G150), .ZN(new_n361));
  OAI22_X1  g0161(.A1(new_n287), .A2(new_n360), .B1(new_n361), .B2(new_n262), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n210), .B1(new_n201), .B2(new_n203), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n281), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n357), .A2(new_n359), .A3(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n347), .A2(KEYINPUT72), .A3(new_n352), .A4(new_n314), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n353), .A2(new_n331), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n354), .A2(new_n365), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(G232), .A2(G1698), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n322), .A2(G238), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n319), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n371), .B(new_n326), .C1(G107), .C2(new_n319), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n345), .A2(G244), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n372), .A2(new_n302), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G190), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n285), .A2(G77), .ZN(new_n377));
  XNOR2_X1  g0177(.A(new_n377), .B(KEYINPUT73), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n305), .A2(new_n210), .ZN(new_n379));
  NOR3_X1   g0179(.A1(new_n355), .A2(new_n379), .A3(new_n350), .ZN(new_n380));
  NAND2_X1  g0180(.A1(G20), .A2(G77), .ZN(new_n381));
  XNOR2_X1  g0181(.A(KEYINPUT15), .B(G87), .ZN(new_n382));
  OAI221_X1 g0182(.A(new_n381), .B1(new_n287), .B2(new_n262), .C1(new_n360), .C2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n380), .B1(new_n281), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n374), .A2(G200), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n376), .A2(new_n378), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n375), .A2(new_n314), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n384), .A2(new_n378), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n374), .A2(new_n331), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  OR2_X1    g0191(.A1(new_n365), .A2(KEYINPUT9), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n365), .A2(KEYINPUT9), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n392), .A2(new_n393), .B1(G200), .B2(new_n353), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT10), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT74), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n353), .B2(new_n337), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n347), .A2(KEYINPUT74), .A3(new_n352), .A4(G190), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AND3_X1   g0199(.A1(new_n394), .A2(new_n395), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n395), .B1(new_n394), .B2(new_n399), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n368), .B(new_n391), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n356), .A2(G68), .A3(new_n292), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n265), .A2(G50), .B1(G20), .B2(new_n270), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(new_n350), .B2(new_n360), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT11), .ZN(new_n406));
  AND3_X1   g0206(.A1(new_n405), .A2(new_n406), .A3(new_n281), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n406), .B1(new_n405), .B2(new_n281), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n403), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n285), .A2(G68), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n410), .B(KEYINPUT12), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n412), .A2(KEYINPUT76), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT76), .ZN(new_n414));
  NOR3_X1   g0214(.A1(new_n409), .A2(new_n414), .A3(new_n411), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n345), .A2(G238), .ZN(new_n417));
  NOR2_X1   g0217(.A1(G226), .A2(G1698), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n418), .B1(new_n234), .B2(G1698), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n419), .A2(new_n319), .B1(G33), .B2(G97), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n417), .B(new_n302), .C1(new_n304), .C2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT13), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n420), .A2(new_n304), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT13), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n423), .A2(new_n424), .A3(new_n302), .A4(new_n417), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n422), .A2(new_n425), .A3(G179), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n331), .B1(new_n422), .B2(new_n425), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT75), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT14), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n426), .B1(new_n427), .B2(new_n431), .ZN(new_n432));
  AOI211_X1 g0232(.A(new_n331), .B(new_n430), .C1(new_n422), .C2(new_n425), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n416), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AND2_X1   g0234(.A1(new_n422), .A2(new_n425), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(G190), .ZN(new_n436));
  INV_X1    g0236(.A(G200), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n436), .B(new_n412), .C1(new_n437), .C2(new_n435), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  NOR3_X1   g0239(.A1(new_n342), .A2(new_n402), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT5), .ZN(new_n442));
  AND2_X1   g0242(.A1(KEYINPUT69), .A2(G41), .ZN(new_n443));
  NOR2_X1   g0243(.A1(KEYINPUT69), .A2(G41), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n303), .A2(KEYINPUT5), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n445), .A2(G45), .A3(new_n291), .A4(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n447), .A2(G264), .A3(new_n304), .ZN(new_n448));
  OAI211_X1 g0248(.A(G257), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n449));
  OAI211_X1 g0249(.A(G250), .B(new_n322), .C1(new_n252), .C2(new_n253), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G294), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n326), .ZN(new_n453));
  AND3_X1   g0253(.A1(new_n448), .A2(new_n453), .A3(KEYINPUT93), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT93), .B1(new_n448), .B2(new_n453), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n304), .A2(G274), .A3(new_n446), .ZN(new_n456));
  AOI21_X1  g0256(.A(KEYINPUT5), .B1(new_n299), .B2(new_n300), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n283), .A2(G45), .A3(new_n284), .ZN(new_n458));
  OAI21_X1  g0258(.A(KEYINPUT83), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(G45), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n289), .A2(new_n290), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT83), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n461), .A2(new_n462), .A3(new_n445), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n456), .B1(new_n459), .B2(new_n463), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n454), .A2(new_n455), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n456), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n457), .A2(new_n458), .A3(KEYINPUT83), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n462), .B1(new_n461), .B2(new_n445), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n469), .A2(new_n448), .A3(new_n453), .ZN(new_n470));
  OAI22_X1  g0270(.A1(new_n465), .A2(G200), .B1(G190), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT95), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n285), .A2(G107), .ZN(new_n473));
  OR2_X1    g0273(.A1(new_n473), .A2(KEYINPUT25), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(KEYINPUT25), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G107), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n291), .A2(G33), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n356), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n476), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT24), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n319), .A2(new_n210), .A3(G87), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT22), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT22), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n319), .A2(new_n484), .A3(new_n210), .A4(G87), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(G116), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n360), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT23), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n489), .B1(new_n210), .B2(G107), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n477), .A2(KEYINPUT23), .A3(G20), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n481), .B1(new_n486), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n486), .A2(new_n481), .A3(new_n492), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n480), .B1(new_n496), .B2(new_n281), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n471), .A2(new_n472), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n448), .A2(new_n453), .ZN(new_n499));
  NOR3_X1   g0299(.A1(new_n499), .A2(G190), .A3(new_n464), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT93), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n448), .A2(new_n453), .A3(KEYINPUT93), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n502), .A2(new_n469), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n500), .B1(new_n504), .B2(new_n437), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n486), .A2(new_n481), .A3(new_n492), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n281), .B1(new_n506), .B2(new_n493), .ZN(new_n507));
  INV_X1    g0307(.A(new_n479), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n508), .A2(G107), .B1(new_n474), .B2(new_n475), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(KEYINPUT95), .B1(new_n505), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n498), .A2(new_n511), .ZN(new_n512));
  AND2_X1   g0312(.A1(KEYINPUT4), .A2(G244), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n322), .B(new_n513), .C1(new_n252), .C2(new_n253), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G283), .ZN(new_n515));
  INV_X1    g0315(.A(G244), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n516), .B1(new_n247), .B2(new_n248), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n514), .B(new_n515), .C1(new_n517), .C2(KEYINPUT4), .ZN(new_n518));
  OAI21_X1  g0318(.A(G250), .B1(new_n252), .B2(new_n253), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n322), .B1(new_n519), .B2(KEYINPUT4), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n326), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n447), .A2(G257), .A3(new_n304), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n469), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT85), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n469), .A2(new_n521), .A3(KEYINPUT85), .A4(new_n522), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n525), .A2(new_n331), .A3(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n522), .ZN(new_n528));
  NOR3_X1   g0328(.A1(new_n528), .A2(new_n464), .A3(KEYINPUT84), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT84), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n530), .B1(new_n469), .B2(new_n522), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n314), .B(new_n521), .C1(new_n529), .C2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT6), .ZN(new_n533));
  NOR3_X1   g0333(.A1(new_n533), .A2(G97), .A3(G107), .ZN(new_n534));
  INV_X1    g0334(.A(G97), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n535), .A2(KEYINPUT6), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT81), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n537), .A2(G107), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n477), .A2(KEYINPUT81), .ZN(new_n539));
  OAI22_X1  g0339(.A1(new_n534), .A2(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(G97), .A2(G107), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT6), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n533), .A2(G97), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n477), .A2(KEYINPUT81), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n537), .A2(G107), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n542), .A2(new_n543), .A3(new_n544), .A4(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n540), .A2(G20), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n265), .A2(G77), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n547), .A2(KEYINPUT82), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n258), .A2(new_n249), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G107), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT82), .B1(new_n547), .B2(new_n548), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n281), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n285), .A2(G97), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n555), .B1(new_n508), .B2(G97), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n527), .A2(new_n532), .A3(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n521), .B1(new_n529), .B2(new_n531), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(G200), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n528), .A2(new_n464), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT85), .B1(new_n561), .B2(new_n521), .ZN(new_n562));
  INV_X1    g0362(.A(new_n526), .ZN(new_n563));
  OAI21_X1  g0363(.A(G190), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n554), .A2(new_n556), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n560), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT88), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n210), .B(G68), .C1(new_n252), .C2(new_n253), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT19), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n360), .B2(new_n535), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  OR2_X1    g0371(.A1(KEYINPUT87), .A2(G87), .ZN(new_n572));
  NAND2_X1  g0372(.A1(KEYINPUT87), .A2(G87), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n572), .A2(new_n541), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n210), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n293), .B1(new_n571), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n382), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n579), .A2(new_n285), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n567), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n577), .A2(new_n570), .A3(new_n568), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n281), .ZN(new_n583));
  INV_X1    g0383(.A(new_n580), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n583), .A2(KEYINPUT88), .A3(new_n584), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n581), .A2(new_n585), .B1(new_n579), .B2(new_n508), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(G274), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n283), .A2(G45), .A3(new_n588), .A4(new_n284), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n304), .B(new_n589), .C1(new_n461), .C2(G250), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(KEYINPUT86), .ZN(new_n591));
  INV_X1    g0391(.A(G250), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n326), .B1(new_n458), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT86), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n593), .A2(new_n594), .A3(new_n589), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(G238), .B(new_n322), .C1(new_n252), .C2(new_n253), .ZN(new_n597));
  OAI211_X1 g0397(.A(G244), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n597), .B(new_n598), .C1(new_n261), .C2(new_n487), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n326), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n596), .A2(new_n314), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(G169), .B1(new_n596), .B2(new_n600), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI221_X4 g0403(.A(new_n337), .B1(new_n326), .B2(new_n599), .C1(new_n591), .C2(new_n595), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n437), .B1(new_n596), .B2(new_n600), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n478), .A2(G87), .A3(new_n293), .A4(new_n285), .ZN(new_n607));
  XNOR2_X1  g0407(.A(new_n607), .B(KEYINPUT89), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n608), .B1(new_n585), .B2(new_n581), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n587), .A2(new_n603), .B1(new_n606), .B2(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n512), .A2(new_n558), .A3(new_n566), .A4(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT91), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n447), .A2(G270), .A3(new_n304), .ZN(new_n613));
  OAI211_X1 g0413(.A(G264), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n614));
  OAI211_X1 g0414(.A(G257), .B(new_n322), .C1(new_n252), .C2(new_n253), .ZN(new_n615));
  INV_X1    g0415(.A(G303), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n614), .B(new_n615), .C1(new_n616), .C2(new_n319), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n326), .ZN(new_n618));
  AND4_X1   g0418(.A1(G179), .A2(new_n469), .A3(new_n613), .A4(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n459), .A2(new_n463), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n620), .A2(new_n466), .B1(new_n326), .B2(new_n617), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n331), .B1(new_n621), .B2(new_n613), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n619), .B1(new_n622), .B2(KEYINPUT21), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n478), .A2(G116), .A3(new_n293), .A4(new_n285), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n286), .A2(new_n487), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n515), .B(new_n210), .C1(G33), .C2(new_n535), .ZN(new_n627));
  AOI221_X4 g0427(.A(KEYINPUT90), .B1(new_n487), .B2(G20), .C1(new_n279), .C2(new_n280), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT90), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n487), .A2(G20), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n629), .B1(new_n281), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n627), .B1(new_n628), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT20), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI211_X1 g0434(.A(KEYINPUT20), .B(new_n627), .C1(new_n628), .C2(new_n631), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n626), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n612), .B1(new_n623), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n469), .A2(new_n613), .A3(new_n618), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n638), .A2(KEYINPUT21), .A3(G169), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n621), .A2(G179), .A3(new_n613), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n626), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n281), .A2(new_n630), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(KEYINPUT90), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n281), .A2(new_n629), .A3(new_n630), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(KEYINPUT20), .B1(new_n646), .B2(new_n627), .ZN(new_n647));
  INV_X1    g0447(.A(new_n635), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n642), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n641), .A2(KEYINPUT91), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n637), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n502), .A2(G179), .A3(new_n469), .A4(new_n503), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n470), .A2(G169), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT94), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n652), .A2(KEYINPUT94), .A3(new_n653), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(new_n510), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT21), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n638), .A2(G169), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(new_n636), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT92), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n649), .A2(G169), .A3(new_n638), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n664), .A2(KEYINPUT92), .A3(new_n659), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n638), .A2(G200), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n621), .A2(G190), .A3(new_n613), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(new_n668), .A3(new_n636), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n651), .A2(new_n658), .A3(new_n666), .A4(new_n669), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n441), .A2(new_n611), .A3(new_n670), .ZN(G372));
  INV_X1    g0471(.A(new_n368), .ZN(new_n672));
  INV_X1    g0472(.A(new_n434), .ZN(new_n673));
  INV_X1    g0473(.A(new_n390), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n673), .B1(new_n438), .B2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n341), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n335), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n400), .A2(new_n401), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n672), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n591), .A2(new_n595), .B1(new_n326), .B2(new_n599), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n314), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(G169), .B2(new_n680), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(new_n586), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n527), .A2(new_n532), .A3(new_n557), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n610), .A2(new_n684), .A3(KEYINPUT26), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT26), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n596), .A2(G190), .A3(new_n600), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n680), .B2(new_n437), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT89), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n607), .B(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(KEYINPUT88), .B1(new_n583), .B2(new_n584), .ZN(new_n691));
  AOI211_X1 g0491(.A(new_n567), .B(new_n580), .C1(new_n582), .C2(new_n281), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OAI22_X1  g0493(.A1(new_n682), .A2(new_n586), .B1(new_n688), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n686), .B1(new_n694), .B2(new_n558), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n683), .B1(new_n685), .B2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n641), .A2(new_n649), .ZN(new_n698));
  AOI211_X1 g0498(.A(new_n662), .B(KEYINPUT21), .C1(new_n622), .C2(new_n649), .ZN(new_n699));
  AOI21_X1  g0499(.A(KEYINPUT92), .B1(new_n664), .B2(new_n659), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT96), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n666), .A2(KEYINPUT96), .A3(new_n698), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n510), .A2(new_n654), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT97), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n611), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n703), .A2(new_n704), .A3(KEYINPUT97), .A4(new_n705), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n697), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n679), .B1(new_n710), .B2(new_n441), .ZN(G369));
  INV_X1    g0511(.A(new_n669), .ZN(new_n712));
  AOI21_X1  g0512(.A(KEYINPUT91), .B1(new_n641), .B2(new_n649), .ZN(new_n713));
  AOI211_X1 g0513(.A(new_n612), .B(new_n636), .C1(new_n639), .C2(new_n640), .ZN(new_n714));
  OAI22_X1  g0514(.A1(new_n713), .A2(new_n714), .B1(new_n699), .B2(new_n700), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n210), .A2(G13), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n291), .A2(new_n716), .ZN(new_n717));
  OR2_X1    g0517(.A1(new_n717), .A2(KEYINPUT27), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(KEYINPUT27), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(G213), .A3(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(G343), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI211_X1 g0522(.A(new_n712), .B(new_n715), .C1(new_n649), .C2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n722), .ZN(new_n724));
  AOI211_X1 g0524(.A(new_n636), .B(new_n724), .C1(new_n703), .C2(new_n704), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(G330), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n657), .ZN(new_n729));
  AOI21_X1  g0529(.A(KEYINPUT94), .B1(new_n652), .B2(new_n653), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n729), .A2(new_n730), .A3(new_n497), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n731), .B1(new_n510), .B2(new_n722), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n512), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(new_n658), .B2(new_n724), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n728), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n722), .B1(new_n651), .B2(new_n666), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n732), .A2(new_n736), .A3(new_n512), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n510), .A2(new_n654), .A3(new_n724), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n735), .A2(new_n740), .ZN(G399));
  INV_X1    g0541(.A(new_n213), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n301), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n574), .A2(G116), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n744), .A2(G1), .A3(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n217), .ZN(new_n748));
  AOI22_X1  g0548(.A1(new_n747), .A2(KEYINPUT98), .B1(new_n748), .B2(new_n743), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n749), .B1(KEYINPUT98), .B2(new_n747), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT28), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n715), .A2(new_n731), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n696), .B1(new_n611), .B2(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n753), .A2(KEYINPUT29), .A3(new_n724), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n706), .A2(new_n707), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n566), .A2(new_n610), .A3(new_n558), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n756), .B1(new_n498), .B2(new_n511), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n755), .A2(new_n757), .A3(new_n709), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n722), .B1(new_n758), .B2(new_n696), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n754), .B1(new_n759), .B2(KEYINPUT29), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n715), .A2(new_n731), .A3(new_n712), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n757), .A2(new_n761), .A3(new_n724), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT30), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n562), .A2(new_n563), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n619), .A2(new_n502), .A3(new_n503), .A4(new_n680), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n525), .A2(new_n526), .ZN(new_n767));
  AND3_X1   g0567(.A1(new_n502), .A2(new_n680), .A3(new_n503), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n767), .A2(new_n768), .A3(KEYINPUT30), .A4(new_n619), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n638), .A2(new_n314), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT99), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(new_n596), .B2(new_n600), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n680), .A2(new_n771), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n773), .A2(new_n559), .A3(new_n504), .A4(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n766), .A2(new_n769), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n722), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(KEYINPUT31), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT31), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n776), .A2(new_n779), .A3(new_n722), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n727), .B1(new_n762), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n760), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT100), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n760), .A2(KEYINPUT100), .A3(new_n783), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n751), .B1(new_n788), .B2(G1), .ZN(G364));
  NAND2_X1  g0589(.A1(new_n728), .A2(KEYINPUT101), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT101), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(new_n726), .B2(new_n727), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n209), .B1(new_n716), .B2(G45), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n743), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n795), .B1(new_n726), .B2(new_n727), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n790), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n213), .A2(new_n319), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n798), .A2(new_n207), .B1(G116), .B2(new_n213), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n245), .A2(G45), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n213), .A2(new_n254), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(new_n460), .B2(new_n748), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n799), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(G13), .A2(G33), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(G20), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n280), .B1(G20), .B2(new_n331), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n795), .B1(new_n803), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n337), .A2(G20), .ZN(new_n811));
  AOI21_X1  g0611(.A(G179), .B1(new_n811), .B2(KEYINPUT102), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(KEYINPUT102), .B2(new_n811), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n437), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G283), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR4_X1   g0617(.A1(new_n210), .A2(new_n337), .A3(new_n437), .A4(G179), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n254), .B1(new_n819), .B2(new_n616), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n811), .A2(new_n437), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n315), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  XNOR2_X1  g0623(.A(KEYINPUT33), .B(G317), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n820), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(G294), .ZN(new_n826));
  INV_X1    g0626(.A(G179), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n827), .A2(new_n437), .A3(G190), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(G20), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n825), .B1(new_n826), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n813), .A2(G200), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n817), .B(new_n831), .C1(G329), .C2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n315), .A2(G20), .ZN(new_n834));
  NOR3_X1   g0634(.A1(new_n834), .A2(new_n337), .A3(G200), .ZN(new_n835));
  NOR3_X1   g0635(.A1(new_n834), .A2(new_n337), .A3(new_n437), .ZN(new_n836));
  AOI22_X1  g0636(.A1(G322), .A2(new_n835), .B1(new_n836), .B2(G326), .ZN(new_n837));
  INV_X1    g0637(.A(G311), .ZN(new_n838));
  NOR3_X1   g0638(.A1(new_n834), .A2(G190), .A3(G200), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n833), .B(new_n837), .C1(new_n838), .C2(new_n840), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n572), .A2(new_n573), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n319), .B1(new_n819), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n835), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n269), .A2(new_n844), .B1(new_n840), .B2(new_n350), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n843), .B(new_n845), .C1(G50), .C2(new_n836), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n830), .A2(new_n535), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(new_n823), .B2(G68), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT103), .Z(new_n849));
  NAND2_X1  g0649(.A1(new_n814), .A2(G107), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n846), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n832), .A2(G159), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT32), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n841), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n810), .B1(new_n854), .B2(new_n807), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT104), .ZN(new_n856));
  INV_X1    g0656(.A(new_n726), .ZN(new_n857));
  INV_X1    g0657(.A(new_n806), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n797), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(G396));
  NAND2_X1  g0661(.A1(new_n388), .A2(new_n722), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n386), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n390), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n674), .A2(new_n724), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n391), .A2(new_n724), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n759), .A2(new_n867), .B1(new_n710), .B2(new_n868), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n869), .A2(new_n783), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n795), .B1(new_n869), .B2(new_n783), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n807), .A2(new_n804), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n795), .B1(G77), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n807), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n836), .A2(G137), .B1(G150), .B2(new_n823), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n877), .B(KEYINPUT105), .ZN(new_n878));
  INV_X1    g0678(.A(G143), .ZN(new_n879));
  OAI221_X1 g0679(.A(new_n878), .B1(new_n879), .B2(new_n844), .C1(new_n263), .C2(new_n840), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT34), .ZN(new_n881));
  OR2_X1    g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n880), .A2(new_n881), .ZN(new_n883));
  OAI221_X1 g0683(.A(new_n319), .B1(new_n830), .B2(new_n269), .C1(new_n819), .C2(new_n358), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n815), .A2(new_n270), .ZN(new_n885));
  AOI211_X1 g0685(.A(new_n884), .B(new_n885), .C1(G132), .C2(new_n832), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n882), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n836), .ZN(new_n888));
  OAI22_X1  g0688(.A1(new_n826), .A2(new_n844), .B1(new_n888), .B2(new_n616), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(G116), .B2(new_n839), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n254), .B1(new_n819), .B2(new_n477), .ZN(new_n891));
  AOI211_X1 g0691(.A(new_n847), .B(new_n891), .C1(G283), .C2(new_n823), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n832), .A2(G311), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n814), .A2(G87), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n890), .A2(new_n892), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n876), .B1(new_n887), .B2(new_n895), .ZN(new_n896));
  AOI211_X1 g0696(.A(new_n875), .B(new_n896), .C1(new_n804), .C2(new_n866), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n872), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(G384));
  NOR2_X1   g0699(.A1(new_n216), .A2(new_n487), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n540), .A2(new_n546), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT35), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n903), .B1(new_n902), .B2(new_n901), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n904), .B(KEYINPUT36), .ZN(new_n905));
  OR3_X1    g0705(.A1(new_n217), .A2(new_n350), .A3(new_n271), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n201), .A2(G68), .ZN(new_n907));
  AOI211_X1 g0707(.A(G13), .B(new_n291), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT38), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT108), .ZN(new_n911));
  INV_X1    g0711(.A(new_n720), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT107), .B1(new_n298), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT107), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n914), .B(new_n720), .C1(new_n282), .C2(new_n297), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT37), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n333), .A2(new_n340), .A3(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n911), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n333), .A2(new_n340), .A3(new_n917), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n273), .B1(new_n259), .B2(G68), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n293), .B1(new_n921), .B2(KEYINPUT16), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n296), .B1(new_n922), .B2(new_n278), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n914), .B1(new_n923), .B2(new_n720), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n298), .A2(KEYINPUT107), .A3(new_n912), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n920), .A2(KEYINPUT108), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n926), .A2(new_n333), .A3(new_n340), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n919), .A2(new_n927), .B1(new_n928), .B2(KEYINPUT37), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n926), .B1(new_n335), .B2(new_n341), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n910), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n922), .B1(KEYINPUT16), .B2(new_n921), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n297), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n933), .A2(new_n912), .B1(new_n923), .B2(new_n339), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n332), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n917), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n916), .A2(new_n911), .A3(new_n918), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT108), .B1(new_n920), .B2(new_n926), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n933), .A2(new_n912), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n335), .B2(new_n341), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n940), .A2(new_n943), .A3(KEYINPUT38), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n931), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT39), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n673), .A2(new_n724), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n936), .B1(new_n919), .B2(new_n927), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n910), .B1(new_n950), .B2(new_n942), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n944), .A2(new_n951), .A3(KEYINPUT39), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n947), .A2(new_n949), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n944), .A2(new_n951), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n416), .A2(new_n722), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n434), .A2(new_n438), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n955), .B1(new_n434), .B2(new_n438), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n868), .B1(new_n758), .B2(new_n696), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n865), .B(KEYINPUT106), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n954), .B(new_n959), .C1(new_n960), .C2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n335), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n720), .ZN(new_n965));
  AND3_X1   g0765(.A1(new_n953), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n440), .B(new_n754), .C1(new_n759), .C2(KEYINPUT29), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n967), .A2(new_n679), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n966), .B(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n867), .B1(new_n956), .B2(new_n957), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(new_n762), .B2(new_n781), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n954), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT40), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n973), .B(new_n970), .C1(new_n762), .C2(new_n781), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n972), .A2(new_n973), .B1(new_n945), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n441), .B1(new_n762), .B2(new_n781), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n976), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n977), .A2(G330), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n969), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n291), .B2(new_n716), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n969), .A2(new_n979), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n909), .B1(new_n981), .B2(new_n982), .ZN(G367));
  INV_X1    g0783(.A(new_n231), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n808), .B1(new_n213), .B2(new_n382), .C1(new_n984), .C2(new_n801), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n795), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n879), .A2(new_n888), .B1(new_n844), .B2(new_n361), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n830), .A2(new_n270), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n319), .B1(new_n819), .B2(new_n269), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n988), .B(new_n989), .C1(G159), .C2(new_n823), .ZN(new_n990));
  INV_X1    g0790(.A(G137), .ZN(new_n991));
  INV_X1    g0791(.A(new_n832), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n990), .B1(new_n350), .B2(new_n815), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n987), .B(new_n993), .C1(new_n202), .C2(new_n839), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT110), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n818), .A2(G116), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT46), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n995), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n888), .B2(new_n838), .C1(new_n816), .C2(new_n840), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n835), .A2(G303), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(KEYINPUT111), .B(KEYINPUT46), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n823), .A2(G294), .B1(new_n996), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n319), .B1(new_n829), .B2(G107), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n818), .A2(KEYINPUT110), .A3(KEYINPUT46), .A4(G116), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1000), .A2(new_n1002), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(G317), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n535), .A2(new_n815), .B1(new_n992), .B2(new_n1006), .ZN(new_n1007));
  NOR3_X1   g0807(.A1(new_n999), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n994), .A2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT47), .Z(new_n1010));
  AOI21_X1  g0810(.A(new_n986), .B1(new_n1010), .B2(new_n807), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n610), .B1(new_n609), .B2(new_n724), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n683), .A2(new_n693), .A3(new_n722), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1012), .A2(new_n806), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n566), .B(new_n558), .C1(new_n565), .C2(new_n724), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n684), .A2(new_n722), .ZN(new_n1017));
  AND2_X1   g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n737), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(KEYINPUT42), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n558), .B1(new_n1016), .B2(new_n658), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n724), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1023), .A2(KEYINPUT109), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1019), .A2(KEYINPUT42), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n1023), .B2(KEYINPUT109), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n1024), .A2(new_n1026), .B1(KEYINPUT43), .B2(new_n1027), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1027), .A2(KEYINPUT43), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1028), .B(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n735), .A2(new_n1018), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1030), .B(new_n1031), .Z(new_n1032));
  AND2_X1   g0832(.A1(new_n739), .A2(new_n1018), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT44), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n739), .A2(new_n1018), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT45), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n735), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1034), .A2(new_n735), .A3(new_n1036), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n734), .A2(new_n736), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n737), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1042), .A2(new_n790), .A3(new_n792), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1041), .A2(new_n728), .A3(new_n737), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n788), .B1(new_n1040), .B2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n743), .B(KEYINPUT41), .Z(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n794), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1015), .B1(new_n1032), .B2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT112), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(G387));
  INV_X1    g0852(.A(KEYINPUT115), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1045), .B1(new_n786), .B2(new_n787), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1054), .A2(new_n744), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n786), .A2(new_n1045), .A3(new_n787), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1045), .A2(new_n793), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n734), .A2(new_n858), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n237), .A2(new_n460), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n1060), .A2(new_n801), .B1(new_n745), .B2(new_n798), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n287), .A2(G50), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1062), .B(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1064), .A2(new_n745), .A3(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1061), .A2(new_n1066), .B1(new_n477), .B2(new_n742), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n795), .B1(new_n1067), .B2(new_n809), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n839), .A2(G68), .B1(new_n294), .B2(new_n823), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT114), .Z(new_n1070));
  NAND2_X1  g0870(.A1(new_n579), .A2(new_n829), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n819), .A2(new_n350), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1072), .A2(new_n254), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1071), .B(new_n1073), .C1(new_n844), .C2(new_n358), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(G159), .B2(new_n836), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(G97), .A2(new_n814), .B1(new_n832), .B2(G150), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1070), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n319), .B1(new_n832), .B2(G326), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n819), .A2(new_n826), .B1(new_n816), .B2(new_n830), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n836), .A2(G322), .B1(G311), .B2(new_n823), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1080), .B1(new_n616), .B2(new_n840), .C1(new_n1006), .C2(new_n844), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT48), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n1082), .B2(new_n1081), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT49), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1078), .B1(new_n487), .B2(new_n815), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1077), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1068), .B1(new_n1088), .B2(new_n807), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1058), .B1(new_n1059), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1053), .B1(new_n1057), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1057), .A2(new_n1053), .A3(new_n1090), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(G393));
  INV_X1    g0894(.A(new_n1040), .ZN(new_n1095));
  OR2_X1    g0895(.A1(new_n1095), .A2(KEYINPUT116), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(KEYINPUT116), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1096), .A2(new_n794), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n744), .B1(new_n1095), .B2(new_n1054), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n1054), .B2(new_n1095), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n242), .A2(new_n801), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n808), .B1(new_n535), .B2(new_n213), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n795), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(G150), .A2(new_n836), .B1(new_n835), .B2(G159), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT51), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n840), .A2(new_n287), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n822), .A2(new_n201), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n830), .A2(new_n350), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n319), .B1(new_n819), .B2(new_n270), .ZN(new_n1109));
  NOR4_X1   g0909(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n832), .A2(G143), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1110), .A2(new_n894), .A3(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n830), .A2(new_n487), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n254), .B1(new_n819), .B2(new_n816), .C1(new_n616), .C2(new_n822), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n1113), .B(new_n1114), .C1(G294), .C2(new_n839), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n832), .A2(G322), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1115), .A2(new_n850), .A3(new_n1116), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(G311), .A2(new_n835), .B1(new_n836), .B2(G317), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT52), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n1105), .A2(new_n1112), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1103), .B1(new_n1120), .B2(new_n807), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1018), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1121), .B1(new_n1122), .B2(new_n858), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1098), .A2(new_n1100), .A3(new_n1123), .ZN(G390));
  AOI211_X1 g0924(.A(new_n727), .B(new_n866), .C1(new_n762), .C2(new_n781), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n959), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n928), .A2(KEYINPUT37), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n938), .B2(new_n939), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n930), .ZN(new_n1130));
  AOI21_X1  g0930(.A(KEYINPUT38), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NOR3_X1   g0931(.A1(new_n950), .A2(new_n910), .A3(new_n942), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n948), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n753), .A2(new_n724), .A3(new_n867), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n958), .B1(new_n1134), .B2(new_n961), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT117), .ZN(new_n1136));
  NOR3_X1   g0936(.A1(new_n1133), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n658), .B(new_n666), .C1(new_n713), .C2(new_n714), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n566), .A2(new_n610), .A3(new_n558), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1138), .A2(new_n512), .A3(new_n1139), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n722), .B(new_n866), .C1(new_n1140), .C2(new_n696), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n959), .B1(new_n1141), .B2(new_n962), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n949), .B1(new_n931), .B2(new_n944), .ZN(new_n1143));
  AOI21_X1  g0943(.A(KEYINPUT117), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1137), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n959), .B1(new_n960), .B2(new_n962), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1146), .A2(new_n948), .B1(new_n947), .B2(new_n952), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1127), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1136), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1142), .A2(KEYINPUT117), .A3(new_n1143), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n944), .A2(new_n951), .A3(KEYINPUT39), .ZN(new_n1152));
  AOI21_X1  g0952(.A(KEYINPUT39), .B1(new_n931), .B2(new_n944), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n961), .B1(new_n710), .B2(new_n868), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n949), .B1(new_n1155), .B2(new_n959), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1151), .B(new_n1126), .C1(new_n1154), .C2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1148), .A2(new_n1157), .ZN(new_n1158));
  NOR3_X1   g0958(.A1(new_n611), .A2(new_n670), .A3(new_n722), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n776), .A2(new_n779), .A3(new_n722), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n779), .B1(new_n776), .B2(new_n722), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n440), .B(G330), .C1(new_n1159), .C2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT118), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n782), .A2(KEYINPUT118), .A3(new_n440), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n967), .A2(new_n679), .A3(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1125), .A2(new_n959), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1155), .B1(new_n1127), .B2(new_n1169), .ZN(new_n1170));
  OAI211_X1 g0970(.A(KEYINPUT119), .B(G330), .C1(new_n1159), .C2(new_n1162), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n867), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n782), .A2(KEYINPUT119), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n958), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1134), .A2(new_n961), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n1125), .B2(new_n959), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1168), .B1(new_n1170), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1158), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1148), .A2(new_n1178), .A3(new_n1157), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(new_n743), .A3(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1148), .A2(new_n794), .A3(new_n1157), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n795), .B1(new_n294), .B2(new_n874), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n487), .A2(new_n844), .B1(new_n888), .B2(new_n816), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G97), .B2(new_n839), .ZN(new_n1186));
  INV_X1    g0986(.A(G87), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n254), .B1(new_n819), .B2(new_n1187), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1108), .B(new_n1188), .C1(G107), .C2(new_n823), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n885), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n832), .A2(G294), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1186), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(G128), .A2(new_n836), .B1(new_n835), .B2(G132), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n819), .A2(KEYINPUT53), .A3(new_n361), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT53), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(new_n818), .B2(G150), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n1194), .A2(new_n254), .A3(new_n1196), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(G125), .A2(new_n832), .B1(new_n814), .B2(new_n202), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1193), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n823), .A2(G137), .B1(G159), .B2(new_n829), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(KEYINPUT54), .B(G143), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1200), .B1(new_n840), .B2(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT120), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1192), .B1(new_n1199), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1184), .B1(new_n1204), .B2(new_n807), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n1154), .B2(new_n805), .ZN(new_n1206));
  AND2_X1   g1006(.A1(new_n1183), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1182), .A2(new_n1207), .ZN(G378));
  INV_X1    g1008(.A(new_n1168), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1181), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT57), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n953), .A2(new_n963), .A3(new_n965), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n945), .A2(KEYINPUT40), .A3(new_n971), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n957), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n434), .A2(new_n438), .A3(new_n955), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n866), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n944), .B2(new_n951), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1213), .B(G330), .C1(new_n1218), .C2(KEYINPUT40), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n365), .A2(new_n912), .ZN(new_n1220));
  AND3_X1   g1020(.A1(new_n678), .A2(new_n368), .A3(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1220), .B1(new_n678), .B2(new_n368), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  OR3_X1    g1024(.A1(new_n1221), .A2(new_n1222), .A3(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1224), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1219), .A2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1227), .B1(new_n975), .B2(G330), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1212), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1219), .A2(new_n1228), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n975), .A2(G330), .A3(new_n1227), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n966), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1211), .B1(new_n1231), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1210), .A2(new_n1235), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n1181), .A2(new_n1209), .B1(new_n1234), .B2(new_n1231), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1236), .B(new_n743), .C1(KEYINPUT57), .C2(new_n1237), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n966), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n1154), .A2(new_n949), .B1(new_n964), .B2(new_n720), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1232), .A2(new_n1233), .B1(new_n1240), .B2(new_n963), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n794), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n795), .B1(new_n202), .B2(new_n874), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n829), .A2(G150), .ZN(new_n1244));
  INV_X1    g1044(.A(G132), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n1244), .B1(new_n819), .B2(new_n1201), .C1(new_n1245), .C2(new_n822), .ZN(new_n1246));
  INV_X1    g1046(.A(G125), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n1247), .A2(new_n888), .B1(new_n840), .B2(new_n991), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1246), .B(new_n1248), .C1(G128), .C2(new_n835), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  OR2_X1    g1050(.A1(new_n1250), .A2(KEYINPUT59), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(KEYINPUT59), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n261), .B(new_n303), .C1(new_n815), .C2(new_n263), .ZN(new_n1253));
  XOR2_X1   g1053(.A(KEYINPUT121), .B(G124), .Z(new_n1254));
  AOI21_X1  g1054(.A(new_n1253), .B1(new_n832), .B2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1251), .A2(new_n1252), .A3(new_n1255), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(G107), .A2(new_n835), .B1(new_n836), .B2(G116), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1257), .B1(new_n382), .B2(new_n840), .ZN(new_n1258));
  NOR4_X1   g1058(.A1(new_n1072), .A2(new_n988), .A3(new_n319), .A4(new_n301), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n814), .A2(G58), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n823), .A2(G97), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n1258), .B(new_n1262), .C1(G283), .C2(new_n832), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(KEYINPUT58), .ZN(new_n1264));
  OAI221_X1 g1064(.A(new_n358), .B1(G33), .B2(G41), .C1(new_n319), .C2(new_n301), .ZN(new_n1265));
  OR2_X1    g1065(.A1(new_n1263), .A2(KEYINPUT58), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1256), .A2(new_n1264), .A3(new_n1265), .A4(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1243), .B1(new_n1267), .B2(new_n807), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(new_n1227), .B2(new_n805), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1242), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1238), .A2(new_n1271), .ZN(G375));
  NAND2_X1  g1072(.A1(new_n1170), .A2(new_n1177), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n958), .A2(new_n804), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n795), .B1(G68), .B2(new_n874), .ZN(new_n1275));
  XOR2_X1   g1075(.A(new_n1275), .B(KEYINPUT122), .Z(new_n1276));
  OAI22_X1  g1076(.A1(new_n1245), .A2(new_n888), .B1(new_n844), .B2(new_n991), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(G150), .B2(new_n839), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n832), .A2(G128), .ZN(new_n1279));
  OAI221_X1 g1079(.A(new_n319), .B1(new_n819), .B2(new_n263), .C1(new_n822), .C2(new_n1201), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(G50), .B2(new_n829), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1278), .A2(new_n1260), .A3(new_n1279), .A4(new_n1281), .ZN(new_n1282));
  OAI22_X1  g1082(.A1(new_n816), .A2(new_n844), .B1(new_n888), .B2(new_n826), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1283), .B1(G107), .B2(new_n839), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n319), .B1(new_n814), .B2(G77), .ZN(new_n1285));
  XOR2_X1   g1085(.A(new_n1285), .B(KEYINPUT123), .Z(new_n1286));
  OAI221_X1 g1086(.A(new_n1071), .B1(new_n819), .B2(new_n535), .C1(new_n487), .C2(new_n822), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(G303), .B2(new_n832), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1284), .A2(new_n1286), .A3(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1282), .A2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1276), .B1(new_n1290), .B2(new_n807), .ZN(new_n1291));
  AOI22_X1  g1091(.A1(new_n1273), .A2(new_n794), .B1(new_n1274), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1179), .A2(new_n1048), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1273), .A2(new_n1209), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1292), .B1(new_n1293), .B2(new_n1294), .ZN(G381));
  XNOR2_X1  g1095(.A(G375), .B(KEYINPUT124), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1092), .A2(new_n860), .A3(new_n1093), .ZN(new_n1297));
  OR2_X1    g1097(.A1(G381), .A2(G384), .ZN(new_n1298));
  NOR4_X1   g1098(.A1(new_n1297), .A2(G390), .A3(new_n1298), .A4(G378), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1051), .A2(new_n1296), .A3(new_n1299), .ZN(G407));
  INV_X1    g1100(.A(G378), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1296), .A2(G213), .A3(new_n721), .A4(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(G407), .A2(G213), .A3(new_n1302), .ZN(G409));
  INV_X1    g1103(.A(new_n1050), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1093), .ZN(new_n1305));
  OAI21_X1  g1105(.A(G396), .B1(new_n1305), .B2(new_n1091), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1297), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT112), .ZN(new_n1308));
  AOI21_X1  g1108(.A(G390), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  AND2_X1   g1109(.A1(new_n1098), .A2(new_n1123), .ZN(new_n1310));
  AOI22_X1  g1110(.A1(new_n1297), .A2(new_n1306), .B1(new_n1310), .B2(new_n1100), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1304), .B1(new_n1309), .B2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1307), .A2(G390), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT112), .B1(new_n1306), .B2(new_n1297), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n1313), .B(new_n1050), .C1(G390), .C2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1312), .A2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n721), .A2(G213), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1179), .A2(new_n743), .ZN(new_n1318));
  NOR3_X1   g1118(.A1(new_n1273), .A2(KEYINPUT60), .A3(new_n1209), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(KEYINPUT60), .B1(new_n1273), .B2(new_n1209), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1318), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1292), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n898), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1321), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1325), .A2(new_n1319), .ZN(new_n1326));
  OAI211_X1 g1126(.A(G384), .B(new_n1292), .C1(new_n1326), .C2(new_n1318), .ZN(new_n1327));
  AND2_X1   g1127(.A1(new_n1324), .A2(new_n1327), .ZN(new_n1328));
  AND3_X1   g1128(.A1(new_n1238), .A2(G378), .A3(new_n1271), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1047), .B1(new_n1231), .B2(new_n1234), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1210), .A2(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1270), .B1(KEYINPUT125), .B2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT125), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1210), .A2(new_n1330), .A3(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(G378), .B1(new_n1332), .B2(new_n1334), .ZN(new_n1335));
  OAI211_X1 g1135(.A(new_n1317), .B(new_n1328), .C1(new_n1329), .C2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT62), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1238), .A2(G378), .A3(new_n1271), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1331), .A2(KEYINPUT125), .ZN(new_n1340));
  AND3_X1   g1140(.A1(new_n1340), .A2(new_n1271), .A3(new_n1334), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1339), .B1(new_n1341), .B2(G378), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1342), .A2(KEYINPUT62), .A3(new_n1317), .A4(new_n1328), .ZN(new_n1343));
  AND3_X1   g1143(.A1(new_n1338), .A2(KEYINPUT127), .A3(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT127), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1336), .A2(new_n1345), .A3(new_n1337), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1342), .A2(new_n1317), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1324), .A2(new_n1327), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n721), .A2(G213), .A3(G2897), .ZN(new_n1349));
  XNOR2_X1  g1149(.A(new_n1348), .B(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1347), .A2(new_n1350), .ZN(new_n1351));
  XNOR2_X1  g1151(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1346), .A2(new_n1351), .A3(new_n1352), .ZN(new_n1353));
  OAI21_X1  g1153(.A(new_n1316), .B1(new_n1344), .B2(new_n1353), .ZN(new_n1354));
  XNOR2_X1  g1154(.A(new_n1336), .B(KEYINPUT63), .ZN(new_n1355));
  AOI21_X1  g1155(.A(KEYINPUT61), .B1(new_n1347), .B2(new_n1350), .ZN(new_n1356));
  NAND4_X1  g1156(.A1(new_n1355), .A2(new_n1312), .A3(new_n1315), .A4(new_n1356), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1354), .A2(new_n1357), .ZN(G405));
  NAND2_X1  g1158(.A1(G375), .A2(new_n1301), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1359), .A2(new_n1339), .ZN(new_n1360));
  XNOR2_X1  g1160(.A(new_n1360), .B(new_n1328), .ZN(new_n1361));
  XNOR2_X1  g1161(.A(new_n1316), .B(new_n1361), .ZN(G402));
endmodule


