//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 0 1 0 1 1 0 1 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 1 0 1 0 1 0 1 0 1 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT30), .ZN(new_n188));
  XNOR2_X1  g002(.A(G143), .B(G146), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n189), .A2(KEYINPUT0), .A3(G128), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT0), .B(G128), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n189), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G137), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(KEYINPUT11), .A3(G134), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G137), .ZN(new_n196));
  AND2_X1   g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G131), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT11), .ZN(new_n199));
  OAI211_X1 g013(.A(KEYINPUT64), .B(new_n199), .C1(new_n195), .C2(G137), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n193), .A2(G134), .ZN(new_n202));
  AOI21_X1  g016(.A(KEYINPUT64), .B1(new_n202), .B2(new_n199), .ZN(new_n203));
  OAI211_X1 g017(.A(new_n197), .B(new_n198), .C1(new_n201), .C2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n199), .B1(new_n195), .B2(G137), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(new_n200), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n210), .A2(KEYINPUT65), .A3(new_n198), .A4(new_n197), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n206), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n197), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G131), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n192), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n198), .B1(new_n202), .B2(new_n196), .ZN(new_n216));
  INV_X1    g030(.A(G128), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n218));
  INV_X1    g032(.A(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G143), .ZN(new_n220));
  INV_X1    g034(.A(G143), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G146), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n218), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n221), .A2(KEYINPUT1), .A3(G146), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n223), .B(new_n224), .C1(G128), .C2(new_n189), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  AOI211_X1 g040(.A(new_n216), .B(new_n226), .C1(new_n206), .C2(new_n211), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n188), .B1(new_n215), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n225), .A2(KEYINPUT67), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n220), .A2(new_n222), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(new_n217), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n231), .A2(new_n232), .A3(new_n224), .A4(new_n223), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n216), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n212), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n206), .A2(new_n211), .B1(G131), .B2(new_n213), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n236), .B(KEYINPUT30), .C1(new_n237), .C2(new_n192), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT66), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT2), .ZN(new_n240));
  INV_X1    g054(.A(G113), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(KEYINPUT66), .A2(KEYINPUT2), .A3(G113), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n240), .A2(new_n241), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(G116), .B(G119), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n244), .A2(new_n245), .A3(new_n247), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n228), .A2(new_n238), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n215), .ZN(new_n253));
  INV_X1    g067(.A(new_n251), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n254), .A3(new_n236), .ZN(new_n255));
  NOR2_X1   g069(.A1(G237), .A2(G953), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G210), .ZN(new_n257));
  XOR2_X1   g071(.A(new_n257), .B(KEYINPUT27), .Z(new_n258));
  XNOR2_X1  g072(.A(new_n258), .B(KEYINPUT26), .ZN(new_n259));
  INV_X1    g073(.A(G101), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n259), .B(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n252), .A2(new_n255), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT68), .ZN(new_n263));
  AND3_X1   g077(.A1(new_n262), .A2(new_n263), .A3(KEYINPUT31), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT28), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n236), .B1(new_n237), .B2(new_n192), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n265), .B1(new_n266), .B2(new_n251), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n251), .B1(new_n215), .B2(new_n227), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n253), .A2(KEYINPUT28), .A3(new_n254), .A4(new_n236), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n261), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT31), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n252), .A2(new_n273), .A3(new_n255), .A4(new_n261), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n263), .B1(new_n262), .B2(KEYINPUT31), .ZN(new_n276));
  NOR3_X1   g090(.A1(new_n264), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(G472), .A2(G902), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n187), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n275), .ZN(new_n281));
  INV_X1    g095(.A(new_n276), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n262), .A2(new_n263), .A3(KEYINPUT31), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(KEYINPUT32), .A3(new_n278), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n266), .A2(new_n251), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(new_n255), .A3(KEYINPUT69), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT69), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n266), .A2(new_n288), .A3(new_n251), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n267), .B1(new_n290), .B2(new_n265), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT29), .ZN(new_n292));
  NOR3_X1   g106(.A1(new_n291), .A2(new_n292), .A3(new_n271), .ZN(new_n293));
  INV_X1    g107(.A(G902), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n292), .B1(new_n270), .B2(new_n271), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n261), .B1(new_n252), .B2(new_n255), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(G472), .B1(new_n293), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n280), .A2(new_n285), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G119), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n300), .A2(G128), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n301), .B1(KEYINPUT70), .B2(KEYINPUT23), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n217), .A2(G119), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT23), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT70), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n306), .B1(new_n300), .B2(G128), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n302), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n301), .A2(new_n303), .ZN(new_n309));
  XOR2_X1   g123(.A(KEYINPUT24), .B(G110), .Z(new_n310));
  OAI22_X1  g124(.A1(new_n308), .A2(G110), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(G125), .B(G140), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT16), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT71), .ZN(new_n314));
  INV_X1    g128(.A(G140), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G125), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n314), .B1(new_n316), .B2(KEYINPUT16), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT16), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n318), .A2(new_n315), .A3(KEYINPUT71), .A4(G125), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n313), .A2(new_n317), .A3(G146), .A4(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n312), .A2(new_n219), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n311), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n322), .B(KEYINPUT72), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n309), .A2(new_n310), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n308), .A2(G110), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n313), .A2(new_n317), .A3(new_n319), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n219), .ZN(new_n327));
  AOI211_X1 g141(.A(new_n324), .B(new_n325), .C1(new_n320), .C2(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G953), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(G221), .A3(G234), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(KEYINPUT22), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n332), .B(G137), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n333), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n335), .B1(new_n323), .B2(new_n328), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n334), .A2(new_n294), .A3(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT25), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT73), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n337), .B(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G217), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n342), .B1(G234), .B2(new_n294), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n334), .A2(new_n336), .ZN(new_n346));
  NOR3_X1   g160(.A1(new_n346), .A2(G902), .A3(new_n343), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n299), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT74), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT74), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n299), .A2(new_n348), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(G110), .B(G140), .ZN(new_n354));
  INV_X1    g168(.A(G227), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n355), .A2(G953), .ZN(new_n356));
  XOR2_X1   g170(.A(new_n354), .B(new_n356), .Z(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT78), .ZN(new_n359));
  INV_X1    g173(.A(G104), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT3), .B1(new_n360), .B2(G107), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT3), .ZN(new_n362));
  INV_X1    g176(.A(G107), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(new_n363), .A3(G104), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n360), .A2(G107), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n361), .A2(new_n364), .A3(new_n260), .A4(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n363), .A2(G104), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n360), .A2(G107), .ZN(new_n368));
  OAI21_X1  g182(.A(G101), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(KEYINPUT76), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n363), .A2(G104), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n365), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(KEYINPUT76), .B1(new_n373), .B2(G101), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n371), .A2(new_n225), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT77), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n374), .B1(new_n370), .B2(KEYINPUT76), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT77), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(new_n225), .ZN(new_n380));
  AOI21_X1  g194(.A(KEYINPUT10), .B1(new_n377), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n234), .A2(KEYINPUT10), .A3(new_n378), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n361), .A2(new_n364), .A3(new_n365), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT4), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(G101), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(KEYINPUT75), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT75), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n383), .A2(new_n387), .A3(new_n384), .A4(G101), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n192), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n384), .B1(new_n383), .B2(G101), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n366), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n389), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n382), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n359), .B1(new_n381), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT10), .ZN(new_n396));
  AND4_X1   g210(.A1(new_n379), .A2(new_n371), .A3(new_n225), .A4(new_n375), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n379), .B1(new_n378), .B2(new_n225), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n386), .A2(new_n388), .B1(new_n366), .B2(new_n391), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n396), .B1(new_n229), .B2(new_n233), .ZN(new_n401));
  AOI22_X1  g215(.A1(new_n390), .A2(new_n400), .B1(new_n401), .B2(new_n378), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n399), .A2(new_n402), .A3(KEYINPUT78), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n237), .B1(new_n395), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n399), .A2(new_n402), .A3(new_n237), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n358), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n357), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT12), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n378), .A2(new_n225), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n411), .B1(new_n377), .B2(new_n380), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n410), .B1(new_n412), .B2(new_n237), .ZN(new_n413));
  INV_X1    g227(.A(new_n378), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n226), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n415), .B1(new_n397), .B2(new_n398), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n212), .A2(new_n214), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n416), .A2(KEYINPUT12), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n413), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n409), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n407), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G469), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n421), .A2(new_n422), .A3(new_n294), .ZN(new_n423));
  NAND2_X1  g237(.A1(G469), .A2(G902), .ZN(new_n424));
  NOR3_X1   g238(.A1(new_n381), .A2(new_n394), .A3(new_n359), .ZN(new_n425));
  AOI21_X1  g239(.A(KEYINPUT78), .B1(new_n399), .B2(new_n402), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n417), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NOR3_X1   g241(.A1(new_n412), .A2(new_n410), .A3(new_n237), .ZN(new_n428));
  AOI21_X1  g242(.A(KEYINPUT12), .B1(new_n416), .B2(new_n417), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n405), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n427), .A2(new_n409), .B1(new_n430), .B2(new_n358), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(G469), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n423), .A2(new_n424), .A3(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT9), .B(G234), .ZN(new_n434));
  OAI21_X1  g248(.A(G221), .B1(new_n434), .B2(G902), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G475), .ZN(new_n437));
  XNOR2_X1  g251(.A(G113), .B(G122), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n438), .B(new_n360), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT85), .ZN(new_n440));
  AOI21_X1  g254(.A(KEYINPUT19), .B1(new_n312), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G125), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G140), .ZN(new_n443));
  AND4_X1   g257(.A1(new_n440), .A2(new_n316), .A3(new_n443), .A4(KEYINPUT19), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n219), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT86), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n256), .A2(G143), .A3(G214), .ZN(new_n447));
  AOI21_X1  g261(.A(G143), .B1(new_n256), .B2(G214), .ZN(new_n448));
  OAI21_X1  g262(.A(G131), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G237), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(new_n330), .A3(G214), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n221), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n256), .A2(G143), .A3(G214), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n198), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT86), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n456), .B(new_n219), .C1(new_n441), .C2(new_n444), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n446), .A2(new_n320), .A3(new_n455), .A4(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n312), .B(new_n219), .ZN(new_n459));
  AND2_X1   g273(.A1(KEYINPUT18), .A2(G131), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n447), .A2(new_n448), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n460), .B1(new_n461), .B2(KEYINPUT84), .ZN(new_n462));
  AND4_X1   g276(.A1(KEYINPUT84), .A2(new_n452), .A3(new_n460), .A4(new_n453), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n439), .B1(new_n458), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT17), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n449), .A2(new_n466), .A3(new_n454), .ZN(new_n467));
  OAI211_X1 g281(.A(KEYINPUT17), .B(G131), .C1(new_n447), .C2(new_n448), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n327), .A2(new_n467), .A3(new_n320), .A4(new_n468), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n469), .A2(new_n464), .A3(new_n439), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n437), .B(new_n294), .C1(new_n465), .C2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT20), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n316), .A2(new_n443), .A3(new_n440), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT19), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n312), .A2(new_n440), .A3(KEYINPUT19), .ZN(new_n476));
  AOI21_X1  g290(.A(G146), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n320), .B(new_n455), .C1(new_n477), .C2(new_n456), .ZN(new_n478));
  INV_X1    g292(.A(new_n457), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n464), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n439), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n469), .A2(new_n464), .A3(new_n439), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT20), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n484), .A2(new_n485), .A3(new_n437), .A4(new_n294), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n472), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n439), .B1(new_n469), .B2(new_n464), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n294), .B1(new_n470), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT87), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT87), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n491), .B(new_n294), .C1(new_n470), .C2(new_n488), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n490), .A2(G475), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT90), .ZN(new_n495));
  INV_X1    g309(.A(G478), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n496), .A2(KEYINPUT15), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n221), .A2(G128), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n217), .A2(G143), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n195), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n499), .A2(new_n500), .A3(G134), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT13), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n500), .A2(new_n504), .A3(G134), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n502), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n499), .A2(new_n500), .A3(new_n504), .A4(G134), .ZN(new_n507));
  INV_X1    g321(.A(G116), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n508), .A2(G122), .ZN(new_n509));
  INV_X1    g323(.A(G122), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n510), .A2(G116), .ZN(new_n511));
  OAI21_X1  g325(.A(G107), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(G116), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n508), .A2(G122), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n514), .A3(new_n363), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n512), .A2(KEYINPUT88), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(KEYINPUT88), .B1(new_n512), .B2(new_n515), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n506), .B(new_n507), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n515), .B(KEYINPUT89), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n502), .A2(new_n503), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT14), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n513), .B1(new_n511), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n514), .A2(KEYINPUT14), .ZN(new_n523));
  OAI21_X1  g337(.A(G107), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n519), .A2(new_n520), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n518), .A2(new_n525), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n434), .A2(new_n342), .A3(G953), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n518), .A2(new_n525), .A3(new_n527), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n498), .B1(new_n531), .B2(new_n294), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n518), .A2(new_n527), .A3(new_n525), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n527), .B1(new_n518), .B2(new_n525), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n294), .B(new_n498), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n495), .B1(new_n532), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n294), .B1(new_n533), .B2(new_n534), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n497), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(new_n535), .A3(KEYINPUT90), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n330), .A2(G952), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n542), .B1(G234), .B2(G237), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  XOR2_X1   g358(.A(KEYINPUT21), .B(G898), .Z(new_n545));
  NAND2_X1  g359(.A1(G234), .A2(G237), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(G902), .A3(G953), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n544), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n494), .A2(new_n541), .A3(new_n549), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n436), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(G214), .B1(G237), .B2(G902), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n389), .A2(new_n251), .A3(new_n392), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n508), .A2(KEYINPUT5), .A3(G119), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n554), .B1(new_n247), .B2(KEYINPUT5), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(G113), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n378), .A2(new_n250), .A3(new_n556), .ZN(new_n557));
  XOR2_X1   g371(.A(G110), .B(G122), .Z(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n553), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n559), .B1(new_n553), .B2(new_n557), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT6), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n553), .A2(new_n557), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n558), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n565), .A2(KEYINPUT6), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT79), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n226), .A2(new_n442), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(KEYINPUT80), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n192), .A2(G125), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(G224), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(G953), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n571), .B(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n553), .A2(new_n557), .A3(new_n559), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n565), .A2(KEYINPUT6), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT79), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n567), .A2(new_n574), .A3(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(KEYINPUT7), .B1(new_n572), .B2(G953), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n569), .A2(KEYINPUT81), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n570), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n569), .A2(KEYINPUT81), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n580), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n556), .A2(new_n250), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n414), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n557), .ZN(new_n587));
  XOR2_X1   g401(.A(new_n558), .B(KEYINPUT8), .Z(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n571), .ZN(new_n590));
  INV_X1    g404(.A(new_n580), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n560), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n584), .A2(new_n589), .A3(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n579), .A2(new_n294), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT82), .ZN(new_n595));
  OAI21_X1  g409(.A(G210), .B1(G237), .B2(G902), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT82), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n579), .A2(new_n598), .A3(new_n593), .A4(new_n294), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n595), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT83), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n579), .A2(new_n294), .A3(new_n593), .A4(new_n596), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n595), .A2(KEYINPUT83), .A3(new_n597), .A4(new_n599), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n551), .A2(new_n552), .A3(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n353), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(new_n260), .ZN(G3));
  NOR2_X1   g422(.A1(new_n264), .A2(new_n276), .ZN(new_n609));
  AOI21_X1  g423(.A(G902), .B1(new_n609), .B2(new_n281), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT91), .ZN(new_n611));
  INV_X1    g425(.A(G472), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n284), .A2(new_n294), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n614), .A2(KEYINPUT91), .A3(G472), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n348), .A2(new_n436), .A3(new_n613), .A4(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT92), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n533), .A2(new_n534), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n618), .A2(KEYINPUT93), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT93), .ZN(new_n621));
  AOI21_X1  g435(.A(KEYINPUT33), .B1(new_n531), .B2(new_n621), .ZN(new_n622));
  OAI211_X1 g436(.A(G478), .B(new_n294), .C1(new_n620), .C2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n538), .A2(new_n496), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n494), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n594), .A2(new_n597), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n603), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n628), .A2(new_n552), .A3(new_n548), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n617), .A2(new_n626), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT34), .B(G104), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  NAND3_X1  g446(.A1(new_n472), .A2(new_n486), .A3(KEYINPUT94), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT94), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n471), .A2(new_n634), .A3(KEYINPUT20), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n539), .A2(KEYINPUT90), .A3(new_n535), .ZN(new_n637));
  AOI21_X1  g451(.A(KEYINPUT90), .B1(new_n539), .B2(new_n535), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n640), .A2(KEYINPUT95), .A3(new_n548), .A4(new_n493), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT95), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n541), .A2(new_n493), .A3(new_n635), .A4(new_n633), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n642), .B1(new_n643), .B2(new_n549), .ZN(new_n644));
  AND4_X1   g458(.A1(new_n552), .A2(new_n628), .A3(new_n641), .A4(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n617), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G107), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT96), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT35), .ZN(G9));
  AND2_X1   g464(.A1(new_n615), .A2(new_n613), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n335), .A2(KEYINPUT36), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n329), .B(new_n652), .ZN(new_n653));
  OAI211_X1 g467(.A(new_n653), .B(new_n294), .C1(new_n342), .C2(G234), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT97), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n344), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n606), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT37), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G110), .ZN(G12));
  AND3_X1   g474(.A1(new_n299), .A2(new_n436), .A3(new_n656), .ZN(new_n661));
  INV_X1    g475(.A(new_n552), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n662), .B1(new_n627), .B2(new_n603), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n544), .B1(new_n547), .B2(G900), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n643), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n663), .A2(KEYINPUT98), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n663), .A2(new_n666), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT98), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n661), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G128), .ZN(G30));
  XNOR2_X1  g486(.A(new_n664), .B(KEYINPUT39), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n436), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n674), .A2(KEYINPUT40), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(new_n656), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n494), .A2(new_n541), .ZN(new_n677));
  AOI211_X1 g491(.A(new_n662), .B(new_n677), .C1(new_n674), .C2(KEYINPUT40), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT99), .B(KEYINPUT100), .ZN(new_n679));
  XOR2_X1   g493(.A(new_n679), .B(KEYINPUT38), .Z(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n605), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n602), .A2(new_n603), .A3(new_n604), .A4(new_n680), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n280), .A2(new_n285), .ZN(new_n685));
  AOI21_X1  g499(.A(G902), .B1(new_n290), .B2(new_n271), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n252), .A2(new_n255), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n261), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n612), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  OR2_X1    g503(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n676), .A2(new_n678), .A3(new_n684), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G143), .ZN(G45));
  NOR2_X1   g506(.A1(new_n626), .A2(new_n665), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n661), .A2(new_n663), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  AOI21_X1  g509(.A(new_n357), .B1(new_n427), .B2(new_n405), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n408), .B1(new_n418), .B2(new_n413), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n294), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(G469), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n699), .A2(new_n435), .A3(new_n423), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT101), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n699), .A2(KEYINPUT101), .A3(new_n435), .A4(new_n423), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n626), .ZN(new_n705));
  AND3_X1   g519(.A1(new_n663), .A2(new_n548), .A3(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n704), .A2(new_n706), .A3(new_n299), .A4(new_n348), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT41), .B(G113), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G15));
  NAND4_X1  g523(.A1(new_n704), .A2(new_n645), .A3(new_n299), .A4(new_n348), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT102), .B(G116), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G18));
  NAND2_X1  g526(.A1(new_n628), .A2(new_n552), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n700), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n714), .A2(new_n299), .A3(new_n550), .A4(new_n656), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G119), .ZN(G21));
  AOI21_X1  g530(.A(new_n629), .B1(new_n702), .B2(new_n703), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n291), .A2(new_n271), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n262), .B(new_n273), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n279), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g534(.A(KEYINPUT103), .B1(new_n610), .B2(new_n612), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT103), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n614), .A2(new_n722), .A3(G472), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n720), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n677), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n717), .A2(new_n724), .A3(new_n348), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(KEYINPUT104), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G122), .ZN(G24));
  NAND4_X1  g542(.A1(new_n724), .A2(new_n656), .A3(new_n693), .A4(new_n714), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G125), .ZN(G27));
  NAND4_X1  g544(.A1(new_n602), .A2(new_n552), .A3(new_n603), .A4(new_n604), .ZN(new_n731));
  INV_X1    g545(.A(new_n435), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n423), .A2(new_n432), .ZN(new_n733));
  XOR2_X1   g547(.A(new_n424), .B(KEYINPUT105), .Z(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n732), .B1(new_n733), .B2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n731), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n685), .A2(KEYINPUT106), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT106), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n285), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n739), .A2(new_n298), .A3(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n738), .A2(new_n742), .A3(new_n348), .A4(new_n693), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(KEYINPUT42), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT42), .ZN(new_n745));
  INV_X1    g559(.A(new_n349), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n738), .A2(new_n745), .A3(new_n746), .A4(new_n693), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(new_n198), .ZN(G33));
  OR3_X1    g563(.A1(new_n643), .A2(KEYINPUT107), .A3(new_n665), .ZN(new_n750));
  OAI21_X1  g564(.A(KEYINPUT107), .B1(new_n643), .B2(new_n665), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n738), .A2(new_n746), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G134), .ZN(G36));
  NAND2_X1  g567(.A1(new_n427), .A2(new_n409), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n430), .A2(new_n358), .ZN(new_n755));
  AOI21_X1  g569(.A(KEYINPUT45), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(KEYINPUT108), .B1(new_n756), .B2(new_n422), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT108), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n758), .B(G469), .C1(new_n431), .C2(KEYINPUT45), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n431), .A2(KEYINPUT45), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n757), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(KEYINPUT46), .A3(new_n735), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n423), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT109), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(KEYINPUT46), .B1(new_n761), .B2(new_n735), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n762), .A2(KEYINPUT109), .A3(new_n423), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n765), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n769), .A2(new_n435), .A3(new_n673), .ZN(new_n770));
  XOR2_X1   g584(.A(new_n770), .B(KEYINPUT110), .Z(new_n771));
  OR2_X1    g585(.A1(new_n494), .A2(KEYINPUT111), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT43), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n625), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n775), .A2(new_n494), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n772), .B(new_n773), .C1(new_n494), .C2(new_n775), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n651), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n656), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n731), .B1(new_n783), .B2(KEYINPUT44), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n771), .B(new_n784), .C1(KEYINPUT44), .C2(new_n783), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G137), .ZN(G39));
  XNOR2_X1  g600(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n769), .A2(new_n435), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n787), .B1(new_n769), .B2(new_n435), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n731), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n299), .A2(new_n348), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n790), .A2(new_n693), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G140), .ZN(G42));
  NAND2_X1  g608(.A1(new_n721), .A2(new_n723), .ZN(new_n795));
  INV_X1    g609(.A(new_n720), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n795), .A2(new_n348), .A3(new_n725), .A4(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n629), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n704), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n707), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT113), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n532), .A2(new_n536), .ZN(new_n802));
  OR3_X1    g616(.A1(new_n494), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n801), .B1(new_n494), .B2(new_n802), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n803), .A2(new_n626), .A3(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n549), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n605), .A2(new_n807), .A3(new_n552), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n616), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n710), .A2(new_n715), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n800), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n724), .A2(new_n656), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n812), .A2(new_n693), .A3(new_n738), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n814));
  INV_X1    g628(.A(new_n636), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n493), .A2(new_n802), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n815), .A2(new_n664), .A3(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n814), .A2(KEYINPUT114), .A3(new_n552), .A4(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT114), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n820), .B1(new_n731), .B2(new_n817), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n819), .A2(new_n661), .A3(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n606), .ZN(new_n823));
  INV_X1    g637(.A(new_n352), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n351), .B1(new_n299), .B2(new_n348), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n657), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n823), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n811), .A2(new_n813), .A3(new_n822), .A4(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n744), .A2(new_n747), .A3(new_n752), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT115), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n656), .A2(new_n665), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n713), .A2(new_n677), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n690), .A2(new_n736), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n671), .A2(new_n694), .A3(new_n834), .A4(new_n729), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n835), .B(new_n836), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n744), .A2(new_n747), .A3(new_n752), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n606), .B1(new_n353), .B2(new_n657), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n726), .A2(new_n707), .A3(new_n710), .A4(new_n715), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n839), .A2(new_n840), .A3(new_n809), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT115), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n822), .A2(new_n813), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n838), .A2(new_n841), .A3(new_n842), .A4(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n831), .A2(new_n837), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n809), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n710), .A2(new_n715), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n849), .A2(new_n850), .A3(new_n707), .A4(new_n726), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n851), .A2(new_n843), .A3(new_n839), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n837), .A2(new_n852), .A3(KEYINPUT53), .A4(new_n838), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT116), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n829), .A2(new_n830), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT116), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n855), .A2(new_n856), .A3(KEYINPUT53), .A4(new_n837), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(KEYINPUT54), .B1(new_n848), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT117), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n699), .A2(new_n423), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n861), .A2(new_n435), .ZN(new_n862));
  INV_X1    g676(.A(new_n787), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n762), .A2(KEYINPUT109), .A3(new_n423), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT109), .B1(new_n762), .B2(new_n423), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n864), .A2(new_n865), .A3(new_n766), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n863), .B1(new_n866), .B2(new_n732), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n769), .A2(new_n435), .A3(new_n787), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n862), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n544), .B1(new_n777), .B2(new_n778), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n724), .A2(new_n348), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(new_n791), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n860), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n348), .A2(new_n543), .ZN(new_n874));
  NOR4_X1   g688(.A1(new_n690), .A2(new_n731), .A3(new_n874), .A4(new_n700), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n625), .A2(new_n494), .ZN(new_n876));
  NOR4_X1   g690(.A1(new_n731), .A2(new_n780), .A3(new_n544), .A4(new_n700), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n875), .A2(new_n876), .B1(new_n877), .B2(new_n812), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT118), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n682), .A2(new_n662), .A3(new_n683), .ZN(new_n881));
  INV_X1    g695(.A(new_n700), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n724), .A2(new_n348), .A3(new_n882), .A4(new_n870), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT50), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n682), .A2(new_n662), .A3(new_n683), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT50), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n886), .A2(new_n883), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n880), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n881), .A2(new_n884), .A3(KEYINPUT50), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n887), .B1(new_n886), .B2(new_n883), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n890), .A2(KEYINPUT118), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n879), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n862), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n894), .B1(new_n788), .B2(new_n789), .ZN(new_n895));
  INV_X1    g709(.A(new_n872), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n895), .A2(KEYINPUT117), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n873), .A2(new_n893), .A3(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT51), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n899), .B1(new_n890), .B2(new_n891), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n878), .B(new_n901), .C1(new_n869), .C2(new_n872), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n871), .A2(new_n714), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n742), .A2(new_n348), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT119), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n905), .A2(new_n877), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n791), .A2(new_n882), .A3(new_n870), .ZN(new_n908));
  OAI21_X1  g722(.A(KEYINPUT119), .B1(new_n908), .B2(new_n904), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n907), .A2(new_n909), .A3(KEYINPUT48), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n542), .B1(new_n875), .B2(new_n705), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n911), .B1(KEYINPUT48), .B2(new_n909), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n902), .A2(new_n903), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n900), .A2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT120), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n838), .A2(new_n841), .A3(new_n844), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n835), .B(KEYINPUT52), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n847), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n853), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n921), .A2(KEYINPUT54), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n900), .A2(KEYINPUT120), .A3(new_n914), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n859), .A2(new_n917), .A3(new_n923), .A4(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(G952), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n330), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n345), .A2(new_n347), .A3(new_n662), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n861), .A2(KEYINPUT49), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n861), .A2(KEYINPUT49), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n932), .A2(new_n690), .A3(new_n732), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n933), .A2(new_n683), .A3(new_n682), .A4(new_n776), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n928), .A2(new_n934), .ZN(G75));
  AOI21_X1  g749(.A(new_n294), .B1(new_n920), .B2(new_n853), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT56), .B1(new_n936), .B2(G210), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n567), .A2(new_n578), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(new_n574), .Z(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT55), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(KEYINPUT121), .B1(new_n937), .B2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT121), .ZN(new_n943));
  INV_X1    g757(.A(G210), .ZN(new_n944));
  AOI211_X1 g758(.A(new_n944), .B(new_n294), .C1(new_n920), .C2(new_n853), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n943), .B(new_n940), .C1(new_n945), .C2(KEYINPUT56), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n942), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n926), .A2(G953), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT123), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT56), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n945), .B2(KEYINPUT122), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n921), .A2(KEYINPUT122), .A3(G210), .A4(G902), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n941), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n949), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n947), .A2(new_n954), .ZN(G51));
  INV_X1    g769(.A(new_n949), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n735), .A2(KEYINPUT57), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n735), .A2(KEYINPUT57), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT54), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n959), .B1(new_n920), .B2(new_n853), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n957), .B(new_n958), .C1(new_n922), .C2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n421), .ZN(new_n962));
  INV_X1    g776(.A(new_n761), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n936), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n956), .B1(new_n962), .B2(new_n964), .ZN(G54));
  NAND3_X1  g779(.A1(new_n936), .A2(KEYINPUT58), .A3(G475), .ZN(new_n966));
  OR2_X1    g780(.A1(new_n966), .A2(new_n484), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n484), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n956), .B1(new_n967), .B2(new_n968), .ZN(G60));
  NOR2_X1   g783(.A1(new_n620), .A2(new_n622), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(G478), .A2(G902), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT59), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n971), .B(new_n973), .C1(new_n922), .C2(new_n960), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n949), .ZN(new_n975));
  INV_X1    g789(.A(new_n858), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n846), .A2(new_n847), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n959), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n973), .B1(new_n978), .B2(new_n922), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n975), .B1(new_n979), .B2(new_n970), .ZN(G63));
  NAND2_X1  g794(.A1(G217), .A2(G902), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT60), .Z(new_n982));
  AND2_X1   g796(.A1(new_n921), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n956), .B1(new_n983), .B2(new_n653), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n346), .B(KEYINPUT124), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n984), .B(KEYINPUT61), .C1(new_n983), .C2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT61), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n983), .A2(new_n985), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n921), .A2(new_n982), .ZN(new_n989));
  INV_X1    g803(.A(new_n653), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n949), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n987), .B1(new_n988), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n986), .A2(new_n992), .ZN(G66));
  AOI21_X1  g807(.A(new_n330), .B1(new_n545), .B2(G224), .ZN(new_n994));
  INV_X1    g808(.A(new_n841), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n994), .B1(new_n995), .B2(new_n330), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n938), .B1(G898), .B2(new_n330), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT125), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n996), .B(new_n998), .ZN(G69));
  AND3_X1   g813(.A1(new_n671), .A2(new_n694), .A3(new_n729), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n793), .A2(new_n1000), .A3(new_n838), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n771), .A2(new_n905), .A3(new_n833), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n1001), .A2(new_n785), .A3(new_n330), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n228), .A2(new_n238), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n441), .A2(new_n444), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  AND2_X1   g820(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(G900), .ZN(new_n1008));
  OAI21_X1  g822(.A(G953), .B1(new_n1008), .B2(G227), .ZN(new_n1009));
  OR4_X1    g823(.A1(new_n353), .A2(new_n674), .A3(new_n731), .A4(new_n806), .ZN(new_n1010));
  NAND2_X1  g824(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1000), .A2(new_n691), .A3(new_n1011), .ZN(new_n1012));
  NOR2_X1   g826(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n785), .A2(new_n793), .A3(new_n1010), .A4(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1006), .B1(new_n1015), .B2(new_n330), .ZN(new_n1016));
  OAI21_X1  g830(.A(G953), .B1(new_n355), .B2(new_n1008), .ZN(new_n1017));
  AOI22_X1  g831(.A1(new_n1007), .A2(new_n1009), .B1(new_n1016), .B2(new_n1017), .ZN(G72));
  NAND2_X1  g832(.A1(G472), .A2(G902), .ZN(new_n1019));
  XOR2_X1   g833(.A(new_n1019), .B(KEYINPUT63), .Z(new_n1020));
  XNOR2_X1  g834(.A(new_n1020), .B(KEYINPUT127), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1001), .A2(new_n785), .A3(new_n1002), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n1021), .B1(new_n1022), .B2(new_n995), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n687), .A2(new_n261), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n956), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1021), .B1(new_n1015), .B2(new_n995), .ZN(new_n1026));
  INV_X1    g840(.A(new_n688), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n1027), .A2(new_n1024), .ZN(new_n1029));
  OAI211_X1 g843(.A(new_n1020), .B(new_n1029), .C1(new_n848), .C2(new_n858), .ZN(new_n1030));
  AND3_X1   g844(.A1(new_n1025), .A2(new_n1028), .A3(new_n1030), .ZN(G57));
endmodule


