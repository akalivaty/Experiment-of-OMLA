

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726;

  XNOR2_X1 U365 ( .A(n694), .B(n695), .ZN(n345) );
  BUF_X1 U366 ( .A(n682), .Z(n693) );
  AND2_X1 U367 ( .A1(n599), .A2(n632), .ZN(n714) );
  NOR2_X1 U368 ( .A1(n532), .A2(n533), .ZN(n623) );
  AND2_X1 U369 ( .A1(n403), .A2(n564), .ZN(n587) );
  BUF_X1 U370 ( .A(G143), .Z(n343) );
  NOR2_X1 U371 ( .A1(G953), .A2(G237), .ZN(n499) );
  XNOR2_X1 U372 ( .A(G104), .B(G107), .ZN(n470) );
  NOR2_X1 U373 ( .A1(n610), .A2(n344), .ZN(n594) );
  NAND2_X1 U374 ( .A1(n591), .A2(n592), .ZN(n344) );
  XNOR2_X2 U375 ( .A(n469), .B(n468), .ZN(n712) );
  XNOR2_X2 U376 ( .A(n430), .B(n570), .ZN(n665) );
  XNOR2_X2 U377 ( .A(n432), .B(n431), .ZN(n540) );
  XNOR2_X2 U378 ( .A(n540), .B(n356), .ZN(n558) );
  NOR2_X1 U379 ( .A1(n345), .A2(n697), .ZN(G66) );
  XOR2_X1 U380 ( .A(KEYINPUT98), .B(n343), .Z(n498) );
  INV_X1 U381 ( .A(n623), .ZN(n625) );
  XNOR2_X2 U382 ( .A(n360), .B(n357), .ZN(n723) );
  AND2_X2 U383 ( .A1(n562), .A2(n561), .ZN(n360) );
  XNOR2_X2 U384 ( .A(n480), .B(n479), .ZN(n536) );
  INV_X1 U385 ( .A(n581), .ZN(n417) );
  XNOR2_X1 U386 ( .A(n492), .B(n491), .ZN(n365) );
  NOR2_X1 U387 ( .A1(n417), .A2(n584), .ZN(n610) );
  XNOR2_X1 U388 ( .A(n673), .B(n436), .ZN(n674) );
  XNOR2_X1 U389 ( .A(n700), .B(n494), .ZN(n673) );
  XNOR2_X1 U390 ( .A(n365), .B(n503), .ZN(n361) );
  XOR2_X1 U391 ( .A(G110), .B(KEYINPUT16), .Z(n492) );
  INV_X2 U392 ( .A(G143), .ZN(n426) );
  XNOR2_X1 U393 ( .A(n482), .B(KEYINPUT96), .ZN(n585) );
  XOR2_X1 U394 ( .A(KEYINPUT42), .B(n524), .Z(n725) );
  XNOR2_X1 U395 ( .A(n361), .B(n493), .ZN(n700) );
  XNOR2_X1 U396 ( .A(n412), .B(KEYINPUT0), .ZN(n346) );
  INV_X1 U397 ( .A(n549), .ZN(n347) );
  XNOR2_X1 U398 ( .A(n412), .B(KEYINPUT0), .ZN(n571) );
  NOR2_X1 U399 ( .A1(n531), .A2(n558), .ZN(n622) );
  XNOR2_X2 U400 ( .A(n509), .B(n354), .ZN(n469) );
  XNOR2_X2 U401 ( .A(n487), .B(G134), .ZN(n509) );
  XNOR2_X1 U402 ( .A(n534), .B(KEYINPUT104), .ZN(n655) );
  XNOR2_X1 U403 ( .A(G137), .B(KEYINPUT71), .ZN(n468) );
  XNOR2_X1 U404 ( .A(n385), .B(n351), .ZN(n527) );
  OR2_X1 U405 ( .A1(n684), .A2(G902), .ZN(n385) );
  INV_X1 U406 ( .A(KEYINPUT64), .ZN(n411) );
  XNOR2_X1 U407 ( .A(n421), .B(n370), .ZN(n369) );
  INV_X1 U408 ( .A(KEYINPUT47), .ZN(n370) );
  INV_X1 U409 ( .A(n621), .ZN(n368) );
  NAND2_X1 U410 ( .A1(n423), .A2(n422), .ZN(n364) );
  INV_X1 U411 ( .A(G900), .ZN(n422) );
  XNOR2_X1 U412 ( .A(n424), .B(KEYINPUT106), .ZN(n423) );
  NOR2_X1 U413 ( .A1(n554), .A2(n715), .ZN(n424) );
  XNOR2_X1 U414 ( .A(n467), .B(KEYINPUT21), .ZN(n637) );
  XNOR2_X1 U415 ( .A(n486), .B(n485), .ZN(n490) );
  XNOR2_X1 U416 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n485) );
  XOR2_X1 U417 ( .A(KEYINPUT18), .B(KEYINPUT87), .Z(n486) );
  XNOR2_X1 U418 ( .A(G902), .B(KEYINPUT15), .ZN(n603) );
  OR2_X1 U419 ( .A1(G237), .A2(G902), .ZN(n495) );
  XNOR2_X1 U420 ( .A(n371), .B(G472), .ZN(n537) );
  OR2_X1 U421 ( .A1(n604), .A2(G902), .ZN(n371) );
  XOR2_X1 U422 ( .A(n537), .B(KEYINPUT6), .Z(n569) );
  XNOR2_X1 U423 ( .A(KEYINPUT3), .B(G119), .ZN(n443) );
  XNOR2_X1 U424 ( .A(n434), .B(n468), .ZN(n366) );
  XOR2_X1 U425 ( .A(G119), .B(G110), .Z(n434) );
  XNOR2_X1 U426 ( .A(G128), .B(KEYINPUT24), .ZN(n458) );
  XNOR2_X1 U427 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n510) );
  XNOR2_X1 U428 ( .A(G122), .B(KEYINPUT102), .ZN(n507) );
  XOR2_X1 U429 ( .A(KEYINPUT100), .B(KEYINPUT103), .Z(n508) );
  XNOR2_X1 U430 ( .A(G113), .B(G131), .ZN(n497) );
  XOR2_X1 U431 ( .A(KEYINPUT70), .B(KEYINPUT10), .Z(n457) );
  XNOR2_X1 U432 ( .A(n349), .B(G140), .ZN(n401) );
  XOR2_X1 U433 ( .A(G122), .B(G104), .Z(n503) );
  XOR2_X1 U434 ( .A(KEYINPUT12), .B(KEYINPUT97), .Z(n501) );
  XNOR2_X1 U435 ( .A(n712), .B(n478), .ZN(n677) );
  XNOR2_X1 U436 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U437 ( .A(n382), .B(n381), .ZN(n663) );
  INV_X1 U438 ( .A(KEYINPUT52), .ZN(n381) );
  BUF_X1 U439 ( .A(n564), .Z(n362) );
  XNOR2_X1 U440 ( .A(n395), .B(n394), .ZN(n667) );
  INV_X1 U441 ( .A(KEYINPUT41), .ZN(n394) );
  INV_X1 U442 ( .A(KEYINPUT34), .ZN(n408) );
  XOR2_X1 U443 ( .A(n518), .B(G478), .Z(n533) );
  NOR2_X1 U444 ( .A1(n689), .A2(G902), .ZN(n518) );
  NOR2_X1 U445 ( .A1(n715), .A2(G952), .ZN(n697) );
  NOR2_X1 U446 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U447 ( .A1(n369), .A2(n368), .ZN(n543) );
  NAND2_X1 U448 ( .A1(n581), .A2(n404), .ZN(n635) );
  XNOR2_X1 U449 ( .A(n438), .B(n425), .ZN(n554) );
  INV_X1 U450 ( .A(KEYINPUT91), .ZN(n425) );
  XNOR2_X1 U451 ( .A(n493), .B(n448), .ZN(n372) );
  XNOR2_X1 U452 ( .A(G137), .B(G146), .ZN(n448) );
  XOR2_X1 U453 ( .A(G140), .B(G110), .Z(n471) );
  XNOR2_X1 U454 ( .A(n473), .B(n472), .ZN(n474) );
  INV_X1 U455 ( .A(KEYINPUT92), .ZN(n472) );
  XNOR2_X1 U456 ( .A(G101), .B(G146), .ZN(n473) );
  XNOR2_X1 U457 ( .A(n437), .B(KEYINPUT14), .ZN(n439) );
  NAND2_X1 U458 ( .A1(G234), .A2(G237), .ZN(n437) );
  XNOR2_X1 U459 ( .A(n536), .B(n535), .ZN(n564) );
  XNOR2_X1 U460 ( .A(n416), .B(n415), .ZN(n538) );
  INV_X1 U461 ( .A(KEYINPUT72), .ZN(n415) );
  INV_X1 U462 ( .A(n635), .ZN(n403) );
  NAND2_X1 U463 ( .A1(n367), .A2(n553), .ZN(n442) );
  XNOR2_X1 U464 ( .A(n364), .B(n363), .ZN(n367) );
  INV_X1 U465 ( .A(KEYINPUT107), .ZN(n363) );
  XNOR2_X1 U466 ( .A(n375), .B(n489), .ZN(n494) );
  XNOR2_X1 U467 ( .A(n490), .B(n488), .ZN(n375) );
  AND2_X1 U468 ( .A1(n601), .A2(n428), .ZN(n427) );
  INV_X1 U469 ( .A(KEYINPUT85), .ZN(n431) );
  INV_X1 U470 ( .A(n362), .ZN(n634) );
  AND2_X1 U471 ( .A1(n581), .A2(n481), .ZN(n482) );
  NOR2_X1 U472 ( .A1(n568), .A2(n536), .ZN(n481) );
  XNOR2_X1 U473 ( .A(n460), .B(n366), .ZN(n402) );
  XNOR2_X1 U474 ( .A(n397), .B(n516), .ZN(n689) );
  XNOR2_X1 U475 ( .A(n515), .B(n398), .ZN(n397) );
  XNOR2_X1 U476 ( .A(n517), .B(KEYINPUT101), .ZN(n398) );
  XNOR2_X1 U477 ( .A(n504), .B(n386), .ZN(n684) );
  XNOR2_X1 U478 ( .A(n505), .B(n506), .ZN(n386) );
  NOR2_X1 U479 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U480 ( .A(n359), .B(KEYINPUT40), .ZN(n724) );
  INV_X1 U481 ( .A(KEYINPUT35), .ZN(n405) );
  NAND2_X1 U482 ( .A1(n407), .A2(n350), .ZN(n406) );
  AND2_X1 U483 ( .A1(n413), .A2(n352), .ZN(n617) );
  INV_X1 U484 ( .A(KEYINPUT105), .ZN(n414) );
  XNOR2_X1 U485 ( .A(n379), .B(n378), .ZN(n584) );
  INV_X1 U486 ( .A(KEYINPUT83), .ZN(n378) );
  INV_X1 U487 ( .A(n697), .ZN(n376) );
  XNOR2_X1 U488 ( .A(n680), .B(n681), .ZN(n377) );
  XNOR2_X1 U489 ( .A(n388), .B(n387), .ZN(G75) );
  XNOR2_X1 U490 ( .A(KEYINPUT121), .B(KEYINPUT53), .ZN(n387) );
  NAND2_X1 U491 ( .A1(n389), .A2(n429), .ZN(n388) );
  AND2_X1 U492 ( .A1(n672), .A2(n706), .ZN(n389) );
  INV_X1 U493 ( .A(n568), .ZN(n404) );
  AND2_X1 U494 ( .A1(G210), .A2(n495), .ZN(n348) );
  XOR2_X2 U495 ( .A(G146), .B(G125), .Z(n349) );
  XOR2_X1 U496 ( .A(n567), .B(KEYINPUT78), .Z(n350) );
  XOR2_X1 U497 ( .A(KEYINPUT13), .B(G475), .Z(n351) );
  NOR2_X1 U498 ( .A1(n581), .A2(n640), .ZN(n352) );
  OR2_X1 U499 ( .A1(n667), .A2(n649), .ZN(n353) );
  XOR2_X1 U500 ( .A(KEYINPUT4), .B(G131), .Z(n354) );
  XNOR2_X1 U501 ( .A(KEYINPUT82), .B(KEYINPUT39), .ZN(n355) );
  XNOR2_X1 U502 ( .A(KEYINPUT77), .B(KEYINPUT19), .ZN(n356) );
  XOR2_X1 U503 ( .A(KEYINPUT67), .B(KEYINPUT32), .Z(n357) );
  XNOR2_X1 U504 ( .A(n449), .B(n372), .ZN(n451) );
  XOR2_X1 U505 ( .A(G101), .B(G113), .Z(n444) );
  NAND2_X1 U506 ( .A1(n346), .A2(n665), .ZN(n409) );
  XNOR2_X1 U507 ( .A(n409), .B(n408), .ZN(n407) );
  XNOR2_X2 U508 ( .A(n358), .B(KEYINPUT2), .ZN(n602) );
  NAND2_X1 U509 ( .A1(n410), .A2(n598), .ZN(n358) );
  NAND2_X1 U510 ( .A1(n545), .A2(n544), .ZN(n393) );
  NAND2_X1 U511 ( .A1(n551), .A2(n623), .ZN(n359) );
  NOR2_X2 U512 ( .A1(n617), .A2(n723), .ZN(n399) );
  NAND2_X1 U513 ( .A1(n538), .A2(n640), .ZN(n521) );
  NAND2_X1 U514 ( .A1(n682), .A2(G475), .ZN(n686) );
  AND2_X2 U515 ( .A1(n427), .A2(n602), .ZN(n682) );
  XNOR2_X1 U516 ( .A(n390), .B(KEYINPUT81), .ZN(n599) );
  XNOR2_X1 U517 ( .A(n373), .B(n609), .ZN(G57) );
  NOR2_X2 U518 ( .A1(n607), .A2(n697), .ZN(n373) );
  XNOR2_X1 U519 ( .A(n374), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U520 ( .A1(n676), .A2(n697), .ZN(n374) );
  NOR2_X2 U521 ( .A1(n531), .A2(n667), .ZN(n524) );
  NAND2_X1 U522 ( .A1(n523), .A2(n522), .ZN(n531) );
  NOR2_X1 U523 ( .A1(n563), .A2(n569), .ZN(n562) );
  XNOR2_X1 U524 ( .A(n583), .B(n414), .ZN(n413) );
  NOR2_X2 U525 ( .A1(n563), .A2(n362), .ZN(n583) );
  XNOR2_X1 U526 ( .A(n402), .B(n711), .ZN(n463) );
  NAND2_X1 U527 ( .A1(n600), .A2(n410), .ZN(n601) );
  NOR2_X2 U528 ( .A1(n484), .A2(n519), .ZN(n528) );
  AND2_X1 U529 ( .A1(n377), .A2(n376), .ZN(G54) );
  NAND2_X1 U530 ( .A1(n583), .A2(n582), .ZN(n379) );
  XNOR2_X1 U531 ( .A(n380), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U532 ( .A1(n687), .A2(n697), .ZN(n380) );
  NAND2_X1 U533 ( .A1(n353), .A2(n383), .ZN(n382) );
  XNOR2_X1 U534 ( .A(n384), .B(KEYINPUT118), .ZN(n383) );
  NAND2_X1 U535 ( .A1(n662), .A2(n665), .ZN(n384) );
  NAND2_X1 U536 ( .A1(n391), .A2(n633), .ZN(n390) );
  XNOR2_X1 U537 ( .A(n393), .B(n392), .ZN(n391) );
  INV_X1 U538 ( .A(KEYINPUT48), .ZN(n392) );
  INV_X1 U539 ( .A(n559), .ZN(n653) );
  NAND2_X1 U540 ( .A1(n559), .A2(n396), .ZN(n395) );
  INV_X1 U541 ( .A(n657), .ZN(n396) );
  NAND2_X1 U542 ( .A1(n399), .A2(n572), .ZN(n566) );
  NAND2_X1 U543 ( .A1(n576), .A2(n399), .ZN(n577) );
  INV_X1 U544 ( .A(n346), .ZN(n588) );
  XNOR2_X2 U545 ( .A(n400), .B(KEYINPUT22), .ZN(n563) );
  NAND2_X1 U546 ( .A1(n571), .A2(n560), .ZN(n400) );
  XNOR2_X2 U547 ( .A(n401), .B(n457), .ZN(n711) );
  XNOR2_X2 U548 ( .A(n464), .B(n465), .ZN(n581) );
  XNOR2_X2 U549 ( .A(n406), .B(n405), .ZN(n722) );
  XNOR2_X2 U550 ( .A(n496), .B(n355), .ZN(n551) );
  NOR2_X1 U551 ( .A1(n580), .A2(n579), .ZN(n596) );
  NAND2_X1 U552 ( .A1(n410), .A2(n706), .ZN(n707) );
  XNOR2_X2 U553 ( .A(n597), .B(KEYINPUT45), .ZN(n410) );
  XNOR2_X2 U554 ( .A(n411), .B(G953), .ZN(n715) );
  NOR2_X2 U555 ( .A1(n558), .A2(n557), .ZN(n412) );
  NAND2_X1 U556 ( .A1(n418), .A2(n417), .ZN(n416) );
  XNOR2_X1 U557 ( .A(n420), .B(n419), .ZN(n418) );
  INV_X1 U558 ( .A(KEYINPUT73), .ZN(n419) );
  NOR2_X2 U559 ( .A1(n519), .A2(n637), .ZN(n420) );
  NAND2_X1 U560 ( .A1(n622), .A2(n655), .ZN(n421) );
  INV_X1 U561 ( .A(n517), .ZN(n491) );
  XNOR2_X2 U562 ( .A(G116), .B(G107), .ZN(n517) );
  XNOR2_X2 U563 ( .A(n426), .B(G128), .ZN(n487) );
  NAND2_X1 U564 ( .A1(n602), .A2(n601), .ZN(n429) );
  INV_X1 U565 ( .A(n603), .ZN(n428) );
  NAND2_X1 U566 ( .A1(n587), .A2(n569), .ZN(n430) );
  NAND2_X1 U567 ( .A1(n530), .A2(n650), .ZN(n432) );
  XNOR2_X2 U568 ( .A(n433), .B(n348), .ZN(n530) );
  NAND2_X1 U569 ( .A1(n673), .A2(n603), .ZN(n433) );
  XNOR2_X1 U570 ( .A(n675), .B(n674), .ZN(n676) );
  NOR2_X1 U571 ( .A1(G902), .A2(n695), .ZN(n464) );
  XNOR2_X2 U572 ( .A(n442), .B(KEYINPUT79), .ZN(n519) );
  NAND2_X1 U573 ( .A1(n724), .A2(n725), .ZN(n526) );
  XNOR2_X1 U574 ( .A(KEYINPUT62), .B(KEYINPUT110), .ZN(n435) );
  XNOR2_X1 U575 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n436) );
  XNOR2_X1 U576 ( .A(KEYINPUT65), .B(KEYINPUT46), .ZN(n525) );
  XNOR2_X1 U577 ( .A(n526), .B(n525), .ZN(n545) );
  XNOR2_X1 U578 ( .A(n511), .B(n510), .ZN(n512) );
  AND2_X1 U579 ( .A1(n559), .A2(n404), .ZN(n560) );
  INV_X1 U580 ( .A(KEYINPUT1), .ZN(n535) );
  XNOR2_X1 U581 ( .A(n604), .B(n435), .ZN(n605) );
  XNOR2_X1 U582 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U583 ( .A(n606), .B(n605), .ZN(n607) );
  XNOR2_X1 U584 ( .A(n686), .B(n685), .ZN(n687) );
  XNOR2_X1 U585 ( .A(n608), .B(KEYINPUT63), .ZN(n609) );
  XNOR2_X1 U586 ( .A(n691), .B(n690), .ZN(n692) );
  NAND2_X1 U587 ( .A1(n439), .A2(G902), .ZN(n438) );
  NAND2_X1 U588 ( .A1(n439), .A2(G952), .ZN(n440) );
  XNOR2_X1 U589 ( .A(n440), .B(KEYINPUT88), .ZN(n664) );
  NOR2_X1 U590 ( .A1(n664), .A2(G953), .ZN(n441) );
  XNOR2_X1 U591 ( .A(n441), .B(KEYINPUT89), .ZN(n553) );
  XOR2_X1 U592 ( .A(KEYINPUT30), .B(KEYINPUT108), .Z(n453) );
  XNOR2_X1 U593 ( .A(n444), .B(n443), .ZN(n493) );
  XOR2_X1 U594 ( .A(G116), .B(KEYINPUT76), .Z(n446) );
  NAND2_X1 U595 ( .A1(n499), .A2(G210), .ZN(n445) );
  XNOR2_X1 U596 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U597 ( .A(n447), .B(KEYINPUT5), .Z(n449) );
  INV_X1 U598 ( .A(n469), .ZN(n450) );
  XNOR2_X1 U599 ( .A(n451), .B(n450), .ZN(n604) );
  NAND2_X1 U600 ( .A1(G214), .A2(n495), .ZN(n650) );
  NAND2_X1 U601 ( .A1(n537), .A2(n650), .ZN(n452) );
  XNOR2_X1 U602 ( .A(n453), .B(n452), .ZN(n483) );
  NAND2_X1 U603 ( .A1(G234), .A2(n603), .ZN(n454) );
  XNOR2_X1 U604 ( .A(KEYINPUT20), .B(n454), .ZN(n466) );
  NAND2_X1 U605 ( .A1(n466), .A2(G217), .ZN(n455) );
  XNOR2_X1 U606 ( .A(n455), .B(KEYINPUT94), .ZN(n456) );
  XNOR2_X1 U607 ( .A(KEYINPUT25), .B(n456), .ZN(n465) );
  XOR2_X1 U608 ( .A(KEYINPUT23), .B(KEYINPUT93), .Z(n459) );
  XNOR2_X1 U609 ( .A(n459), .B(n458), .ZN(n460) );
  NAND2_X1 U610 ( .A1(n715), .A2(G234), .ZN(n461) );
  XOR2_X1 U611 ( .A(KEYINPUT8), .B(n461), .Z(n514) );
  NAND2_X1 U612 ( .A1(G221), .A2(n514), .ZN(n462) );
  XNOR2_X1 U613 ( .A(n463), .B(n462), .ZN(n695) );
  NAND2_X1 U614 ( .A1(n466), .A2(G221), .ZN(n467) );
  XOR2_X1 U615 ( .A(n637), .B(KEYINPUT95), .Z(n568) );
  NAND2_X1 U616 ( .A1(G227), .A2(n715), .ZN(n477) );
  XNOR2_X1 U617 ( .A(n471), .B(n470), .ZN(n475) );
  XNOR2_X1 U618 ( .A(n477), .B(n476), .ZN(n478) );
  NOR2_X1 U619 ( .A1(G902), .A2(n677), .ZN(n480) );
  XNOR2_X1 U620 ( .A(KEYINPUT74), .B(G469), .ZN(n479) );
  NAND2_X1 U621 ( .A1(n483), .A2(n585), .ZN(n484) );
  XOR2_X1 U622 ( .A(n487), .B(n349), .Z(n489) );
  NAND2_X1 U623 ( .A1(G224), .A2(n715), .ZN(n488) );
  INV_X1 U624 ( .A(n530), .ZN(n549) );
  XNOR2_X1 U625 ( .A(KEYINPUT38), .B(n549), .ZN(n651) );
  NAND2_X1 U626 ( .A1(n528), .A2(n651), .ZN(n496) );
  XNOR2_X1 U627 ( .A(n498), .B(n497), .ZN(n506) );
  NAND2_X1 U628 ( .A1(G214), .A2(n499), .ZN(n500) );
  XNOR2_X1 U629 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U630 ( .A(n502), .B(KEYINPUT11), .Z(n505) );
  XNOR2_X1 U631 ( .A(n503), .B(n711), .ZN(n504) );
  XNOR2_X1 U632 ( .A(n527), .B(KEYINPUT99), .ZN(n532) );
  XNOR2_X1 U633 ( .A(n508), .B(n507), .ZN(n513) );
  INV_X1 U634 ( .A(n509), .ZN(n511) );
  XOR2_X1 U635 ( .A(n513), .B(n512), .Z(n516) );
  NAND2_X1 U636 ( .A1(G217), .A2(n514), .ZN(n515) );
  NAND2_X1 U637 ( .A1(n651), .A2(n650), .ZN(n657) );
  NOR2_X1 U638 ( .A1(n533), .A2(n527), .ZN(n559) );
  BUF_X1 U639 ( .A(n537), .Z(n640) );
  XNOR2_X1 U640 ( .A(KEYINPUT109), .B(KEYINPUT28), .ZN(n520) );
  XNOR2_X1 U641 ( .A(n521), .B(n520), .ZN(n523) );
  INV_X1 U642 ( .A(n536), .ZN(n522) );
  NAND2_X1 U643 ( .A1(n533), .A2(n527), .ZN(n567) );
  NAND2_X1 U644 ( .A1(n347), .A2(n528), .ZN(n529) );
  NOR2_X1 U645 ( .A1(n567), .A2(n529), .ZN(n621) );
  NAND2_X1 U646 ( .A1(n533), .A2(n532), .ZN(n628) );
  NAND2_X1 U647 ( .A1(n625), .A2(n628), .ZN(n534) );
  INV_X1 U648 ( .A(n569), .ZN(n582) );
  NOR2_X1 U649 ( .A1(n625), .A2(n582), .ZN(n539) );
  NAND2_X1 U650 ( .A1(n539), .A2(n538), .ZN(n546) );
  NOR2_X1 U651 ( .A1(n546), .A2(n540), .ZN(n541) );
  XOR2_X1 U652 ( .A(KEYINPUT36), .B(n541), .Z(n542) );
  NOR2_X1 U653 ( .A1(n634), .A2(n542), .ZN(n630) );
  NOR2_X1 U654 ( .A1(n543), .A2(n630), .ZN(n544) );
  NOR2_X1 U655 ( .A1(n362), .A2(n546), .ZN(n547) );
  NAND2_X1 U656 ( .A1(n547), .A2(n650), .ZN(n548) );
  XNOR2_X1 U657 ( .A(n548), .B(KEYINPUT43), .ZN(n550) );
  NAND2_X1 U658 ( .A1(n550), .A2(n549), .ZN(n633) );
  INV_X1 U659 ( .A(n628), .ZN(n618) );
  NAND2_X1 U660 ( .A1(n618), .A2(n551), .ZN(n632) );
  AND2_X1 U661 ( .A1(n632), .A2(KEYINPUT80), .ZN(n552) );
  AND2_X1 U662 ( .A1(n599), .A2(n552), .ZN(n598) );
  INV_X1 U663 ( .A(n553), .ZN(n556) );
  XOR2_X1 U664 ( .A(KEYINPUT90), .B(G898), .Z(n704) );
  NAND2_X1 U665 ( .A1(G953), .A2(n704), .ZN(n698) );
  NOR2_X1 U666 ( .A1(n554), .A2(n698), .ZN(n555) );
  NOR2_X1 U667 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U668 ( .A1(n634), .A2(n581), .ZN(n561) );
  INV_X1 U669 ( .A(KEYINPUT69), .ZN(n572) );
  AND2_X1 U670 ( .A1(KEYINPUT44), .A2(KEYINPUT66), .ZN(n565) );
  NAND2_X1 U671 ( .A1(n566), .A2(n565), .ZN(n578) );
  XOR2_X1 U672 ( .A(KEYINPUT33), .B(KEYINPUT75), .Z(n570) );
  XNOR2_X1 U673 ( .A(n722), .B(n572), .ZN(n574) );
  INV_X1 U674 ( .A(KEYINPUT44), .ZN(n573) );
  NAND2_X1 U675 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U676 ( .A1(n575), .A2(KEYINPUT66), .ZN(n576) );
  NAND2_X1 U677 ( .A1(n578), .A2(n577), .ZN(n580) );
  NOR2_X1 U678 ( .A1(KEYINPUT44), .A2(KEYINPUT66), .ZN(n579) );
  NOR2_X1 U679 ( .A1(n640), .A2(n588), .ZN(n586) );
  NAND2_X1 U680 ( .A1(n586), .A2(n585), .ZN(n612) );
  NAND2_X1 U681 ( .A1(n640), .A2(n587), .ZN(n645) );
  NOR2_X1 U682 ( .A1(n645), .A2(n588), .ZN(n589) );
  XNOR2_X1 U683 ( .A(n589), .B(KEYINPUT31), .ZN(n627) );
  NAND2_X1 U684 ( .A1(n612), .A2(n627), .ZN(n590) );
  NAND2_X1 U685 ( .A1(n590), .A2(n655), .ZN(n592) );
  OR2_X1 U686 ( .A1(n722), .A2(n573), .ZN(n591) );
  XNOR2_X1 U687 ( .A(n594), .B(KEYINPUT84), .ZN(n595) );
  NAND2_X1 U688 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U689 ( .A1(n714), .A2(KEYINPUT80), .ZN(n600) );
  NAND2_X1 U690 ( .A1(n682), .A2(G472), .ZN(n606) );
  INV_X1 U691 ( .A(KEYINPUT86), .ZN(n608) );
  XOR2_X1 U692 ( .A(G101), .B(n610), .Z(G3) );
  NOR2_X1 U693 ( .A1(n625), .A2(n612), .ZN(n611) );
  XOR2_X1 U694 ( .A(G104), .B(n611), .Z(G6) );
  NOR2_X1 U695 ( .A1(n612), .A2(n628), .ZN(n616) );
  XOR2_X1 U696 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n614) );
  XNOR2_X1 U697 ( .A(G107), .B(KEYINPUT111), .ZN(n613) );
  XNOR2_X1 U698 ( .A(n614), .B(n613), .ZN(n615) );
  XNOR2_X1 U699 ( .A(n616), .B(n615), .ZN(G9) );
  XOR2_X1 U700 ( .A(G110), .B(n617), .Z(G12) );
  XOR2_X1 U701 ( .A(G128), .B(KEYINPUT29), .Z(n620) );
  NAND2_X1 U702 ( .A1(n622), .A2(n618), .ZN(n619) );
  XNOR2_X1 U703 ( .A(n620), .B(n619), .ZN(G30) );
  XOR2_X1 U704 ( .A(n343), .B(n621), .Z(G45) );
  NAND2_X1 U705 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U706 ( .A(G146), .B(n624), .ZN(G48) );
  NOR2_X1 U707 ( .A1(n625), .A2(n627), .ZN(n626) );
  XOR2_X1 U708 ( .A(G113), .B(n626), .Z(G15) );
  NOR2_X1 U709 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U710 ( .A(G116), .B(n629), .Z(G18) );
  XNOR2_X1 U711 ( .A(G125), .B(n630), .ZN(n631) );
  XNOR2_X1 U712 ( .A(n631), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U713 ( .A(G134), .B(n632), .ZN(G36) );
  XNOR2_X1 U714 ( .A(G140), .B(n633), .ZN(G42) );
  NAND2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U716 ( .A(KEYINPUT50), .B(n636), .Z(n643) );
  NAND2_X1 U717 ( .A1(n637), .A2(n417), .ZN(n638) );
  XNOR2_X1 U718 ( .A(KEYINPUT49), .B(n638), .ZN(n639) );
  NOR2_X1 U719 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U720 ( .A(KEYINPUT112), .B(n641), .Z(n642) );
  NOR2_X1 U721 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U722 ( .A(KEYINPUT113), .B(n644), .ZN(n646) );
  NAND2_X1 U723 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U724 ( .A(n647), .B(KEYINPUT114), .ZN(n648) );
  XNOR2_X1 U725 ( .A(n648), .B(KEYINPUT51), .ZN(n649) );
  NOR2_X1 U726 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U727 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U728 ( .A(KEYINPUT115), .B(n654), .Z(n660) );
  INV_X1 U729 ( .A(n655), .ZN(n656) );
  XNOR2_X1 U730 ( .A(KEYINPUT116), .B(n658), .ZN(n659) );
  NOR2_X1 U731 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U732 ( .A(KEYINPUT117), .B(n661), .ZN(n662) );
  NOR2_X1 U733 ( .A1(n664), .A2(n663), .ZN(n670) );
  INV_X1 U734 ( .A(n665), .ZN(n666) );
  NOR2_X1 U735 ( .A1(n667), .A2(n666), .ZN(n668) );
  XOR2_X1 U736 ( .A(KEYINPUT119), .B(n668), .Z(n669) );
  XNOR2_X1 U737 ( .A(n671), .B(KEYINPUT120), .ZN(n672) );
  NAND2_X1 U738 ( .A1(n682), .A2(G210), .ZN(n675) );
  XNOR2_X1 U739 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n679) );
  XNOR2_X1 U740 ( .A(n677), .B(KEYINPUT57), .ZN(n678) );
  XNOR2_X1 U741 ( .A(n679), .B(n678), .ZN(n681) );
  NAND2_X1 U742 ( .A1(n693), .A2(G469), .ZN(n680) );
  XOR2_X1 U743 ( .A(KEYINPUT59), .B(KEYINPUT68), .Z(n683) );
  NAND2_X1 U744 ( .A1(n693), .A2(G478), .ZN(n691) );
  INV_X1 U745 ( .A(KEYINPUT123), .ZN(n688) );
  XNOR2_X1 U746 ( .A(n689), .B(n688), .ZN(n690) );
  NOR2_X1 U747 ( .A1(n697), .A2(n692), .ZN(G63) );
  NAND2_X1 U748 ( .A1(G217), .A2(n693), .ZN(n694) );
  INV_X1 U749 ( .A(n698), .ZN(n699) );
  NOR2_X1 U750 ( .A1(n700), .A2(n699), .ZN(n710) );
  XOR2_X1 U751 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n702) );
  NAND2_X1 U752 ( .A1(G224), .A2(G953), .ZN(n701) );
  XNOR2_X1 U753 ( .A(n702), .B(n701), .ZN(n703) );
  NOR2_X1 U754 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U755 ( .A(n705), .B(KEYINPUT125), .ZN(n708) );
  INV_X1 U756 ( .A(G953), .ZN(n706) );
  NAND2_X1 U757 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U758 ( .A(n710), .B(n709), .ZN(G69) );
  XOR2_X1 U759 ( .A(n712), .B(n711), .Z(n713) );
  XOR2_X1 U760 ( .A(KEYINPUT126), .B(n713), .Z(n717) );
  XOR2_X1 U761 ( .A(n717), .B(n714), .Z(n716) );
  NAND2_X1 U762 ( .A1(n716), .A2(n715), .ZN(n721) );
  XNOR2_X1 U763 ( .A(G227), .B(n717), .ZN(n718) );
  NAND2_X1 U764 ( .A1(n718), .A2(G900), .ZN(n719) );
  NAND2_X1 U765 ( .A1(n719), .A2(G953), .ZN(n720) );
  NAND2_X1 U766 ( .A1(n721), .A2(n720), .ZN(G72) );
  XNOR2_X1 U767 ( .A(n722), .B(G122), .ZN(G24) );
  XOR2_X1 U768 ( .A(n723), .B(G119), .Z(G21) );
  XNOR2_X1 U769 ( .A(n724), .B(G131), .ZN(G33) );
  XOR2_X1 U770 ( .A(n725), .B(G137), .Z(n726) );
  XNOR2_X1 U771 ( .A(KEYINPUT127), .B(n726), .ZN(G39) );
endmodule

