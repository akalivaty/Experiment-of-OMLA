//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 1 1 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999;
  INV_X1    g000(.A(G125), .ZN(new_n187));
  NOR3_X1   g001(.A1(new_n187), .A2(KEYINPUT16), .A3(G140), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n187), .A2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(G125), .A2(G140), .ZN(new_n192));
  AND2_X1   g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT16), .ZN(new_n194));
  OAI211_X1 g008(.A(G146), .B(new_n189), .C1(new_n193), .C2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n191), .A2(new_n192), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT75), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  AND2_X1   g012(.A1(KEYINPUT64), .A2(G146), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT64), .A2(G146), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n191), .A2(KEYINPUT75), .A3(new_n192), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n198), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XOR2_X1   g018(.A(KEYINPUT24), .B(G110), .Z(new_n205));
  XNOR2_X1  g019(.A(new_n205), .B(KEYINPUT74), .ZN(new_n206));
  INV_X1    g020(.A(G119), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G128), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G119), .ZN(new_n210));
  AND2_X1   g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n206), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT23), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n209), .A2(KEYINPUT23), .A3(G119), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(new_n208), .A3(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(G110), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n195), .B(new_n204), .C1(new_n212), .C2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G146), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n194), .B1(new_n191), .B2(new_n192), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n219), .B1(new_n220), .B2(new_n188), .ZN(new_n221));
  AOI22_X1  g035(.A1(new_n206), .A2(new_n211), .B1(new_n221), .B2(new_n195), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n216), .A2(G110), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n218), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT22), .B(G137), .ZN(new_n226));
  INV_X1    g040(.A(G953), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n227), .A2(G221), .A3(G234), .ZN(new_n228));
  XOR2_X1   g042(.A(new_n226), .B(new_n228), .Z(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n225), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n218), .A2(new_n224), .A3(new_n229), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT25), .B1(new_n233), .B2(G902), .ZN(new_n234));
  INV_X1    g048(.A(G217), .ZN(new_n235));
  INV_X1    g049(.A(G902), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n235), .B1(G234), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT25), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n231), .A2(new_n238), .A3(new_n236), .A4(new_n232), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n234), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  OR3_X1    g054(.A1(new_n233), .A2(G902), .A3(new_n237), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(G472), .A2(G902), .ZN(new_n243));
  OR2_X1    g057(.A1(KEYINPUT67), .A2(G116), .ZN(new_n244));
  NAND2_X1  g058(.A1(KEYINPUT67), .A2(G116), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G119), .ZN(new_n247));
  INV_X1    g061(.A(G116), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n248), .A2(G119), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT2), .B(G113), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n247), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n207), .B1(new_n244), .B2(new_n245), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n251), .B1(new_n254), .B2(new_n249), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n253), .A2(new_n255), .A3(KEYINPUT68), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT11), .ZN(new_n261));
  INV_X1    g075(.A(G134), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n261), .B1(new_n262), .B2(G137), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(G137), .ZN(new_n264));
  INV_X1    g078(.A(G137), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(KEYINPUT11), .A3(G134), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n263), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G131), .ZN(new_n268));
  INV_X1    g082(.A(G131), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n263), .A2(new_n266), .A3(new_n269), .A4(new_n264), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT65), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n270), .A2(new_n271), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n268), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT0), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n275), .A2(new_n209), .ZN(new_n276));
  OR2_X1    g090(.A1(KEYINPUT64), .A2(G146), .ZN(new_n277));
  INV_X1    g091(.A(G143), .ZN(new_n278));
  NAND2_X1  g092(.A1(KEYINPUT64), .A2(G146), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n278), .A2(G146), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n276), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n275), .A2(new_n209), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n278), .B1(new_n277), .B2(new_n279), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n219), .A2(G143), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n283), .A2(new_n284), .B1(new_n287), .B2(new_n276), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n274), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT30), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n270), .B(new_n271), .ZN(new_n291));
  OAI21_X1  g105(.A(G143), .B1(new_n199), .B2(new_n200), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n209), .A2(KEYINPUT1), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n292), .B(new_n293), .C1(G143), .C2(new_n219), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n209), .B1(new_n292), .B2(KEYINPUT1), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n281), .B1(new_n201), .B2(new_n278), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n265), .A2(G134), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n269), .B1(new_n264), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT66), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n299), .B(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n291), .A2(new_n297), .A3(new_n301), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n289), .A2(new_n290), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n290), .B1(new_n289), .B2(new_n302), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n260), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(G237), .A2(G953), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G210), .ZN(new_n307));
  XOR2_X1   g121(.A(new_n307), .B(KEYINPUT70), .Z(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n308), .B(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT26), .B(G101), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n310), .B(new_n311), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n253), .A2(KEYINPUT68), .A3(new_n255), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT68), .B1(new_n253), .B2(new_n255), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(new_n289), .A3(new_n302), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n305), .A2(new_n312), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT31), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT31), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n305), .A2(new_n319), .A3(new_n312), .A4(new_n316), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n289), .A2(new_n302), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n260), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT71), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(new_n324), .A3(new_n316), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n325), .B(KEYINPUT28), .C1(new_n324), .C2(new_n323), .ZN(new_n326));
  INV_X1    g140(.A(new_n316), .ZN(new_n327));
  OR2_X1    g141(.A1(new_n327), .A2(KEYINPUT28), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n312), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n243), .B1(new_n321), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(KEYINPUT32), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT32), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n332), .B(new_n243), .C1(new_n321), .C2(new_n329), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT72), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n323), .A2(new_n335), .A3(new_n316), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n322), .A2(KEYINPUT72), .A3(new_n260), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(KEYINPUT28), .A3(new_n337), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n338), .A2(new_n328), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n339), .A2(KEYINPUT73), .A3(KEYINPUT29), .A4(new_n312), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n338), .A2(KEYINPUT29), .A3(new_n328), .A4(new_n312), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT73), .ZN(new_n342));
  AOI21_X1  g156(.A(G902), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n326), .A2(new_n312), .A3(new_n328), .ZN(new_n344));
  INV_X1    g158(.A(new_n312), .ZN(new_n345));
  INV_X1    g159(.A(new_n305), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n345), .B1(new_n346), .B2(new_n327), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT29), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n344), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n340), .A2(new_n343), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G472), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n242), .B1(new_n334), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G221), .ZN(new_n353));
  XOR2_X1   g167(.A(KEYINPUT9), .B(G234), .Z(new_n354));
  AOI21_X1  g168(.A(new_n353), .B1(new_n354), .B2(new_n236), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n209), .B1(new_n282), .B2(KEYINPUT1), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n294), .B1(new_n287), .B2(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(G104), .B(G107), .ZN(new_n358));
  INV_X1    g172(.A(G101), .ZN(new_n359));
  OAI21_X1  g173(.A(KEYINPUT81), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G104), .ZN(new_n361));
  OAI21_X1  g175(.A(KEYINPUT3), .B1(new_n361), .B2(G107), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT3), .ZN(new_n363));
  INV_X1    g177(.A(G107), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(new_n364), .A3(G104), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n361), .A2(G107), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n362), .A2(new_n365), .A3(new_n359), .A4(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT81), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n364), .A2(G104), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n361), .A2(G107), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n368), .B(G101), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n360), .A2(new_n367), .A3(new_n371), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n357), .A2(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n297), .A2(new_n372), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n274), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(KEYINPUT12), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT77), .B(G140), .ZN(new_n378));
  XNOR2_X1  g192(.A(KEYINPUT76), .B(G110), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n378), .B(new_n379), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n227), .A2(G227), .ZN(new_n381));
  XOR2_X1   g195(.A(new_n380), .B(new_n381), .Z(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT82), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT10), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n357), .A2(new_n372), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n385), .B1(new_n297), .B2(new_n372), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT79), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n367), .A2(KEYINPUT78), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n362), .A2(new_n365), .A3(new_n366), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G101), .ZN(new_n392));
  AND2_X1   g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n391), .A2(KEYINPUT78), .A3(G101), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT4), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n389), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n394), .A2(KEYINPUT4), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n390), .A2(new_n392), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(KEYINPUT79), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n392), .ZN(new_n400));
  XOR2_X1   g214(.A(KEYINPUT80), .B(KEYINPUT4), .Z(new_n401));
  AOI22_X1  g215(.A1(new_n396), .A2(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n388), .B1(new_n402), .B2(new_n288), .ZN(new_n403));
  INV_X1    g217(.A(new_n274), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n384), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n400), .A2(new_n401), .ZN(new_n406));
  NOR3_X1   g220(.A1(new_n393), .A2(new_n389), .A3(new_n395), .ZN(new_n407));
  AOI21_X1  g221(.A(KEYINPUT79), .B1(new_n397), .B2(new_n398), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n288), .B(new_n406), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT1), .ZN(new_n410));
  OAI21_X1  g224(.A(G128), .B1(new_n285), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n280), .A2(new_n282), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n411), .A2(new_n412), .B1(new_n287), .B2(new_n293), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n360), .A2(new_n367), .A3(new_n371), .ZN(new_n414));
  OAI21_X1  g228(.A(KEYINPUT10), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n357), .A2(new_n372), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n415), .B1(KEYINPUT10), .B2(new_n416), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n409), .A2(new_n384), .A3(new_n404), .A4(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n377), .B(new_n383), .C1(new_n405), .C2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT83), .ZN(new_n421));
  OAI22_X1  g235(.A1(new_n405), .A2(new_n419), .B1(new_n404), .B2(new_n403), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n382), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n409), .A2(new_n404), .A3(new_n417), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT82), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n376), .B1(new_n425), .B2(new_n418), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT83), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n427), .A3(new_n383), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n421), .A2(new_n423), .A3(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G469), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(new_n430), .A3(new_n236), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n425), .A2(new_n418), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n383), .B1(new_n432), .B2(new_n377), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n404), .B1(new_n409), .B2(new_n417), .ZN(new_n434));
  AOI211_X1 g248(.A(new_n434), .B(new_n382), .C1(new_n425), .C2(new_n418), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(G469), .B1(new_n436), .B2(G902), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n355), .B1(new_n431), .B2(new_n437), .ZN(new_n438));
  AND2_X1   g252(.A1(KEYINPUT67), .A2(G116), .ZN(new_n439));
  NOR2_X1   g253(.A1(KEYINPUT67), .A2(G116), .ZN(new_n440));
  OAI21_X1  g254(.A(G122), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT14), .ZN(new_n442));
  OR2_X1    g256(.A1(new_n248), .A2(G122), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n246), .A2(KEYINPUT14), .A3(G122), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(G107), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT92), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n444), .A2(new_n445), .A3(KEYINPUT92), .A4(G107), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n441), .A2(new_n364), .A3(new_n443), .ZN(new_n451));
  XOR2_X1   g265(.A(new_n451), .B(KEYINPUT91), .Z(new_n452));
  XNOR2_X1  g266(.A(G128), .B(G143), .ZN(new_n453));
  OR2_X1    g267(.A1(new_n453), .A2(G134), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(G134), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n450), .A2(new_n452), .A3(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT90), .B(KEYINPUT13), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n209), .A2(G143), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(G134), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n441), .A2(new_n443), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(G107), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n451), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n453), .A2(new_n459), .A3(G134), .A4(new_n460), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n462), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n458), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n354), .ZN(new_n469));
  NOR3_X1   g283(.A1(new_n469), .A2(new_n235), .A3(G953), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n458), .A2(new_n467), .A3(new_n470), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n236), .ZN(new_n475));
  INV_X1    g289(.A(G478), .ZN(new_n476));
  NOR2_X1   g290(.A1(KEYINPUT93), .A2(KEYINPUT15), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(KEYINPUT93), .A2(KEYINPUT15), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n480), .ZN(new_n482));
  INV_X1    g296(.A(new_n473), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n470), .B1(new_n458), .B2(new_n467), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n236), .B(new_n482), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n481), .A2(KEYINPUT94), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT94), .ZN(new_n487));
  INV_X1    g301(.A(new_n485), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n482), .B1(new_n474), .B2(new_n236), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n306), .A2(G143), .A3(G214), .ZN(new_n492));
  AOI21_X1  g306(.A(G143), .B1(new_n306), .B2(G214), .ZN(new_n493));
  OAI21_X1  g307(.A(G131), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n306), .A2(G214), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n278), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n306), .A2(G143), .A3(G214), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n269), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT86), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT87), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n197), .B1(new_n502), .B2(KEYINPUT19), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n193), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(KEYINPUT19), .B1(new_n203), .B2(new_n502), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n202), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n494), .A2(new_n498), .A3(KEYINPUT86), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n501), .A2(new_n195), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n204), .B1(new_n219), .B2(new_n196), .ZN(new_n509));
  NAND2_X1  g323(.A1(KEYINPUT85), .A2(KEYINPUT18), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n496), .B(new_n497), .C1(new_n269), .C2(new_n510), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n509), .B(new_n511), .C1(new_n510), .C2(new_n494), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(G113), .B(G122), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(new_n361), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g331(.A(KEYINPUT17), .B(G131), .C1(new_n492), .C2(new_n493), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n195), .A2(new_n518), .A3(new_n221), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT88), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n195), .A2(new_n518), .A3(new_n221), .A4(KEYINPUT88), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT17), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n494), .A2(new_n498), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT89), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT89), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n494), .A2(new_n498), .A3(new_n526), .A4(new_n523), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n521), .A2(new_n522), .A3(new_n525), .A4(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(new_n515), .A3(new_n512), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n517), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G475), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n531), .A3(new_n236), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT20), .ZN(new_n533));
  AOI21_X1  g347(.A(G475), .B1(new_n517), .B2(new_n529), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT20), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n535), .A3(new_n236), .ZN(new_n536));
  INV_X1    g350(.A(new_n529), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n515), .B1(new_n528), .B2(new_n512), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n236), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g353(.A1(new_n533), .A2(new_n536), .B1(G475), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n227), .A2(G952), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n542), .B1(G234), .B2(G237), .ZN(new_n543));
  XOR2_X1   g357(.A(KEYINPUT21), .B(G898), .Z(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  AOI211_X1 g359(.A(new_n236), .B(new_n227), .C1(G234), .C2(G237), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n543), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NOR3_X1   g361(.A1(new_n491), .A2(new_n541), .A3(new_n547), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n260), .B(new_n406), .C1(new_n407), .C2(new_n408), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n247), .A2(KEYINPUT5), .A3(new_n250), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n550), .B(G113), .C1(KEYINPUT5), .C2(new_n250), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n551), .A2(new_n253), .A3(new_n372), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  XOR2_X1   g367(.A(G110), .B(G122), .Z(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n554), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n549), .A2(new_n552), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n555), .A2(KEYINPUT6), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n413), .A2(new_n187), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n559), .B1(new_n187), .B2(new_n288), .ZN(new_n560));
  INV_X1    g374(.A(G224), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n561), .A2(G953), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n560), .B(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT6), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n553), .A2(new_n564), .A3(new_n554), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n558), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(G210), .B1(G237), .B2(G902), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT7), .B1(new_n561), .B2(G953), .ZN(new_n568));
  OAI21_X1  g382(.A(KEYINPUT84), .B1(new_n288), .B2(new_n187), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n560), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n552), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n571), .B1(new_n402), .B2(new_n260), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n570), .B1(new_n572), .B2(new_n556), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT84), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n560), .B1(new_n574), .B2(new_n568), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n554), .B(KEYINPUT8), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n551), .A2(new_n253), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n414), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n576), .B1(new_n578), .B2(new_n552), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(G902), .B1(new_n573), .B2(new_n580), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n566), .A2(new_n567), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n567), .B1(new_n566), .B2(new_n581), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(G214), .B1(G237), .B2(G902), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n352), .A2(new_n438), .A3(new_n548), .A4(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(G101), .ZN(G3));
  INV_X1    g403(.A(new_n547), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n566), .A2(new_n581), .ZN(new_n591));
  INV_X1    g405(.A(new_n567), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n566), .A2(new_n567), .A3(new_n581), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(KEYINPUT95), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(G478), .B1(new_n474), .B2(new_n236), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT96), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT33), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(KEYINPUT96), .A2(KEYINPUT33), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n599), .B(new_n600), .C1(new_n483), .C2(new_n484), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n472), .A2(new_n597), .A3(new_n598), .A4(new_n473), .ZN(new_n602));
  AOI21_X1  g416(.A(G902), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n596), .B1(new_n603), .B2(G478), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n604), .A2(new_n540), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT95), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n566), .A2(new_n606), .A3(new_n581), .A4(new_n567), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n607), .A2(new_n585), .ZN(new_n608));
  AND4_X1   g422(.A1(new_n590), .A2(new_n595), .A3(new_n605), .A4(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n242), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n236), .B1(new_n321), .B2(new_n329), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(G472), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n330), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n438), .A2(new_n611), .A3(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(new_n361), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT97), .B(KEYINPUT34), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G6));
  INV_X1    g434(.A(KEYINPUT98), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n534), .A2(new_n535), .A3(new_n236), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n535), .B1(new_n534), .B2(new_n236), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n533), .A2(KEYINPUT98), .A3(new_n536), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n539), .A2(G475), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n491), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(new_n547), .B(KEYINPUT99), .Z(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  AND4_X1   g444(.A1(new_n595), .A2(new_n628), .A3(new_n608), .A4(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n616), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT35), .B(G107), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G9));
  NAND4_X1  g449(.A1(new_n438), .A2(new_n615), .A3(new_n587), .A4(new_n548), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n237), .A2(G902), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT100), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n218), .B2(new_n224), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n230), .A2(KEYINPUT36), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n218), .A2(new_n638), .A3(new_n224), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n641), .B1(new_n640), .B2(new_n642), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n637), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT101), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n240), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n646), .B1(new_n240), .B2(new_n645), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n636), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(KEYINPUT37), .B(G110), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G12));
  INV_X1    g466(.A(G900), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n546), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n543), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n628), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n649), .B1(new_n334), .B2(new_n351), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n607), .A2(new_n585), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n659), .B1(new_n584), .B2(KEYINPUT95), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n657), .A2(new_n658), .A3(new_n438), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G128), .ZN(G30));
  XNOR2_X1  g476(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n584), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n593), .A2(new_n594), .ZN(new_n665));
  INV_X1    g479(.A(new_n663), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n240), .A2(new_n645), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n586), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n336), .A2(new_n337), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n236), .B1(new_n672), .B2(new_n312), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n312), .B1(new_n346), .B2(new_n327), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g489(.A(G472), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n334), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n540), .B1(new_n486), .B2(new_n490), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n668), .A2(new_n670), .A3(new_n677), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT103), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n656), .B(KEYINPUT39), .Z(new_n681));
  AOI211_X1 g495(.A(new_n355), .B(new_n681), .C1(new_n431), .C2(new_n437), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT40), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G143), .ZN(G45));
  INV_X1    g501(.A(new_n656), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n604), .A2(new_n540), .A3(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n595), .A2(new_n608), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(KEYINPUT105), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n595), .A2(new_n608), .A3(new_n689), .A4(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n691), .A2(new_n438), .A3(new_n658), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  NAND2_X1  g509(.A1(new_n429), .A2(new_n236), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(G469), .ZN(new_n697));
  INV_X1    g511(.A(new_n355), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n697), .A2(new_n698), .A3(new_n431), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n352), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n700), .A2(new_n610), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT41), .B(G113), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G15));
  NOR2_X1   g517(.A1(new_n700), .A2(new_n632), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n248), .ZN(G18));
  NAND4_X1  g519(.A1(new_n699), .A2(new_n548), .A3(new_n660), .A4(new_n658), .ZN(new_n706));
  XOR2_X1   g520(.A(KEYINPUT106), .B(G119), .Z(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G21));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n338), .A2(new_n709), .A3(new_n328), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n709), .B1(new_n338), .B2(new_n328), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n710), .A2(new_n711), .A3(new_n312), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n243), .B1(new_n712), .B2(new_n321), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n611), .A3(new_n613), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n713), .A2(KEYINPUT108), .A3(new_n611), .A4(new_n613), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n660), .A2(new_n630), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n718), .A2(new_n719), .A3(new_n699), .A4(new_n678), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G122), .ZN(G24));
  NAND4_X1  g535(.A1(new_n660), .A2(new_n698), .A3(new_n431), .A4(new_n697), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n713), .A2(new_n613), .A3(new_n669), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n689), .ZN(new_n725));
  OAI21_X1  g539(.A(KEYINPUT109), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT109), .ZN(new_n727));
  INV_X1    g541(.A(new_n689), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n723), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n699), .A2(new_n727), .A3(new_n729), .A4(new_n660), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G125), .ZN(G27));
  INV_X1    g546(.A(KEYINPUT42), .ZN(new_n733));
  OAI21_X1  g547(.A(KEYINPUT111), .B1(new_n433), .B2(new_n435), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT111), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n735), .B1(new_n426), .B2(new_n383), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n734), .A2(G469), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(G469), .A2(G902), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT110), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n431), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n355), .A2(new_n586), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n352), .A2(new_n740), .A3(new_n584), .A4(new_n741), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n733), .B1(new_n742), .B2(new_n728), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n740), .A2(new_n584), .A3(new_n741), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n744), .A2(KEYINPUT42), .A3(new_n352), .A4(new_n689), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n269), .ZN(G33));
  NAND3_X1  g561(.A1(new_n744), .A2(new_n352), .A3(new_n657), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G134), .ZN(G36));
  NAND3_X1  g563(.A1(new_n734), .A2(KEYINPUT45), .A3(new_n736), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(new_n433), .B2(new_n435), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n750), .A2(G469), .A3(new_n752), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n753), .A2(KEYINPUT46), .A3(new_n739), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT46), .B1(new_n753), .B2(new_n739), .ZN(new_n755));
  INV_X1    g569(.A(new_n431), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n757), .A2(new_n355), .A3(new_n681), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n665), .A2(new_n586), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n601), .A2(new_n602), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(G478), .A3(new_n236), .ZN(new_n761));
  INV_X1    g575(.A(new_n596), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n540), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT43), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n614), .A3(new_n669), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT44), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n758), .A2(new_n759), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G137), .ZN(G39));
  INV_X1    g586(.A(KEYINPUT47), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n773), .B1(new_n757), .B2(new_n355), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n753), .A2(new_n739), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT46), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n753), .A2(KEYINPUT46), .A3(new_n739), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n431), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(KEYINPUT47), .A3(new_n698), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n774), .A2(new_n780), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n334), .A2(new_n351), .A3(new_n242), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n781), .A2(new_n689), .A3(new_n759), .A4(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G140), .ZN(G42));
  NOR2_X1   g598(.A1(G952), .A2(G953), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n699), .A2(new_n759), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n611), .A2(new_n543), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n786), .A2(new_n677), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n542), .B1(new_n788), .B2(new_n605), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n766), .A2(new_n543), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT48), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n791), .A2(new_n792), .A3(new_n352), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n792), .B1(new_n791), .B2(new_n352), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n789), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n697), .A2(new_n431), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT114), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n697), .A2(new_n799), .A3(new_n431), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n355), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n774), .A2(new_n780), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n790), .B1(new_n716), .B2(new_n717), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n759), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n796), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n786), .A2(new_n723), .A3(new_n790), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n763), .A2(new_n541), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n668), .A2(new_n585), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n804), .A2(KEYINPUT50), .A3(new_n699), .A4(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n766), .A2(new_n543), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n812), .A2(new_n810), .A3(new_n699), .A4(new_n718), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT50), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AOI221_X4 g629(.A(new_n808), .B1(new_n788), .B2(new_n809), .C1(new_n811), .C2(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n795), .B1(new_n807), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n756), .B1(new_n775), .B2(new_n776), .ZN(new_n818));
  AOI211_X1 g632(.A(new_n773), .B(new_n355), .C1(new_n818), .C2(new_n778), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT47), .B1(new_n779), .B2(new_n698), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n801), .A2(KEYINPUT115), .A3(new_n355), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT115), .B1(new_n801), .B2(new_n355), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n805), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n811), .A2(new_n815), .ZN(new_n826));
  INV_X1    g640(.A(new_n808), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n788), .A2(new_n809), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n796), .B1(new_n825), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n804), .A2(new_n660), .A3(new_n699), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n817), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT116), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n817), .A2(new_n830), .A3(KEYINPUT116), .A4(new_n831), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n699), .B(new_n352), .C1(new_n631), .C2(new_n609), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n720), .A2(new_n838), .A3(new_n706), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n481), .A2(new_n485), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n540), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n605), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n843), .A2(new_n587), .A3(new_n630), .ZN(new_n844));
  OAI221_X1 g658(.A(new_n588), .B1(new_n616), .B2(new_n844), .C1(new_n649), .C2(new_n636), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n746), .A2(new_n839), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n744), .A2(new_n729), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n840), .A2(new_n688), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n658), .A2(new_n438), .A3(new_n759), .A4(new_n848), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n626), .A2(new_n627), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n748), .B(new_n847), .C1(new_n849), .C2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n694), .A2(new_n661), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(new_n730), .B2(new_n726), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n660), .A2(new_n656), .A3(new_n678), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n669), .B1(new_n334), .B2(new_n676), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n856), .A2(new_n698), .A3(new_n740), .A4(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT52), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n694), .A2(new_n661), .ZN(new_n860));
  AND4_X1   g674(.A1(KEYINPUT52), .A2(new_n731), .A3(new_n860), .A4(new_n858), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n846), .B(new_n853), .C1(new_n859), .C2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n859), .A2(new_n861), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n862), .B(new_n863), .C1(KEYINPUT112), .C2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n731), .A2(new_n860), .A3(new_n858), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT52), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n731), .A2(new_n860), .A3(KEYINPUT52), .A4(new_n858), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n852), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT112), .B1(new_n868), .B2(new_n869), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n846), .B(new_n870), .C1(new_n871), .C2(KEYINPUT53), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n837), .B1(new_n865), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n862), .A2(new_n863), .ZN(new_n874));
  INV_X1    g688(.A(new_n845), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n839), .A2(KEYINPUT113), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT113), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n720), .A2(new_n838), .A3(new_n877), .A4(new_n706), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n863), .B1(new_n743), .B2(new_n745), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n876), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n870), .A2(new_n875), .A3(new_n880), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n874), .A2(new_n837), .A3(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n873), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n785), .B1(new_n836), .B2(new_n883), .ZN(new_n884));
  OR4_X1    g698(.A1(new_n355), .A2(new_n677), .A3(new_n586), .A4(new_n764), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n797), .B(KEYINPUT49), .Z(new_n887));
  INV_X1    g701(.A(new_n668), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n886), .A2(new_n887), .A3(new_n611), .A4(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(KEYINPUT117), .B1(new_n884), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n865), .A2(new_n872), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT54), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n874), .A2(new_n837), .A3(new_n881), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n893), .A2(new_n894), .A3(new_n834), .A4(new_n835), .ZN(new_n895));
  INV_X1    g709(.A(new_n785), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT117), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n897), .A2(new_n898), .A3(new_n889), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n891), .A2(new_n899), .ZN(G75));
  NAND2_X1  g714(.A1(new_n868), .A2(new_n869), .ZN(new_n901));
  AND4_X1   g715(.A1(new_n901), .A2(new_n880), .A3(new_n875), .A4(new_n853), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT53), .B1(new_n870), .B2(new_n846), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n904), .A2(new_n236), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(G210), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT56), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n558), .A2(new_n565), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT118), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n563), .B(KEYINPUT55), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n909), .B(new_n910), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n906), .A2(new_n907), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n911), .B1(new_n906), .B2(new_n907), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n227), .A2(G952), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(G51));
  INV_X1    g729(.A(KEYINPUT119), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n739), .B(KEYINPUT57), .Z(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT54), .B1(new_n902), .B2(new_n903), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n918), .B1(new_n919), .B2(new_n894), .ZN(new_n920));
  INV_X1    g734(.A(new_n429), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n916), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n837), .B1(new_n874), .B2(new_n881), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n917), .B1(new_n882), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n924), .A2(KEYINPUT119), .A3(new_n429), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n753), .B(KEYINPUT120), .Z(new_n926));
  NAND2_X1  g740(.A1(new_n905), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n922), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n914), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(G54));
  NAND3_X1  g744(.A1(new_n905), .A2(KEYINPUT58), .A3(G475), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n931), .A2(new_n529), .A3(new_n517), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n905), .A2(KEYINPUT58), .A3(G475), .A4(new_n530), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n932), .A2(new_n929), .A3(new_n933), .ZN(G60));
  INV_X1    g748(.A(new_n760), .ZN(new_n935));
  XNOR2_X1  g749(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n476), .A2(new_n236), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n936), .B(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n938), .B1(new_n873), .B2(new_n882), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n919), .A2(new_n894), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n940), .A2(new_n760), .A3(new_n938), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT122), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n940), .A2(KEYINPUT122), .A3(new_n760), .A4(new_n938), .ZN(new_n944));
  AOI221_X4 g758(.A(new_n914), .B1(new_n935), .B2(new_n939), .C1(new_n943), .C2(new_n944), .ZN(G63));
  INV_X1    g759(.A(KEYINPUT61), .ZN(new_n946));
  NAND2_X1  g760(.A1(G217), .A2(G902), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT123), .Z(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT60), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n233), .B1(new_n904), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(KEYINPUT124), .B1(new_n950), .B2(new_n929), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n949), .B1(new_n874), .B2(new_n881), .ZN(new_n952));
  INV_X1    g766(.A(new_n233), .ZN(new_n953));
  OAI211_X1 g767(.A(KEYINPUT124), .B(new_n929), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n952), .B1(new_n643), .B2(new_n644), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n946), .B1(new_n951), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n946), .B1(new_n950), .B2(KEYINPUT125), .ZN(new_n958));
  OR3_X1    g772(.A1(new_n952), .A2(KEYINPUT125), .A3(new_n953), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n958), .A2(new_n929), .A3(new_n955), .A4(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n957), .A2(new_n960), .ZN(G66));
  OR2_X1    g775(.A1(new_n839), .A2(new_n845), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n227), .ZN(new_n963));
  OAI21_X1  g777(.A(G953), .B1(new_n545), .B2(new_n561), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n909), .B1(G898), .B2(new_n227), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(G69));
  AND2_X1   g781(.A1(new_n783), .A2(new_n771), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n758), .A2(new_n352), .A3(new_n660), .A4(new_n678), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n855), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n970), .A2(new_n746), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n968), .A2(new_n971), .A3(new_n748), .ZN(new_n972));
  OR2_X1    g786(.A1(new_n972), .A2(G953), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n303), .A2(new_n304), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n504), .A2(new_n505), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n973), .B(new_n976), .C1(new_n653), .C2(new_n227), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n682), .A2(new_n352), .A3(new_n759), .A4(new_n843), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n686), .A2(KEYINPUT62), .A3(new_n855), .ZN(new_n979));
  AOI21_X1  g793(.A(KEYINPUT62), .B1(new_n686), .B2(new_n855), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n978), .B(new_n968), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n981), .A2(new_n227), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n977), .B1(new_n982), .B2(new_n976), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n227), .B1(G227), .B2(G900), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n984), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n977), .B(new_n986), .C1(new_n982), .C2(new_n976), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n985), .A2(new_n987), .ZN(G72));
  XOR2_X1   g802(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n989));
  NAND2_X1  g803(.A1(G472), .A2(G902), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n989), .B(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n991), .B1(new_n972), .B2(new_n962), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n992), .A2(new_n345), .A3(new_n316), .A4(new_n305), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT127), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n347), .A2(new_n994), .A3(new_n317), .ZN(new_n995));
  OR2_X1    g809(.A1(new_n347), .A2(new_n994), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n892), .A2(new_n991), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n993), .A2(new_n929), .A3(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n991), .B1(new_n981), .B2(new_n962), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n998), .B1(new_n675), .B2(new_n999), .ZN(G57));
endmodule


