

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758;

  OR2_X1 U377 ( .A1(n694), .A2(n676), .ZN(n576) );
  XNOR2_X1 U378 ( .A(n478), .B(G122), .ZN(n501) );
  XNOR2_X1 U379 ( .A(n481), .B(n480), .ZN(n736) );
  XNOR2_X1 U380 ( .A(n736), .B(n490), .ZN(n632) );
  BUF_X1 U381 ( .A(n535), .Z(n563) );
  XOR2_X1 U382 ( .A(KEYINPUT7), .B(KEYINPUT100), .Z(n355) );
  NOR2_X2 U383 ( .A1(n538), .A2(n537), .ZN(n658) );
  NAND2_X2 U384 ( .A1(n367), .A2(n639), .ZN(n593) );
  NOR2_X2 U385 ( .A1(G902), .A2(n721), .ZN(n517) );
  XNOR2_X2 U386 ( .A(n585), .B(KEYINPUT33), .ZN(n701) );
  NOR2_X2 U387 ( .A1(n600), .A2(n584), .ZN(n585) );
  NOR2_X1 U388 ( .A1(n476), .A2(n519), .ZN(n544) );
  XNOR2_X1 U389 ( .A(G119), .B(KEYINPUT3), .ZN(n432) );
  NAND2_X1 U390 ( .A1(n389), .A2(n398), .ZN(n641) );
  NAND2_X1 U391 ( .A1(n668), .A2(n617), .ZN(n401) );
  NOR2_X1 U392 ( .A1(n648), .A2(n609), .ZN(n610) );
  OR2_X1 U393 ( .A1(n755), .A2(n591), .ZN(n592) );
  XNOR2_X1 U394 ( .A(n461), .B(n460), .ZN(n578) );
  INV_X1 U395 ( .A(n432), .ZN(n433) );
  XNOR2_X1 U396 ( .A(n465), .B(G110), .ZN(n479) );
  XNOR2_X2 U397 ( .A(G116), .B(G107), .ZN(n422) );
  BUF_X1 U398 ( .A(n586), .Z(n599) );
  OR2_X1 U399 ( .A1(n717), .A2(G902), .ZN(n412) );
  INV_X1 U400 ( .A(n618), .ZN(n400) );
  XNOR2_X1 U401 ( .A(n445), .B(G125), .ZN(n484) );
  INV_X1 U402 ( .A(G146), .ZN(n445) );
  XNOR2_X1 U403 ( .A(n487), .B(G134), .ZN(n513) );
  XNOR2_X1 U404 ( .A(n468), .B(n467), .ZN(n743) );
  XNOR2_X1 U405 ( .A(n403), .B(KEYINPUT30), .ZN(n402) );
  XNOR2_X1 U406 ( .A(n411), .B(KEYINPUT28), .ZN(n522) );
  NOR2_X1 U407 ( .A1(n548), .A2(n679), .ZN(n411) );
  XNOR2_X1 U408 ( .A(n607), .B(KEYINPUT72), .ZN(n409) );
  AND2_X1 U409 ( .A1(n556), .A2(n666), .ZN(n397) );
  NOR2_X1 U410 ( .A1(n405), .A2(n404), .ZN(n546) );
  INV_X1 U411 ( .A(n637), .ZN(n404) );
  AND2_X1 U412 ( .A1(n401), .A2(n400), .ZN(n388) );
  XNOR2_X1 U413 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n483) );
  XNOR2_X1 U414 ( .A(n577), .B(KEYINPUT22), .ZN(n582) );
  NOR2_X1 U415 ( .A1(n676), .A2(n578), .ZN(n681) );
  XNOR2_X1 U416 ( .A(n479), .B(n501), .ZN(n480) );
  XNOR2_X1 U417 ( .A(n425), .B(n477), .ZN(n481) );
  XNOR2_X1 U418 ( .A(n422), .B(KEYINPUT16), .ZN(n425) );
  XOR2_X1 U419 ( .A(n355), .B(n509), .Z(n424) );
  XNOR2_X1 U420 ( .A(KEYINPUT99), .B(KEYINPUT98), .ZN(n509) );
  XNOR2_X1 U421 ( .A(n422), .B(n421), .ZN(n507) );
  INV_X1 U422 ( .A(G122), .ZN(n421) );
  XNOR2_X1 U423 ( .A(n504), .B(n503), .ZN(n624) );
  XNOR2_X1 U424 ( .A(n502), .B(n501), .ZN(n503) );
  NAND2_X1 U425 ( .A1(n370), .A2(n382), .ZN(n372) );
  NAND2_X1 U426 ( .A1(n380), .A2(n588), .ZN(n379) );
  OR2_X1 U427 ( .A1(n599), .A2(n386), .ZN(n385) );
  XNOR2_X1 U428 ( .A(n515), .B(KEYINPUT101), .ZN(n516) );
  OR2_X1 U429 ( .A1(n642), .A2(G902), .ZN(n439) );
  XNOR2_X1 U430 ( .A(n415), .B(n413), .ZN(n726) );
  XNOR2_X1 U431 ( .A(n454), .B(n414), .ZN(n413) );
  XNOR2_X1 U432 ( .A(n743), .B(n390), .ZN(n717) );
  XNOR2_X1 U433 ( .A(n466), .B(n391), .ZN(n390) );
  XNOR2_X1 U434 ( .A(n464), .B(n392), .ZN(n391) );
  NAND2_X1 U435 ( .A1(n361), .A2(n409), .ZN(n408) );
  XOR2_X1 U436 ( .A(G146), .B(G113), .Z(n435) );
  XNOR2_X1 U437 ( .A(G101), .B(G116), .ZN(n434) );
  XNOR2_X1 U438 ( .A(G131), .B(G143), .ZN(n495) );
  INV_X1 U439 ( .A(KEYINPUT64), .ZN(n399) );
  XNOR2_X1 U440 ( .A(n513), .B(n426), .ZN(n468) );
  XNOR2_X1 U441 ( .A(n394), .B(n393), .ZN(n620) );
  INV_X1 U442 ( .A(KEYINPUT48), .ZN(n393) );
  NOR2_X1 U443 ( .A1(n613), .A2(n612), .ZN(n614) );
  INV_X1 U444 ( .A(n587), .ZN(n380) );
  INV_X1 U445 ( .A(n374), .ZN(n370) );
  NAND2_X1 U446 ( .A1(n578), .A2(n520), .ZN(n548) );
  XNOR2_X1 U447 ( .A(n484), .B(n446), .ZN(n744) );
  XOR2_X1 U448 ( .A(G104), .B(G107), .Z(n463) );
  INV_X1 U449 ( .A(KEYINPUT89), .ZN(n392) );
  XNOR2_X1 U450 ( .A(G101), .B(KEYINPUT87), .ZN(n465) );
  XNOR2_X1 U451 ( .A(n506), .B(n505), .ZN(n542) );
  XNOR2_X1 U452 ( .A(n470), .B(n469), .ZN(n603) );
  XNOR2_X1 U453 ( .A(n510), .B(n424), .ZN(n511) );
  XNOR2_X1 U454 ( .A(n624), .B(KEYINPUT59), .ZN(n625) );
  XNOR2_X1 U455 ( .A(n530), .B(n529), .ZN(n756) );
  XNOR2_X1 U456 ( .A(n528), .B(KEYINPUT112), .ZN(n529) );
  NOR2_X1 U457 ( .A1(n538), .A2(n675), .ZN(n530) );
  XNOR2_X1 U458 ( .A(n518), .B(n363), .ZN(n531) );
  NAND2_X1 U459 ( .A1(n377), .A2(n375), .ZN(n755) );
  OR2_X1 U460 ( .A1(n384), .A2(n376), .ZN(n375) );
  NOR2_X1 U461 ( .A1(n381), .A2(n378), .ZN(n377) );
  NAND2_X1 U462 ( .A1(n418), .A2(n357), .ZN(n639) );
  XNOR2_X1 U463 ( .A(n420), .B(n419), .ZN(n418) );
  INV_X1 U464 ( .A(KEYINPUT104), .ZN(n419) );
  XNOR2_X1 U465 ( .A(n726), .B(n725), .ZN(n727) );
  XNOR2_X1 U466 ( .A(n719), .B(n718), .ZN(n720) );
  AND2_X1 U467 ( .A1(n401), .A2(n365), .ZN(n356) );
  AND2_X1 U468 ( .A1(n587), .A2(KEYINPUT35), .ZN(n382) );
  AND2_X1 U469 ( .A1(n578), .A2(n679), .ZN(n357) );
  AND2_X1 U470 ( .A1(n680), .A2(n578), .ZN(n358) );
  XNOR2_X1 U471 ( .A(n494), .B(KEYINPUT39), .ZN(n557) );
  AND2_X1 U472 ( .A1(n755), .A2(n591), .ZN(n359) );
  AND2_X1 U473 ( .A1(n371), .A2(n379), .ZN(n360) );
  AND2_X1 U474 ( .A1(n658), .A2(n410), .ZN(n361) );
  NOR2_X1 U475 ( .A1(n559), .A2(n368), .ZN(n362) );
  XOR2_X1 U476 ( .A(KEYINPUT109), .B(KEYINPUT40), .Z(n363) );
  XNOR2_X1 U477 ( .A(n633), .B(n632), .ZN(n364) );
  AND2_X1 U478 ( .A1(n400), .A2(n399), .ZN(n365) );
  XOR2_X1 U479 ( .A(G131), .B(KEYINPUT127), .Z(n366) );
  NAND2_X1 U480 ( .A1(n388), .A2(n623), .ZN(n387) );
  XNOR2_X1 U481 ( .A(n367), .B(G119), .ZN(G21) );
  XNOR2_X2 U482 ( .A(n580), .B(KEYINPUT32), .ZN(n367) );
  XNOR2_X2 U483 ( .A(n368), .B(n536), .ZN(n573) );
  NAND2_X2 U484 ( .A1(n417), .A2(n690), .ZN(n368) );
  NAND2_X1 U485 ( .A1(n599), .A2(n386), .ZN(n383) );
  NAND2_X1 U486 ( .A1(n369), .A2(n599), .ZN(n371) );
  AND2_X1 U487 ( .A1(n382), .A2(n386), .ZN(n369) );
  NAND2_X1 U488 ( .A1(n701), .A2(n386), .ZN(n374) );
  NAND2_X1 U489 ( .A1(n372), .A2(n360), .ZN(n378) );
  NAND2_X1 U490 ( .A1(n374), .A2(n373), .ZN(n376) );
  AND2_X1 U491 ( .A1(n383), .A2(n588), .ZN(n373) );
  AND2_X1 U492 ( .A1(n384), .A2(n382), .ZN(n381) );
  NOR2_X1 U493 ( .A1(n701), .A2(n385), .ZN(n384) );
  INV_X1 U494 ( .A(KEYINPUT34), .ZN(n386) );
  NAND2_X1 U495 ( .A1(n387), .A2(KEYINPUT64), .ZN(n389) );
  XNOR2_X1 U496 ( .A(n531), .B(n366), .ZN(G33) );
  NAND2_X1 U497 ( .A1(n620), .A2(n565), .ZN(n567) );
  NAND2_X1 U498 ( .A1(n397), .A2(n395), .ZN(n394) );
  XNOR2_X1 U499 ( .A(n532), .B(n396), .ZN(n395) );
  INV_X1 U500 ( .A(KEYINPUT46), .ZN(n396) );
  INV_X1 U501 ( .A(n401), .ZN(n671) );
  NAND2_X1 U502 ( .A1(n356), .A2(n623), .ZN(n398) );
  NAND2_X1 U503 ( .A1(n603), .A2(n402), .ZN(n476) );
  NOR2_X1 U504 ( .A1(n679), .A2(n534), .ZN(n403) );
  XNOR2_X2 U505 ( .A(n433), .B(KEYINPUT68), .ZN(n477) );
  XNOR2_X2 U506 ( .A(G113), .B(G104), .ZN(n478) );
  OR2_X2 U507 ( .A1(n594), .A2(n680), .ZN(n596) );
  NAND2_X1 U508 ( .A1(n408), .A2(n406), .ZN(n405) );
  NAND2_X1 U509 ( .A1(n407), .A2(KEYINPUT47), .ZN(n406) );
  NAND2_X1 U510 ( .A1(n539), .A2(n658), .ZN(n407) );
  INV_X1 U511 ( .A(KEYINPUT47), .ZN(n410) );
  XNOR2_X2 U512 ( .A(G143), .B(G128), .ZN(n487) );
  XNOR2_X2 U513 ( .A(n554), .B(n553), .ZN(n680) );
  XNOR2_X2 U514 ( .A(n412), .B(G469), .ZN(n554) );
  AND2_X1 U515 ( .A1(n508), .A2(G221), .ZN(n414) );
  XNOR2_X1 U516 ( .A(n416), .B(n744), .ZN(n415) );
  XNOR2_X1 U517 ( .A(n452), .B(n447), .ZN(n416) );
  NAND2_X1 U518 ( .A1(n573), .A2(n572), .ZN(n575) );
  INV_X1 U519 ( .A(n535), .ZN(n417) );
  XNOR2_X2 U520 ( .A(n493), .B(n492), .ZN(n535) );
  NAND2_X1 U521 ( .A1(n582), .A2(n581), .ZN(n420) );
  XNOR2_X1 U522 ( .A(n593), .B(n583), .ZN(n589) );
  XNOR2_X2 U523 ( .A(n439), .B(n640), .ZN(n679) );
  XNOR2_X1 U524 ( .A(KEYINPUT81), .B(KEYINPUT56), .ZN(n423) );
  AND2_X1 U525 ( .A1(n627), .A2(G953), .ZN(n730) );
  INV_X1 U526 ( .A(KEYINPUT84), .ZN(n583) );
  INV_X1 U527 ( .A(KEYINPUT10), .ZN(n446) );
  INV_X1 U528 ( .A(KEYINPUT94), .ZN(n469) );
  BUF_X1 U529 ( .A(n668), .Z(n731) );
  XNOR2_X1 U530 ( .A(n717), .B(n716), .ZN(n718) );
  XNOR2_X1 U531 ( .A(n728), .B(n727), .ZN(n729) );
  XNOR2_X1 U532 ( .A(G131), .B(KEYINPUT4), .ZN(n426) );
  XOR2_X1 U533 ( .A(KEYINPUT73), .B(KEYINPUT96), .Z(n428) );
  XNOR2_X1 U534 ( .A(G137), .B(KEYINPUT5), .ZN(n427) );
  XNOR2_X1 U535 ( .A(n428), .B(n427), .ZN(n430) );
  NOR2_X1 U536 ( .A1(G953), .A2(G237), .ZN(n498) );
  NAND2_X1 U537 ( .A1(n498), .A2(G210), .ZN(n429) );
  XNOR2_X1 U538 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U539 ( .A(n468), .B(n431), .ZN(n438) );
  XNOR2_X1 U540 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U541 ( .A(n477), .B(n436), .ZN(n437) );
  XNOR2_X1 U542 ( .A(n438), .B(n437), .ZN(n642) );
  INV_X1 U543 ( .A(G472), .ZN(n640) );
  INV_X1 U544 ( .A(G902), .ZN(n441) );
  INV_X1 U545 ( .A(G237), .ZN(n440) );
  NAND2_X1 U546 ( .A1(n441), .A2(n440), .ZN(n491) );
  NAND2_X1 U547 ( .A1(n491), .A2(G214), .ZN(n690) );
  XNOR2_X1 U548 ( .A(G902), .B(KEYINPUT15), .ZN(n618) );
  NAND2_X1 U549 ( .A1(G234), .A2(n618), .ZN(n442) );
  XNOR2_X1 U550 ( .A(KEYINPUT20), .B(n442), .ZN(n455) );
  AND2_X1 U551 ( .A1(n455), .A2(G221), .ZN(n444) );
  XNOR2_X1 U552 ( .A(KEYINPUT93), .B(KEYINPUT21), .ZN(n443) );
  XNOR2_X1 U553 ( .A(n444), .B(n443), .ZN(n676) );
  XNOR2_X1 U554 ( .A(KEYINPUT69), .B(KEYINPUT76), .ZN(n447) );
  INV_X2 U555 ( .A(G953), .ZN(n747) );
  NAND2_X1 U556 ( .A1(n747), .A2(G234), .ZN(n449) );
  XNOR2_X1 U557 ( .A(KEYINPUT67), .B(KEYINPUT8), .ZN(n448) );
  XNOR2_X1 U558 ( .A(n449), .B(n448), .ZN(n508) );
  XOR2_X1 U559 ( .A(KEYINPUT24), .B(KEYINPUT90), .Z(n451) );
  XNOR2_X1 U560 ( .A(G128), .B(KEYINPUT23), .ZN(n450) );
  XNOR2_X1 U561 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U562 ( .A(G119), .B(G110), .ZN(n453) );
  XOR2_X1 U563 ( .A(G137), .B(G140), .Z(n467) );
  XNOR2_X1 U564 ( .A(n453), .B(n467), .ZN(n454) );
  NOR2_X1 U565 ( .A1(G902), .A2(n726), .ZN(n461) );
  XNOR2_X1 U566 ( .A(KEYINPUT75), .B(KEYINPUT91), .ZN(n457) );
  NAND2_X1 U567 ( .A1(G217), .A2(n455), .ZN(n456) );
  XNOR2_X1 U568 ( .A(n457), .B(n456), .ZN(n459) );
  XOR2_X1 U569 ( .A(KEYINPUT92), .B(KEYINPUT25), .Z(n458) );
  XNOR2_X1 U570 ( .A(n459), .B(n458), .ZN(n460) );
  NAND2_X1 U571 ( .A1(G227), .A2(n747), .ZN(n462) );
  XNOR2_X1 U572 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U573 ( .A(G146), .B(n479), .ZN(n466) );
  NAND2_X1 U574 ( .A1(n681), .A2(n554), .ZN(n470) );
  NAND2_X1 U575 ( .A1(G234), .A2(G237), .ZN(n471) );
  XNOR2_X1 U576 ( .A(n471), .B(KEYINPUT14), .ZN(n472) );
  NAND2_X1 U577 ( .A1(G952), .A2(n472), .ZN(n708) );
  NOR2_X1 U578 ( .A1(G953), .A2(n708), .ZN(n570) );
  NAND2_X1 U579 ( .A1(G902), .A2(n472), .ZN(n568) );
  NOR2_X1 U580 ( .A1(G900), .A2(n568), .ZN(n473) );
  NAND2_X1 U581 ( .A1(G953), .A2(n473), .ZN(n474) );
  XOR2_X1 U582 ( .A(KEYINPUT106), .B(n474), .Z(n475) );
  NOR2_X1 U583 ( .A1(n570), .A2(n475), .ZN(n519) );
  AND2_X1 U584 ( .A1(n747), .A2(G224), .ZN(n482) );
  XNOR2_X1 U585 ( .A(n483), .B(n482), .ZN(n485) );
  XNOR2_X1 U586 ( .A(n485), .B(n484), .ZN(n489) );
  XNOR2_X1 U587 ( .A(KEYINPUT77), .B(KEYINPUT4), .ZN(n486) );
  XNOR2_X1 U588 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U589 ( .A(n489), .B(n488), .ZN(n490) );
  NAND2_X1 U590 ( .A1(n632), .A2(n618), .ZN(n493) );
  NAND2_X1 U591 ( .A1(n491), .A2(G210), .ZN(n492) );
  XNOR2_X1 U592 ( .A(n563), .B(KEYINPUT38), .ZN(n691) );
  NAND2_X1 U593 ( .A1(n544), .A2(n691), .ZN(n494) );
  XOR2_X1 U594 ( .A(KEYINPUT97), .B(G140), .Z(n496) );
  XNOR2_X1 U595 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U596 ( .A(n744), .B(n497), .ZN(n504) );
  XOR2_X1 U597 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n500) );
  NAND2_X1 U598 ( .A1(G214), .A2(n498), .ZN(n499) );
  XNOR2_X1 U599 ( .A(n500), .B(n499), .ZN(n502) );
  NOR2_X1 U600 ( .A1(G902), .A2(n624), .ZN(n506) );
  XNOR2_X1 U601 ( .A(KEYINPUT13), .B(G475), .ZN(n505) );
  XNOR2_X1 U602 ( .A(n507), .B(KEYINPUT9), .ZN(n512) );
  NAND2_X1 U603 ( .A1(G217), .A2(n508), .ZN(n510) );
  XNOR2_X1 U604 ( .A(n512), .B(n511), .ZN(n514) );
  XNOR2_X1 U605 ( .A(n514), .B(n513), .ZN(n721) );
  INV_X1 U606 ( .A(G478), .ZN(n515) );
  XNOR2_X2 U607 ( .A(n517), .B(n516), .ZN(n540) );
  NAND2_X1 U608 ( .A1(n542), .A2(n540), .ZN(n660) );
  INV_X1 U609 ( .A(n660), .ZN(n657) );
  NAND2_X1 U610 ( .A1(n557), .A2(n657), .ZN(n518) );
  NOR2_X1 U611 ( .A1(n676), .A2(n519), .ZN(n520) );
  XNOR2_X1 U612 ( .A(n554), .B(KEYINPUT108), .ZN(n521) );
  NAND2_X1 U613 ( .A1(n522), .A2(n521), .ZN(n538) );
  NAND2_X1 U614 ( .A1(n691), .A2(n690), .ZN(n523) );
  XNOR2_X1 U615 ( .A(n523), .B(KEYINPUT110), .ZN(n697) );
  INV_X1 U616 ( .A(n542), .ZN(n524) );
  NAND2_X1 U617 ( .A1(n540), .A2(n524), .ZN(n526) );
  INV_X1 U618 ( .A(KEYINPUT103), .ZN(n525) );
  XNOR2_X1 U619 ( .A(n526), .B(n525), .ZN(n694) );
  NOR2_X1 U620 ( .A1(n697), .A2(n694), .ZN(n527) );
  XNOR2_X1 U621 ( .A(n527), .B(KEYINPUT41), .ZN(n675) );
  XNOR2_X1 U622 ( .A(KEYINPUT111), .B(KEYINPUT42), .ZN(n528) );
  NAND2_X1 U623 ( .A1(n531), .A2(n756), .ZN(n532) );
  NOR2_X1 U624 ( .A1(n542), .A2(n540), .ZN(n654) );
  NOR2_X1 U625 ( .A1(n654), .A2(n657), .ZN(n533) );
  XNOR2_X1 U626 ( .A(KEYINPUT102), .B(n533), .ZN(n696) );
  INV_X1 U627 ( .A(n696), .ZN(n607) );
  INV_X1 U628 ( .A(n690), .ZN(n534) );
  XNOR2_X1 U629 ( .A(KEYINPUT74), .B(KEYINPUT19), .ZN(n536) );
  INV_X1 U630 ( .A(n573), .ZN(n537) );
  AND2_X1 U631 ( .A1(n607), .A2(KEYINPUT72), .ZN(n539) );
  INV_X1 U632 ( .A(n540), .ZN(n541) );
  NAND2_X1 U633 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U634 ( .A(n543), .B(KEYINPUT105), .ZN(n587) );
  NAND2_X1 U635 ( .A1(n544), .A2(n587), .ZN(n545) );
  OR2_X1 U636 ( .A1(n563), .A2(n545), .ZN(n637) );
  XOR2_X1 U637 ( .A(KEYINPUT71), .B(n546), .Z(n556) );
  INV_X1 U638 ( .A(KEYINPUT6), .ZN(n547) );
  XNOR2_X1 U639 ( .A(n679), .B(n547), .ZN(n584) );
  INV_X1 U640 ( .A(n584), .ZN(n550) );
  NOR2_X1 U641 ( .A1(n660), .A2(n548), .ZN(n549) );
  NAND2_X1 U642 ( .A1(n550), .A2(n549), .ZN(n559) );
  XOR2_X1 U643 ( .A(KEYINPUT85), .B(n362), .Z(n551) );
  XNOR2_X1 U644 ( .A(n551), .B(KEYINPUT36), .ZN(n555) );
  INV_X1 U645 ( .A(KEYINPUT65), .ZN(n552) );
  XNOR2_X1 U646 ( .A(n552), .B(KEYINPUT1), .ZN(n553) );
  NAND2_X1 U647 ( .A1(n555), .A2(n680), .ZN(n666) );
  NAND2_X1 U648 ( .A1(n654), .A2(n557), .ZN(n558) );
  XNOR2_X1 U649 ( .A(n558), .B(KEYINPUT113), .ZN(n754) );
  XOR2_X1 U650 ( .A(KEYINPUT43), .B(KEYINPUT107), .Z(n562) );
  NOR2_X1 U651 ( .A1(n680), .A2(n559), .ZN(n560) );
  NAND2_X1 U652 ( .A1(n560), .A2(n690), .ZN(n561) );
  XNOR2_X1 U653 ( .A(n562), .B(n561), .ZN(n564) );
  AND2_X1 U654 ( .A1(n564), .A2(n563), .ZN(n638) );
  NOR2_X1 U655 ( .A1(n754), .A2(n638), .ZN(n619) );
  AND2_X1 U656 ( .A1(n619), .A2(KEYINPUT2), .ZN(n565) );
  INV_X1 U657 ( .A(KEYINPUT80), .ZN(n566) );
  XNOR2_X1 U658 ( .A(n567), .B(n566), .ZN(n617) );
  OR2_X1 U659 ( .A1(n747), .A2(G898), .ZN(n737) );
  NOR2_X1 U660 ( .A1(n568), .A2(n737), .ZN(n569) );
  OR2_X1 U661 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U662 ( .A(n571), .B(KEYINPUT88), .ZN(n572) );
  XNOR2_X1 U663 ( .A(KEYINPUT66), .B(KEYINPUT0), .ZN(n574) );
  XNOR2_X1 U664 ( .A(n575), .B(n574), .ZN(n586) );
  NOR2_X2 U665 ( .A1(n586), .A2(n576), .ZN(n577) );
  NAND2_X1 U666 ( .A1(n582), .A2(n584), .ZN(n594) );
  INV_X1 U667 ( .A(n594), .ZN(n579) );
  INV_X1 U668 ( .A(n578), .ZN(n597) );
  NAND2_X1 U669 ( .A1(n579), .A2(n358), .ZN(n580) );
  INV_X1 U670 ( .A(n680), .ZN(n581) );
  NAND2_X1 U671 ( .A1(n681), .A2(n680), .ZN(n600) );
  INV_X1 U672 ( .A(KEYINPUT35), .ZN(n588) );
  INV_X1 U673 ( .A(KEYINPUT44), .ZN(n591) );
  NAND2_X1 U674 ( .A1(n589), .A2(n359), .ZN(n590) );
  XNOR2_X1 U675 ( .A(n590), .B(KEYINPUT70), .ZN(n615) );
  XNOR2_X1 U676 ( .A(n592), .B(KEYINPUT83), .ZN(n613) );
  NAND2_X1 U677 ( .A1(n593), .A2(KEYINPUT44), .ZN(n611) );
  INV_X1 U678 ( .A(KEYINPUT82), .ZN(n595) );
  XNOR2_X1 U679 ( .A(n596), .B(n595), .ZN(n598) );
  AND2_X1 U680 ( .A1(n598), .A2(n597), .ZN(n648) );
  INV_X1 U681 ( .A(n599), .ZN(n604) );
  NOR2_X1 U682 ( .A1(n600), .A2(n679), .ZN(n687) );
  NAND2_X1 U683 ( .A1(n604), .A2(n687), .ZN(n602) );
  INV_X1 U684 ( .A(KEYINPUT31), .ZN(n601) );
  XNOR2_X1 U685 ( .A(n602), .B(n601), .ZN(n662) );
  NAND2_X1 U686 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U687 ( .A(KEYINPUT95), .B(n605), .ZN(n606) );
  NAND2_X1 U688 ( .A1(n606), .A2(n679), .ZN(n650) );
  NAND2_X1 U689 ( .A1(n662), .A2(n650), .ZN(n608) );
  AND2_X1 U690 ( .A1(n608), .A2(n607), .ZN(n609) );
  NAND2_X1 U691 ( .A1(n611), .A2(n610), .ZN(n612) );
  NAND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X2 U693 ( .A(n616), .B(KEYINPUT45), .ZN(n668) );
  AND2_X1 U694 ( .A1(n620), .A2(n619), .ZN(n745) );
  NAND2_X1 U695 ( .A1(n668), .A2(n745), .ZN(n622) );
  INV_X1 U696 ( .A(KEYINPUT2), .ZN(n621) );
  NAND2_X1 U697 ( .A1(n622), .A2(n621), .ZN(n623) );
  INV_X2 U698 ( .A(n641), .ZN(n715) );
  NAND2_X1 U699 ( .A1(n715), .A2(G475), .ZN(n626) );
  XNOR2_X1 U700 ( .A(n626), .B(n625), .ZN(n629) );
  INV_X1 U701 ( .A(G952), .ZN(n627) );
  INV_X1 U702 ( .A(n730), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n629), .A2(n628), .ZN(n631) );
  INV_X1 U704 ( .A(KEYINPUT60), .ZN(n630) );
  XNOR2_X1 U705 ( .A(n631), .B(n630), .ZN(G60) );
  NAND2_X1 U706 ( .A1(n715), .A2(G210), .ZN(n634) );
  XOR2_X1 U707 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n633) );
  XNOR2_X1 U708 ( .A(n634), .B(n364), .ZN(n635) );
  NAND2_X1 U709 ( .A1(n635), .A2(n628), .ZN(n636) );
  XNOR2_X1 U710 ( .A(n636), .B(n423), .ZN(G51) );
  XNOR2_X1 U711 ( .A(n637), .B(G143), .ZN(G45) );
  XOR2_X1 U712 ( .A(n638), .B(G140), .Z(G42) );
  XNOR2_X1 U713 ( .A(n639), .B(G110), .ZN(G12) );
  NOR2_X1 U714 ( .A1(n641), .A2(n640), .ZN(n644) );
  XOR2_X1 U715 ( .A(KEYINPUT62), .B(n642), .Z(n643) );
  XNOR2_X1 U716 ( .A(n644), .B(n643), .ZN(n645) );
  NOR2_X1 U717 ( .A1(n645), .A2(n730), .ZN(n647) );
  XOR2_X1 U718 ( .A(KEYINPUT86), .B(KEYINPUT63), .Z(n646) );
  XNOR2_X1 U719 ( .A(n647), .B(n646), .ZN(G57) );
  XOR2_X1 U720 ( .A(G101), .B(n648), .Z(G3) );
  NOR2_X1 U721 ( .A1(n660), .A2(n650), .ZN(n649) );
  XOR2_X1 U722 ( .A(G104), .B(n649), .Z(G6) );
  INV_X1 U723 ( .A(n654), .ZN(n663) );
  NOR2_X1 U724 ( .A1(n663), .A2(n650), .ZN(n652) );
  XNOR2_X1 U725 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n651) );
  XNOR2_X1 U726 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U727 ( .A(G107), .B(n653), .ZN(G9) );
  XOR2_X1 U728 ( .A(G128), .B(KEYINPUT29), .Z(n656) );
  NAND2_X1 U729 ( .A1(n658), .A2(n654), .ZN(n655) );
  XNOR2_X1 U730 ( .A(n656), .B(n655), .ZN(G30) );
  NAND2_X1 U731 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U732 ( .A(n659), .B(G146), .ZN(G48) );
  NOR2_X1 U733 ( .A1(n660), .A2(n662), .ZN(n661) );
  XOR2_X1 U734 ( .A(G113), .B(n661), .Z(G15) );
  NOR2_X1 U735 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U736 ( .A(G116), .B(n664), .Z(G18) );
  XOR2_X1 U737 ( .A(KEYINPUT37), .B(KEYINPUT114), .Z(n665) );
  XNOR2_X1 U738 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U739 ( .A(G125), .B(n667), .ZN(G27) );
  NOR2_X1 U740 ( .A1(n731), .A2(KEYINPUT2), .ZN(n669) );
  XOR2_X1 U741 ( .A(KEYINPUT78), .B(n669), .Z(n674) );
  NOR2_X1 U742 ( .A1(KEYINPUT2), .A2(n745), .ZN(n670) );
  XOR2_X1 U743 ( .A(KEYINPUT79), .B(n670), .Z(n672) );
  NOR2_X1 U744 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U745 ( .A1(n674), .A2(n673), .ZN(n712) );
  NAND2_X1 U746 ( .A1(n578), .A2(n676), .ZN(n677) );
  XOR2_X1 U747 ( .A(KEYINPUT49), .B(n677), .Z(n678) );
  NAND2_X1 U748 ( .A1(n679), .A2(n678), .ZN(n684) );
  NOR2_X1 U749 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U750 ( .A(n682), .B(KEYINPUT50), .ZN(n683) );
  NOR2_X1 U751 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U752 ( .A(KEYINPUT115), .B(n685), .Z(n686) );
  NOR2_X1 U753 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U754 ( .A(KEYINPUT51), .B(n688), .Z(n689) );
  NOR2_X1 U755 ( .A1(n675), .A2(n689), .ZN(n704) );
  NOR2_X1 U756 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U757 ( .A(n692), .B(KEYINPUT116), .ZN(n693) );
  NOR2_X1 U758 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U759 ( .A(KEYINPUT117), .B(n695), .Z(n700) );
  NOR2_X1 U760 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U761 ( .A(KEYINPUT118), .B(n698), .ZN(n699) );
  NOR2_X1 U762 ( .A1(n700), .A2(n699), .ZN(n702) );
  NOR2_X1 U763 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U764 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U765 ( .A(n705), .B(KEYINPUT119), .Z(n706) );
  XNOR2_X1 U766 ( .A(KEYINPUT52), .B(n706), .ZN(n707) );
  NOR2_X1 U767 ( .A1(n708), .A2(n707), .ZN(n710) );
  NOR2_X1 U768 ( .A1(n701), .A2(n675), .ZN(n709) );
  NOR2_X1 U769 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U770 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U771 ( .A1(n713), .A2(G953), .ZN(n714) );
  XNOR2_X1 U772 ( .A(n714), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U773 ( .A1(n715), .A2(G469), .ZN(n719) );
  XOR2_X1 U774 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n716) );
  NOR2_X1 U775 ( .A1(n730), .A2(n720), .ZN(G54) );
  NAND2_X1 U776 ( .A1(n715), .A2(G478), .ZN(n723) );
  XNOR2_X1 U777 ( .A(n721), .B(KEYINPUT120), .ZN(n722) );
  XNOR2_X1 U778 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X1 U779 ( .A1(n730), .A2(n724), .ZN(G63) );
  NAND2_X1 U780 ( .A1(n715), .A2(G217), .ZN(n728) );
  XOR2_X1 U781 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n725) );
  NOR2_X1 U782 ( .A1(n730), .A2(n729), .ZN(G66) );
  NAND2_X1 U783 ( .A1(n731), .A2(n747), .ZN(n735) );
  NAND2_X1 U784 ( .A1(G953), .A2(G224), .ZN(n732) );
  XNOR2_X1 U785 ( .A(KEYINPUT61), .B(n732), .ZN(n733) );
  NAND2_X1 U786 ( .A1(n733), .A2(G898), .ZN(n734) );
  NAND2_X1 U787 ( .A1(n735), .A2(n734), .ZN(n742) );
  XOR2_X1 U788 ( .A(KEYINPUT123), .B(KEYINPUT125), .Z(n740) );
  XOR2_X1 U789 ( .A(n736), .B(KEYINPUT124), .Z(n738) );
  NAND2_X1 U790 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U791 ( .A(n740), .B(n739), .ZN(n741) );
  XNOR2_X1 U792 ( .A(n742), .B(n741), .ZN(G69) );
  XNOR2_X1 U793 ( .A(n744), .B(n743), .ZN(n749) );
  INV_X1 U794 ( .A(n749), .ZN(n746) );
  XNOR2_X1 U795 ( .A(n746), .B(n745), .ZN(n748) );
  NAND2_X1 U796 ( .A1(n748), .A2(n747), .ZN(n753) );
  XNOR2_X1 U797 ( .A(G227), .B(n749), .ZN(n750) );
  NAND2_X1 U798 ( .A1(n750), .A2(G900), .ZN(n751) );
  NAND2_X1 U799 ( .A1(n751), .A2(G953), .ZN(n752) );
  NAND2_X1 U800 ( .A1(n753), .A2(n752), .ZN(G72) );
  XOR2_X1 U801 ( .A(G134), .B(n754), .Z(G36) );
  XNOR2_X1 U802 ( .A(G122), .B(n755), .ZN(G24) );
  INV_X1 U803 ( .A(n756), .ZN(n757) );
  XOR2_X1 U804 ( .A(G137), .B(n757), .Z(n758) );
  XNOR2_X1 U805 ( .A(KEYINPUT126), .B(n758), .ZN(G39) );
endmodule

