//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 0 0 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 1 0 0 1 0 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n566, new_n568, new_n569, new_n570, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n617, new_n618,
    new_n620, new_n621, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  XOR2_X1   g029(.A(G325), .B(KEYINPUT65), .Z(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI21_X1  g032(.A(new_n456), .B1(new_n457), .B2(new_n452), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT66), .ZN(G319));
  NAND2_X1  g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n461), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n473), .A2(new_n464), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n475), .B1(new_n463), .B2(G2104), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n474), .A2(G137), .A3(new_n476), .A4(new_n470), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n478), .A2(G101), .A3(G2104), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n472), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NAND3_X1  g056(.A1(new_n476), .A2(new_n464), .A3(new_n473), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n482), .B(new_n483), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n484), .A2(new_n471), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT71), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n484), .A2(new_n478), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n484), .A2(KEYINPUT70), .A3(new_n478), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G136), .ZN(new_n493));
  NOR2_X1   g068(.A1(G100), .A2(G2105), .ZN(new_n494));
  XNOR2_X1  g069(.A(new_n494), .B(KEYINPUT72), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n495), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n496));
  AND3_X1   g071(.A1(new_n487), .A2(new_n493), .A3(new_n496), .ZN(G162));
  AND2_X1   g072(.A1(G126), .A2(G2105), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n476), .A2(new_n473), .A3(new_n464), .A4(new_n498), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n500), .B(G2104), .C1(G114), .C2(new_n478), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT73), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n499), .A2(new_n501), .A3(KEYINPUT73), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G138), .ZN(new_n507));
  NOR3_X1   g082(.A1(new_n468), .A2(new_n469), .A3(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT3), .B(G2104), .ZN(new_n509));
  AOI21_X1  g084(.A(KEYINPUT4), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT67), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(new_n478), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n513));
  NAND4_X1  g088(.A1(new_n512), .A2(KEYINPUT4), .A3(G138), .A4(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n482), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n506), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(G164));
  NAND2_X1  g093(.A1(KEYINPUT74), .A2(KEYINPUT5), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(KEYINPUT74), .A2(KEYINPUT5), .A3(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT6), .B(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n524), .A2(G543), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n526), .A2(G88), .B1(new_n527), .B2(G50), .ZN(new_n528));
  INV_X1    g103(.A(G62), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n529), .B1(new_n521), .B2(new_n522), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT75), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(G75), .A2(G543), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n533), .B1(new_n530), .B2(new_n531), .ZN(new_n534));
  OAI21_X1  g109(.A(G651), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT76), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n535), .A2(new_n536), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n528), .B1(new_n537), .B2(new_n538), .ZN(G303));
  INV_X1    g114(.A(G303), .ZN(G166));
  XOR2_X1   g115(.A(KEYINPUT78), .B(KEYINPUT7), .Z(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n541), .B(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n526), .A2(G89), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n545));
  XNOR2_X1  g120(.A(KEYINPUT77), .B(G51), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n527), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g122(.A1(new_n543), .A2(new_n544), .A3(new_n545), .A4(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(G168));
  AOI22_X1  g124(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G651), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g127(.A(KEYINPUT79), .B(G90), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n524), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G52), .ZN(new_n555));
  OAI22_X1  g130(.A1(new_n525), .A2(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n552), .A2(new_n556), .ZN(G171));
  AOI22_X1  g132(.A1(new_n526), .A2(G81), .B1(new_n527), .B2(G43), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT80), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n523), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n560));
  OR2_X1    g135(.A1(new_n560), .A2(new_n551), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(G860), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT81), .ZN(G153));
  AND3_X1   g140(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G36), .ZN(G176));
  XOR2_X1   g142(.A(KEYINPUT82), .B(KEYINPUT8), .Z(new_n568));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n568), .B(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(G188));
  NAND2_X1  g146(.A1(new_n527), .A2(G53), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT9), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(new_n523), .ZN(new_n575));
  INV_X1    g150(.A(G65), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n577), .A2(G651), .B1(new_n526), .B2(G91), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n573), .A2(new_n578), .ZN(G299));
  INV_X1    g154(.A(G171), .ZN(G301));
  XNOR2_X1  g155(.A(new_n548), .B(KEYINPUT83), .ZN(G286));
  AOI22_X1  g156(.A1(new_n526), .A2(G87), .B1(new_n527), .B2(G49), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(G288));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n575), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G651), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n527), .A2(G48), .ZN(new_n589));
  INV_X1    g164(.A(G86), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n525), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT84), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NOR3_X1   g168(.A1(new_n525), .A2(KEYINPUT84), .A3(new_n590), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n588), .B(new_n589), .C1(new_n593), .C2(new_n594), .ZN(G305));
  AOI22_X1  g170(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(new_n551), .ZN(new_n597));
  INV_X1    g172(.A(G85), .ZN(new_n598));
  INV_X1    g173(.A(G47), .ZN(new_n599));
  OAI22_X1  g174(.A1(new_n525), .A2(new_n598), .B1(new_n554), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(G290));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NOR2_X1   g178(.A1(G301), .A2(new_n603), .ZN(new_n604));
  AND3_X1   g179(.A1(new_n523), .A2(G92), .A3(new_n524), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT10), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n527), .A2(G54), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n523), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n606), .B(new_n607), .C1(new_n551), .C2(new_n608), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT85), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n604), .B1(new_n610), .B2(new_n603), .ZN(G284));
  XOR2_X1   g186(.A(G284), .B(KEYINPUT86), .Z(G321));
  NOR2_X1   g187(.A1(G299), .A2(G868), .ZN(new_n613));
  INV_X1    g188(.A(G286), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(G297));
  AOI21_X1  g190(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n610), .B1(new_n617), .B2(G860), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT87), .ZN(G148));
  NAND2_X1  g194(.A1(new_n562), .A2(new_n603), .ZN(new_n620));
  AND2_X1   g195(.A1(new_n610), .A2(new_n617), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n603), .ZN(G323));
  XOR2_X1   g197(.A(KEYINPUT88), .B(KEYINPUT11), .Z(new_n623));
  XNOR2_X1  g198(.A(G323), .B(new_n623), .ZN(G282));
  NAND2_X1  g199(.A1(new_n492), .A2(G135), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n485), .A2(G123), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n470), .A2(G111), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n625), .B(new_n626), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n629), .A2(G2096), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(G2096), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n478), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT12), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(G2100), .Z(new_n635));
  NAND3_X1  g210(.A1(new_n630), .A2(new_n631), .A3(new_n635), .ZN(G156));
  XNOR2_X1  g211(.A(G2427), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(KEYINPUT14), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n642), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2443), .B(G2446), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G1341), .B(G1348), .Z(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT89), .ZN(new_n650));
  OAI21_X1  g225(.A(G14), .B1(new_n647), .B2(new_n648), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(G401));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AND2_X1   g230(.A1(new_n655), .A2(KEYINPUT17), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n653), .A2(new_n654), .ZN(new_n657));
  AOI21_X1  g232(.A(KEYINPUT18), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2072), .B(G2078), .Z(new_n659));
  AOI21_X1  g234(.A(new_n659), .B1(new_n655), .B2(KEYINPUT18), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n658), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2096), .B(G2100), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G227));
  XOR2_X1   g238(.A(G1971), .B(G1976), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1956), .B(G2474), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1961), .B(G1966), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  NOR3_X1   g244(.A1(new_n665), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n665), .A2(new_n668), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT20), .Z(new_n672));
  AOI211_X1 g247(.A(new_n670), .B(new_n672), .C1(new_n665), .C2(new_n669), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT91), .ZN(new_n674));
  XOR2_X1   g249(.A(G1981), .B(G1986), .Z(new_n675));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT90), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n677), .B(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n674), .B(new_n680), .Z(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(G229));
  INV_X1    g257(.A(G29), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G33), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n492), .A2(G139), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT25), .ZN(new_n687));
  NAND2_X1  g262(.A1(G115), .A2(G2104), .ZN(new_n688));
  INV_X1    g263(.A(G127), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n688), .B1(new_n465), .B2(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n687), .B1(new_n471), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n684), .B1(new_n693), .B2(new_n683), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(G2072), .Z(new_n695));
  INV_X1    g270(.A(G16), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G4), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(new_n610), .B2(new_n696), .ZN(new_n698));
  INV_X1    g273(.A(G1348), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n695), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n683), .A2(G32), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n492), .A2(G141), .ZN(new_n703));
  NAND3_X1  g278(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT26), .Z(new_n705));
  NAND3_X1  g280(.A1(new_n478), .A2(G105), .A3(G2104), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(new_n485), .B2(G129), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n703), .A2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n702), .B1(new_n710), .B2(new_n683), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT27), .B(G1996), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G27), .ZN(new_n714));
  OR3_X1    g289(.A1(new_n714), .A2(KEYINPUT97), .A3(G29), .ZN(new_n715));
  OAI21_X1  g290(.A(KEYINPUT97), .B1(new_n714), .B2(G29), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n715), .B(new_n716), .C1(G164), .C2(new_n683), .ZN(new_n717));
  INV_X1    g292(.A(G2078), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n696), .A2(G19), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT94), .ZN(new_n721));
  INV_X1    g296(.A(new_n562), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(new_n696), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(G1341), .Z(new_n724));
  INV_X1    g299(.A(G34), .ZN(new_n725));
  AOI21_X1  g300(.A(G29), .B1(new_n725), .B2(KEYINPUT24), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(KEYINPUT24), .B2(new_n725), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n480), .B2(new_n683), .ZN(new_n728));
  INV_X1    g303(.A(G2084), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(G171), .A2(new_n696), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G5), .B2(new_n696), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n730), .B1(new_n733), .B2(G1961), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n696), .A2(G21), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G168), .B2(new_n696), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1966), .ZN(new_n737));
  INV_X1    g312(.A(G1961), .ZN(new_n738));
  OAI22_X1  g313(.A1(new_n732), .A2(new_n738), .B1(new_n729), .B2(new_n728), .ZN(new_n739));
  NOR3_X1   g314(.A1(new_n734), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  NAND4_X1  g315(.A1(new_n713), .A2(new_n719), .A3(new_n724), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT95), .B(KEYINPUT28), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n683), .A2(G26), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n492), .A2(G140), .ZN(new_n745));
  OAI21_X1  g320(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n746));
  INV_X1    g321(.A(G116), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n746), .B1(new_n471), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n485), .B2(G128), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n744), .B1(new_n750), .B2(G29), .ZN(new_n751));
  INV_X1    g326(.A(G2067), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT30), .B(G28), .ZN(new_n754));
  OR2_X1    g329(.A1(KEYINPUT31), .A2(G11), .ZN(new_n755));
  NAND2_X1  g330(.A1(KEYINPUT31), .A2(G11), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n754), .A2(new_n683), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n629), .B2(new_n683), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT96), .Z(new_n759));
  NOR4_X1   g334(.A1(new_n701), .A2(new_n741), .A3(new_n753), .A4(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n683), .A2(G35), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G162), .B2(new_n683), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT29), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n763), .A2(G2090), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n696), .A2(G20), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT23), .Z(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G299), .B2(G16), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT98), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1956), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n763), .B2(G2090), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT99), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n765), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n492), .A2(G131), .ZN(new_n775));
  OAI21_X1  g350(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n776));
  INV_X1    g351(.A(G107), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n776), .B1(new_n471), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n485), .B2(G119), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n781), .A2(new_n683), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G25), .B2(new_n683), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT92), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT35), .B(G1991), .Z(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n784), .A2(new_n786), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n696), .A2(G24), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n601), .B2(new_n696), .ZN(new_n790));
  INV_X1    g365(.A(G1986), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  NOR3_X1   g368(.A1(new_n787), .A2(new_n788), .A3(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n696), .A2(G23), .ZN(new_n796));
  INV_X1    g371(.A(G288), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(new_n696), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT33), .ZN(new_n799));
  INV_X1    g374(.A(G1976), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(G1971), .ZN(new_n802));
  NOR2_X1   g377(.A1(G16), .A2(G22), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G166), .B2(G16), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n801), .B1(new_n802), .B2(new_n805), .ZN(new_n806));
  MUX2_X1   g381(.A(G6), .B(G305), .S(G16), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT93), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT32), .B(G1981), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n806), .B(new_n810), .C1(new_n802), .C2(new_n805), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT34), .ZN(new_n812));
  OAI21_X1  g387(.A(KEYINPUT36), .B1(new_n795), .B2(new_n812), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n811), .B(KEYINPUT34), .Z(new_n814));
  INV_X1    g389(.A(KEYINPUT36), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n814), .A2(new_n815), .A3(new_n794), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n774), .B1(new_n813), .B2(new_n816), .ZN(G311));
  INV_X1    g392(.A(G311), .ZN(G150));
  NAND2_X1  g393(.A1(new_n610), .A2(G559), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT38), .Z(new_n820));
  AOI22_X1  g395(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n821), .A2(new_n551), .ZN(new_n822));
  INV_X1    g397(.A(G93), .ZN(new_n823));
  INV_X1    g398(.A(G55), .ZN(new_n824));
  OAI22_X1  g399(.A1(new_n525), .A2(new_n823), .B1(new_n554), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n562), .B(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n820), .B(new_n828), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n829), .A2(KEYINPUT39), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(KEYINPUT39), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n830), .A2(new_n563), .A3(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n826), .A2(new_n563), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT37), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n834), .ZN(G145));
  NAND2_X1  g410(.A1(new_n492), .A2(G142), .ZN(new_n836));
  INV_X1    g411(.A(new_n633), .ZN(new_n837));
  OAI21_X1  g412(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n838));
  INV_X1    g413(.A(G118), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n838), .B1(new_n471), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(new_n485), .B2(G130), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n836), .A2(new_n837), .A3(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n837), .B1(new_n836), .B2(new_n841), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n780), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n844), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n846), .A2(new_n781), .A3(new_n842), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n709), .A2(new_n750), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n499), .A2(new_n501), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n474), .A2(new_n508), .A3(KEYINPUT4), .A4(new_n476), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT4), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n512), .A2(G138), .A3(new_n513), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n852), .B1(new_n853), .B2(new_n465), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n850), .A2(new_n851), .A3(new_n854), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n703), .A2(new_n745), .A3(new_n708), .A4(new_n749), .ZN(new_n856));
  AND3_X1   g431(.A1(new_n849), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n855), .B1(new_n849), .B2(new_n856), .ZN(new_n858));
  OAI22_X1  g433(.A1(new_n857), .A2(new_n858), .B1(KEYINPUT100), .B2(new_n693), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n849), .A2(new_n856), .ZN(new_n860));
  INV_X1    g435(.A(new_n855), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n849), .A2(new_n855), .A3(new_n856), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT100), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n692), .B(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n862), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n848), .B1(new_n859), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT103), .ZN(new_n868));
  AND2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n629), .B(new_n480), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(G162), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(new_n867), .B2(new_n868), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n859), .A2(new_n866), .A3(new_n848), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(KEYINPUT101), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT101), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n859), .A2(new_n866), .A3(new_n876), .A4(new_n848), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(G37), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n867), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n871), .ZN(new_n882));
  AOI21_X1  g457(.A(KEYINPUT102), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n867), .B1(new_n875), .B2(new_n877), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT102), .ZN(new_n885));
  NOR3_X1   g460(.A1(new_n884), .A2(new_n885), .A3(new_n871), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n879), .B(KEYINPUT40), .C1(new_n883), .C2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n881), .A2(KEYINPUT102), .A3(new_n882), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n885), .B1(new_n884), .B2(new_n871), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(KEYINPUT40), .B1(new_n891), .B2(new_n879), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n888), .A2(new_n892), .ZN(G395));
  XNOR2_X1  g468(.A(G288), .B(new_n601), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n894), .B(KEYINPUT105), .Z(new_n895));
  XOR2_X1   g470(.A(G303), .B(G305), .Z(new_n896));
  OR2_X1    g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n896), .B1(KEYINPUT105), .B2(new_n894), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT42), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n621), .B(new_n828), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n609), .B(G299), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  OR3_X1    g479(.A1(new_n902), .A2(KEYINPUT104), .A3(KEYINPUT41), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT104), .B1(new_n902), .B2(KEYINPUT41), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n902), .A2(KEYINPUT41), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n909), .A2(new_n901), .ZN(new_n910));
  NOR3_X1   g485(.A1(new_n900), .A2(new_n904), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n901), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n912), .B1(new_n903), .B2(new_n901), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n900), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(G868), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n826), .A2(G868), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(G295));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n915), .A2(new_n919), .A3(new_n917), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n919), .B1(new_n915), .B2(new_n917), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(G331));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n923));
  INV_X1    g498(.A(G37), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n828), .A2(KEYINPUT107), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n828), .A2(KEYINPUT107), .ZN(new_n927));
  NAND2_X1  g502(.A1(G301), .A2(new_n548), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(G286), .B2(G301), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NOR3_X1   g505(.A1(new_n926), .A2(new_n927), .A3(new_n930), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n828), .A2(KEYINPUT107), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n929), .B1(new_n932), .B2(new_n925), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n903), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n930), .B1(new_n926), .B2(new_n927), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n932), .A2(new_n925), .A3(new_n929), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(new_n908), .A3(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n934), .A2(new_n899), .A3(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n934), .ZN(new_n939));
  XOR2_X1   g514(.A(new_n902), .B(KEYINPUT41), .Z(new_n940));
  NOR3_X1   g515(.A1(new_n931), .A2(new_n933), .A3(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n924), .B(new_n938), .C1(new_n942), .C2(new_n899), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n923), .B1(new_n943), .B2(KEYINPUT43), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n938), .A2(new_n924), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n899), .B1(new_n934), .B2(new_n937), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n945), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT108), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n945), .A2(KEYINPUT108), .A3(new_n946), .A4(new_n948), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n944), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n938), .A2(new_n924), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT43), .B1(new_n954), .B2(new_n947), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n955), .B1(new_n943), .B2(KEYINPUT43), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n923), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n953), .A2(new_n957), .ZN(G397));
  AOI21_X1  g533(.A(G1384), .B1(new_n516), .B2(new_n850), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n959), .A2(KEYINPUT45), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n472), .A2(new_n477), .A3(G40), .A4(new_n479), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n963), .B(KEYINPUT109), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n965), .A2(new_n710), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n963), .A2(G1996), .ZN(new_n967));
  AOI22_X1  g542(.A1(new_n966), .A2(G1996), .B1(new_n710), .B2(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n750), .A2(G2067), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n752), .B1(new_n745), .B2(new_n749), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n964), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n781), .A2(new_n785), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n780), .A2(new_n786), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n964), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n963), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n601), .B(new_n791), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G1384), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT45), .B1(new_n517), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n855), .A2(KEYINPUT45), .A3(new_n980), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n962), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT53), .B1(new_n984), .B2(new_n718), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT50), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n855), .A2(new_n986), .A3(new_n980), .ZN(new_n987));
  AOI21_X1  g562(.A(G1384), .B1(new_n506), .B2(new_n516), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n962), .B(new_n987), .C1(new_n988), .C2(new_n986), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n985), .B1(new_n738), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n855), .A2(new_n980), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n961), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n517), .A2(KEYINPUT45), .A3(new_n980), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n993), .A2(new_n994), .A3(KEYINPUT53), .A4(new_n718), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n990), .A2(G301), .A3(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n996), .B(KEYINPUT123), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT54), .ZN(new_n998));
  INV_X1    g573(.A(new_n993), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(KEYINPUT121), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(KEYINPUT121), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT122), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT53), .B1(new_n1002), .B2(G2078), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1003), .B1(new_n1002), .B2(G2078), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1001), .A2(new_n982), .A3(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n990), .B1(new_n1000), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n998), .B1(new_n1006), .B2(G171), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n997), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT114), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(new_n989), .B2(G2084), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n986), .B1(new_n517), .B2(new_n980), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n987), .A2(new_n962), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1012), .A2(KEYINPUT114), .A3(new_n729), .A4(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n993), .A2(new_n994), .ZN(new_n1016));
  INV_X1    g591(.A(G1966), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1010), .A2(new_n1015), .A3(new_n1018), .A4(G168), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(G8), .ZN(new_n1020));
  AOI21_X1  g595(.A(G1966), .B1(new_n993), .B2(new_n994), .ZN(new_n1021));
  NOR3_X1   g596(.A1(new_n1011), .A2(new_n1013), .A3(G2084), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1021), .B1(new_n1022), .B2(KEYINPUT114), .ZN(new_n1023));
  AOI21_X1  g598(.A(G168), .B1(new_n1023), .B2(new_n1010), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT51), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1019), .A2(new_n1026), .A3(G8), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G8), .ZN(new_n1029));
  OR2_X1    g604(.A1(new_n989), .A2(G2090), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n802), .B1(new_n981), .B2(new_n983), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1029), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1033), .B1(G166), .B2(new_n1029), .ZN(new_n1034));
  NAND3_X1  g609(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1032), .A2(new_n1036), .ZN(new_n1037));
  OAI221_X1 g612(.A(G8), .B1(G288), .B2(new_n800), .C1(new_n961), .C2(new_n991), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT52), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1039), .A2(KEYINPUT110), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n991), .A2(new_n961), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1043), .A2(new_n1029), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n797), .A2(G1976), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(new_n1045), .A3(new_n1040), .ZN(new_n1046));
  XNOR2_X1  g621(.A(KEYINPUT111), .B(G1976), .ZN(new_n1047));
  OR3_X1    g622(.A1(new_n797), .A2(KEYINPUT52), .A3(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1042), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n588), .A2(new_n589), .ZN(new_n1050));
  OAI21_X1  g625(.A(G1981), .B1(new_n1050), .B2(new_n591), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1051), .B1(G305), .B2(G1981), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT49), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1051), .B(KEYINPUT49), .C1(G1981), .C2(G305), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1054), .A2(new_n1055), .A3(new_n1044), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1049), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1037), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1036), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT112), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n986), .B1(new_n855), .B2(new_n980), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1060), .B1(new_n1061), .B2(new_n961), .ZN(new_n1062));
  OAI211_X1 g637(.A(KEYINPUT112), .B(new_n962), .C1(new_n959), .C2(new_n986), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n988), .A2(new_n986), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1031), .B1(new_n1065), .B2(G2090), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT113), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT113), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1068), .B(new_n1031), .C1(new_n1065), .C2(G2090), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1067), .A2(G8), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1058), .B1(new_n1059), .B2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1006), .A2(G171), .ZN(new_n1072));
  AOI21_X1  g647(.A(G301), .B1(new_n990), .B2(new_n995), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n998), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1008), .A2(new_n1028), .A3(new_n1071), .A4(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g650(.A(KEYINPUT58), .B(G1341), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1043), .A2(new_n1076), .ZN(new_n1077));
  XOR2_X1   g652(.A(KEYINPUT117), .B(G1996), .Z(new_n1078));
  AOI21_X1  g653(.A(new_n1077), .B1(new_n984), .B2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1079), .A2(new_n562), .ZN(new_n1080));
  XNOR2_X1  g655(.A(new_n1080), .B(KEYINPUT59), .ZN(new_n1081));
  INV_X1    g656(.A(G1956), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1065), .A2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1085), .B1(new_n573), .B2(new_n578), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g662(.A(KEYINPUT56), .B(G2072), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n984), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1083), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT61), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1065), .A2(new_n1082), .B1(new_n984), .B2(new_n1088), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1087), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1091), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1081), .B1(new_n1090), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT116), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1090), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1092), .A2(KEYINPUT116), .A3(new_n1087), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1098), .A2(new_n1099), .B1(new_n1094), .B2(new_n1093), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1100), .A2(new_n1101), .A3(KEYINPUT61), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1103));
  AND4_X1   g678(.A1(KEYINPUT116), .A2(new_n1083), .A3(new_n1087), .A4(new_n1089), .ZN(new_n1104));
  AOI21_X1  g679(.A(KEYINPUT116), .B1(new_n1092), .B2(new_n1087), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1103), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT118), .B1(new_n1106), .B2(new_n1091), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1096), .B1(new_n1102), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  OAI211_X1 g685(.A(KEYINPUT119), .B(new_n1096), .C1(new_n1102), .C2(new_n1107), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n989), .A2(new_n699), .B1(new_n752), .B2(new_n1043), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT60), .B1(new_n609), .B2(KEYINPUT120), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n609), .A2(KEYINPUT120), .ZN(new_n1115));
  OR3_X1    g690(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1115), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1116), .B(new_n1117), .C1(KEYINPUT60), .C2(new_n1112), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1110), .A2(new_n1111), .A3(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1103), .B1(new_n1112), .B2(new_n609), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1120), .B1(new_n1105), .B2(new_n1104), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1075), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT62), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1025), .A2(new_n1124), .A3(new_n1027), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1070), .A2(new_n1059), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1126), .A2(new_n1037), .A3(new_n1057), .A4(new_n1073), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1123), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1025), .A2(new_n1124), .A3(new_n1027), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1071), .A2(new_n1129), .A3(KEYINPUT124), .A4(new_n1073), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1028), .A2(KEYINPUT62), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1128), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(KEYINPUT125), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT125), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1128), .A2(new_n1130), .A3(new_n1134), .A4(new_n1131), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1056), .A2(new_n800), .A3(new_n797), .ZN(new_n1136));
  NOR2_X1   g711(.A1(G305), .A2(G1981), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1044), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1057), .A2(new_n1036), .A3(new_n1032), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT115), .ZN(new_n1141));
  OAI21_X1  g716(.A(KEYINPUT63), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1058), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1023), .A2(new_n1010), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1144), .A2(G8), .A3(new_n614), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1141), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1147));
  NOR4_X1   g722(.A1(new_n1058), .A2(new_n1142), .A3(new_n1145), .A4(KEYINPUT115), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1071), .A2(new_n1146), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT63), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1140), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1133), .A2(new_n1135), .A3(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n979), .B1(new_n1122), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n969), .B1(new_n972), .B2(new_n974), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1156), .A2(new_n965), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1157), .A2(KEYINPUT126), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1157), .A2(KEYINPUT126), .ZN(new_n1159));
  XOR2_X1   g734(.A(new_n967), .B(KEYINPUT46), .Z(new_n1160));
  OAI211_X1 g735(.A(new_n1160), .B(new_n971), .C1(new_n710), .C2(new_n965), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1161), .B(KEYINPUT47), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n963), .A2(G1986), .A3(G290), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1163), .B(KEYINPUT48), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1162), .B1(new_n976), .B2(new_n1164), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n1158), .A2(new_n1159), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1155), .A2(new_n1166), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g742(.A1(new_n891), .A2(new_n879), .ZN(new_n1169));
  NOR2_X1   g743(.A1(G227), .A2(new_n458), .ZN(new_n1170));
  INV_X1    g744(.A(new_n1170), .ZN(new_n1171));
  OAI21_X1  g745(.A(KEYINPUT127), .B1(G401), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g746(.A1(new_n1172), .A2(new_n681), .ZN(new_n1173));
  NOR3_X1   g747(.A1(G401), .A2(KEYINPUT127), .A3(new_n1171), .ZN(new_n1174));
  NOR2_X1   g748(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g749(.A1(new_n1169), .A2(new_n956), .A3(new_n1175), .ZN(G225));
  INV_X1    g750(.A(G225), .ZN(G308));
endmodule


