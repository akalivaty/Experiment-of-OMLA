//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 0 0 0 1 0 1 1 0 1 1 0 0 0 1 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 0 0 1 1 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1272, new_n1273,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343;
  INV_X1    g0000(.A(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G58), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT0), .Z(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G107), .A2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n212), .B(new_n213), .C1(new_n201), .C2(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G50), .ZN(new_n217));
  INV_X1    g0017(.A(G226), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n202), .C2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G58), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n208), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT64), .ZN(new_n229));
  OAI21_X1  g0029(.A(G50), .B1(G58), .B2(G68), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n211), .B(new_n225), .C1(new_n229), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G264), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(new_n222), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n235), .B(new_n239), .Z(G358));
  NOR2_X1   g0040(.A1(new_n201), .A2(new_n202), .ZN(new_n241));
  INV_X1    g0041(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(new_n203), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n243), .B(KEYINPUT65), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  INV_X1    g0050(.A(KEYINPUT14), .ZN(new_n251));
  INV_X1    g0051(.A(G41), .ZN(new_n252));
  INV_X1    g0052(.A(G45), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AND2_X1   g0054(.A1(KEYINPUT66), .A2(G1), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT66), .A2(G1), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  OAI211_X1 g0058(.A(G1), .B(G13), .C1(new_n258), .C2(new_n252), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G238), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n254), .A2(new_n263), .A3(G274), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT71), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n264), .B(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G97), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n222), .A2(G1698), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n268), .B1(G226), .B2(G1698), .ZN(new_n269));
  AND2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NOR2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n267), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n262), .A2(new_n266), .A3(new_n275), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT72), .B(KEYINPUT13), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n277), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n262), .A2(new_n266), .A3(new_n275), .A4(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n251), .B1(new_n281), .B2(G169), .ZN(new_n282));
  INV_X1    g0082(.A(G169), .ZN(new_n283));
  AOI211_X1 g0083(.A(KEYINPUT14), .B(new_n283), .C1(new_n278), .C2(new_n280), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT73), .ZN(new_n286));
  OR2_X1    g0086(.A1(new_n280), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n276), .A2(KEYINPUT13), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n280), .A2(new_n286), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n287), .A2(G179), .A3(new_n288), .A4(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g0091(.A(G13), .B(G20), .C1(new_n255), .C2(new_n256), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n201), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT12), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT66), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n263), .ZN(new_n297));
  NAND2_X1  g0097(.A1(KEYINPUT66), .A2(G1), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n227), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n226), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n295), .B1(new_n201), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n301), .ZN(new_n305));
  OAI21_X1  g0105(.A(KEYINPUT68), .B1(new_n258), .B2(G20), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT68), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n307), .A2(new_n227), .A3(G33), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n306), .A2(new_n308), .A3(G77), .ZN(new_n309));
  NOR2_X1   g0109(.A1(G20), .A2(G33), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n310), .A2(G50), .B1(G20), .B2(new_n201), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n305), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n312), .B(KEYINPUT11), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n304), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n291), .A2(new_n315), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n287), .A2(G190), .A3(new_n288), .A4(new_n289), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n281), .A2(G200), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n317), .A2(new_n314), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(KEYINPUT74), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT16), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT3), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n258), .ZN(new_n324));
  NAND2_X1  g0124(.A1(KEYINPUT3), .A2(G33), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(new_n227), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT7), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n324), .A2(KEYINPUT7), .A3(new_n227), .A4(new_n325), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n201), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AND2_X1   g0130(.A1(G58), .A2(G68), .ZN(new_n331));
  NOR2_X1   g0131(.A1(G58), .A2(G68), .ZN(new_n332));
  OAI21_X1  g0132(.A(G20), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n310), .A2(G159), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n322), .B1(new_n330), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT76), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(KEYINPUT7), .B1(new_n272), .B2(new_n227), .ZN(new_n339));
  INV_X1    g0139(.A(new_n329), .ZN(new_n340));
  OAI21_X1  g0140(.A(G68), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT75), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n342), .B1(new_n333), .B2(new_n334), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n335), .A2(KEYINPUT75), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n341), .B(KEYINPUT16), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  OAI211_X1 g0145(.A(KEYINPUT76), .B(new_n322), .C1(new_n330), .C2(new_n335), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n338), .A2(new_n301), .A3(new_n345), .A4(new_n346), .ZN(new_n347));
  XNOR2_X1  g0147(.A(KEYINPUT8), .B(G58), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT77), .ZN(new_n349));
  NOR3_X1   g0149(.A1(new_n299), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  XOR2_X1   g0150(.A(KEYINPUT8), .B(G58), .Z(new_n351));
  OAI21_X1  g0151(.A(G20), .B1(new_n255), .B2(new_n256), .ZN(new_n352));
  AOI21_X1  g0152(.A(KEYINPUT77), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n292), .A2(new_n305), .ZN(new_n354));
  NOR3_X1   g0154(.A1(new_n350), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n292), .A2(new_n351), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT78), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT78), .ZN(new_n358));
  INV_X1    g0158(.A(new_n356), .ZN(new_n359));
  INV_X1    g0159(.A(new_n353), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n351), .A2(new_n352), .A3(KEYINPUT77), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n358), .B(new_n359), .C1(new_n362), .C2(new_n354), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n357), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n347), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n257), .A2(G232), .A3(new_n259), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT80), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n257), .A2(KEYINPUT80), .A3(G232), .A4(new_n259), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n264), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT79), .ZN(new_n372));
  OR2_X1    g0172(.A1(G223), .A2(G1698), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n218), .A2(G1698), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n373), .B(new_n374), .C1(new_n270), .C2(new_n271), .ZN(new_n375));
  NAND2_X1  g0175(.A1(G33), .A2(G87), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n372), .B1(new_n377), .B2(new_n274), .ZN(new_n378));
  AOI211_X1 g0178(.A(KEYINPUT79), .B(new_n259), .C1(new_n375), .C2(new_n376), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n371), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(G179), .ZN(new_n382));
  INV_X1    g0182(.A(new_n264), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n383), .B1(new_n368), .B2(new_n369), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n377), .A2(new_n274), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n381), .A2(new_n382), .B1(new_n283), .B2(new_n386), .ZN(new_n387));
  AND3_X1   g0187(.A1(new_n365), .A2(KEYINPUT18), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(KEYINPUT18), .B1(new_n365), .B2(new_n387), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(G200), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  XOR2_X1   g0192(.A(KEYINPUT81), .B(G190), .Z(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n384), .B(new_n394), .C1(new_n378), .C2(new_n379), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n396), .A2(new_n364), .A3(new_n347), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT17), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n396), .A2(KEYINPUT17), .A3(new_n347), .A4(new_n364), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n390), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n324), .A2(new_n325), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G238), .A2(G1698), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n403), .B(new_n404), .C1(new_n222), .C2(G1698), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n405), .B(new_n274), .C1(G107), .C2(new_n403), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n406), .B(new_n264), .C1(new_n219), .C2(new_n260), .ZN(new_n407));
  INV_X1    g0207(.A(G190), .ZN(new_n408));
  OR2_X1    g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G20), .A2(G77), .ZN(new_n410));
  INV_X1    g0210(.A(new_n310), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n306), .A2(new_n308), .ZN(new_n412));
  XNOR2_X1  g0212(.A(KEYINPUT15), .B(G87), .ZN(new_n413));
  OAI221_X1 g0213(.A(new_n410), .B1(new_n348), .B2(new_n411), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n414), .A2(new_n301), .B1(new_n202), .B2(new_n293), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT70), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n302), .A2(G77), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n415), .A2(new_n417), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT70), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n407), .A2(G200), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n409), .A2(new_n418), .A3(new_n420), .A4(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n321), .A2(new_n402), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n420), .A2(new_n418), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n407), .A2(new_n283), .ZN(new_n425));
  OR2_X1    g0225(.A1(new_n407), .A2(G179), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n227), .B1(new_n332), .B2(new_n217), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT69), .ZN(new_n430));
  XNOR2_X1  g0230(.A(new_n429), .B(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n310), .A2(G150), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n431), .B(new_n432), .C1(new_n412), .C2(new_n348), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n301), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n293), .A2(new_n217), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n302), .A2(G50), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n434), .A2(KEYINPUT9), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(G1698), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(G222), .ZN(new_n439));
  XNOR2_X1  g0239(.A(KEYINPUT67), .B(G223), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n403), .B(new_n439), .C1(new_n440), .C2(new_n438), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n441), .B(new_n274), .C1(G77), .C2(new_n403), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n261), .A2(G226), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(new_n264), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(G200), .ZN(new_n445));
  OR2_X1    g0245(.A1(new_n444), .A2(new_n408), .ZN(new_n446));
  AND3_X1   g0246(.A1(new_n437), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT10), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n433), .A2(new_n301), .B1(new_n217), .B2(new_n293), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT9), .B1(new_n449), .B2(new_n436), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n447), .A2(new_n448), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n437), .A2(new_n445), .A3(new_n446), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT10), .B1(new_n453), .B2(new_n450), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n449), .A2(new_n436), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n444), .A2(new_n283), .ZN(new_n457));
  OR2_X1    g0257(.A1(new_n444), .A2(G179), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n455), .B(new_n459), .C1(new_n320), .C2(KEYINPUT74), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n423), .A2(new_n428), .A3(new_n460), .ZN(new_n461));
  AND2_X1   g0261(.A1(G264), .A2(G1698), .ZN(new_n462));
  AOI21_X1  g0262(.A(KEYINPUT88), .B1(new_n403), .B2(new_n462), .ZN(new_n463));
  OAI211_X1 g0263(.A(KEYINPUT88), .B(new_n462), .C1(new_n270), .C2(new_n271), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G303), .ZN(new_n466));
  OAI22_X1  g0266(.A1(new_n463), .A2(new_n465), .B1(new_n466), .B2(new_n403), .ZN(new_n467));
  OAI211_X1 g0267(.A(G257), .B(new_n438), .C1(new_n270), .C2(new_n271), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT87), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n403), .A2(KEYINPUT87), .A3(G257), .A4(new_n438), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n274), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n297), .A2(new_n298), .ZN(new_n474));
  XNOR2_X1  g0274(.A(KEYINPUT5), .B(G41), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n474), .A2(new_n475), .A3(G45), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n476), .A2(G270), .A3(new_n259), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n253), .B1(new_n297), .B2(new_n298), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n478), .A2(G274), .A3(new_n259), .A4(new_n475), .ZN(new_n479));
  AND2_X1   g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n473), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n474), .A2(G33), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(new_n305), .A3(new_n292), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G116), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G283), .ZN(new_n486));
  INV_X1    g0286(.A(G97), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n486), .B(new_n227), .C1(G33), .C2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G116), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G20), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n301), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT20), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n488), .A2(KEYINPUT20), .A3(new_n301), .A4(new_n490), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n493), .A2(new_n494), .B1(new_n489), .B2(new_n293), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n485), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n481), .A2(G169), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT21), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n497), .A2(KEYINPUT89), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n473), .A2(new_n480), .A3(G179), .ZN(new_n500));
  INV_X1    g0300(.A(new_n496), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n498), .B1(new_n497), .B2(KEYINPUT89), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n481), .A2(new_n394), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n391), .B1(new_n473), .B2(new_n480), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n506), .A2(new_n496), .A3(new_n507), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n504), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT85), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n219), .A2(G1698), .ZN(new_n511));
  OAI221_X1 g0311(.A(new_n511), .B1(G238), .B2(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G116), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n259), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT83), .ZN(new_n515));
  OAI21_X1  g0315(.A(G250), .B1(new_n478), .B2(new_n515), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n515), .B(G45), .C1(new_n255), .C2(new_n256), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n259), .ZN(new_n518));
  OAI21_X1  g0318(.A(KEYINPUT84), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n274), .B1(new_n478), .B2(new_n515), .ZN(new_n520));
  INV_X1    g0320(.A(G250), .ZN(new_n521));
  OAI21_X1  g0321(.A(G45), .B1(new_n255), .B2(new_n256), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n521), .B1(new_n522), .B2(KEYINPUT83), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT84), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n520), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n514), .B1(new_n519), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n478), .A2(G274), .A3(new_n259), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n391), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT19), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n306), .A2(new_n308), .A3(G97), .ZN(new_n530));
  AOI21_X1  g0330(.A(G20), .B1(new_n324), .B2(new_n325), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n529), .A2(new_n530), .B1(new_n531), .B2(G68), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n227), .B1(new_n267), .B2(new_n529), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(G87), .B2(new_n206), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n301), .ZN(new_n536));
  INV_X1    g0336(.A(new_n413), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n537), .A2(new_n292), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(G87), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n536), .B(new_n539), .C1(new_n540), .C2(new_n483), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n510), .B1(new_n528), .B2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n527), .ZN(new_n543));
  AOI211_X1 g0343(.A(new_n543), .B(new_n514), .C1(new_n519), .C2(new_n525), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n544), .A2(KEYINPUT86), .A3(G190), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n519), .A2(new_n525), .ZN(new_n546));
  INV_X1    g0346(.A(new_n514), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n546), .A2(G190), .A3(new_n527), .A4(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT86), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n305), .B1(new_n532), .B2(new_n534), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n483), .A2(new_n540), .ZN(new_n552));
  NOR3_X1   g0352(.A1(new_n551), .A2(new_n538), .A3(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(KEYINPUT85), .B(new_n553), .C1(new_n544), .C2(new_n391), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n542), .A2(new_n545), .A3(new_n550), .A4(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n546), .A2(new_n382), .A3(new_n527), .A4(new_n547), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n484), .A2(new_n537), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n536), .A2(new_n557), .A3(new_n539), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n556), .B(new_n558), .C1(new_n544), .C2(G169), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n227), .B(G87), .C1(new_n270), .C2(new_n271), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT22), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT22), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n403), .A2(new_n563), .A3(new_n227), .A4(G87), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT24), .ZN(new_n566));
  OR3_X1    g0366(.A1(new_n513), .A2(KEYINPUT90), .A3(G20), .ZN(new_n567));
  OAI21_X1  g0367(.A(KEYINPUT90), .B1(new_n513), .B2(G20), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT23), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n227), .B2(G107), .ZN(new_n570));
  INV_X1    g0370(.A(G107), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n571), .A2(KEYINPUT23), .A3(G20), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n567), .A2(new_n568), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n565), .A2(new_n566), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n566), .B1(new_n565), .B2(new_n573), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n301), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n484), .A2(G107), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n292), .A2(G107), .ZN(new_n578));
  XNOR2_X1  g0378(.A(new_n578), .B(KEYINPUT25), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(G250), .B(new_n438), .C1(new_n270), .C2(new_n271), .ZN(new_n581));
  OAI211_X1 g0381(.A(G257), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n582));
  NAND2_X1  g0382(.A1(G33), .A2(G294), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT91), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n581), .A2(new_n582), .A3(KEYINPUT91), .A4(new_n583), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n259), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AND2_X1   g0388(.A1(KEYINPUT5), .A2(G41), .ZN(new_n589));
  NOR2_X1   g0389(.A1(KEYINPUT5), .A2(G41), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(G264), .B(new_n259), .C1(new_n522), .C2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n283), .B1(new_n594), .B2(new_n479), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n592), .A2(KEYINPUT92), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT92), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n476), .A2(new_n597), .A3(G264), .A4(new_n259), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n479), .ZN(new_n600));
  NOR4_X1   g0400(.A1(new_n588), .A2(new_n599), .A3(new_n382), .A4(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n580), .B1(new_n595), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n586), .A2(new_n587), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n274), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n604), .A2(new_n479), .A3(new_n592), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n588), .A2(new_n599), .A3(new_n600), .ZN(new_n606));
  OAI22_X1  g0406(.A1(new_n605), .A2(G190), .B1(new_n606), .B2(G200), .ZN(new_n607));
  INV_X1    g0407(.A(new_n580), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(G107), .B1(new_n339), .B2(new_n340), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT6), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n487), .A2(new_n571), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n611), .B1(new_n612), .B2(new_n205), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n571), .A2(KEYINPUT6), .A3(G97), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G20), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n310), .A2(G77), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n610), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n301), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n292), .A2(G97), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n483), .A2(new_n487), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n619), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n476), .A2(G257), .A3(new_n259), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  OAI211_X1 g0426(.A(G244), .B(new_n438), .C1(new_n270), .C2(new_n271), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT4), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n627), .A2(new_n628), .B1(G33), .B2(G283), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n403), .A2(KEYINPUT4), .A3(G244), .A4(new_n438), .ZN(new_n630));
  OAI211_X1 g0430(.A(G250), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(KEYINPUT82), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT82), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n403), .A2(new_n633), .A3(G250), .A4(G1698), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n629), .A2(new_n630), .A3(new_n632), .A4(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n626), .B1(new_n635), .B2(new_n274), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n636), .A2(new_n382), .A3(new_n479), .ZN(new_n637));
  AOI211_X1 g0437(.A(new_n600), .B(new_n626), .C1(new_n274), .C2(new_n635), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n624), .B(new_n637), .C1(new_n638), .C2(G169), .ZN(new_n639));
  AOI211_X1 g0439(.A(new_n620), .B(new_n622), .C1(new_n618), .C2(new_n301), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n636), .A2(G190), .A3(new_n479), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n640), .B(new_n641), .C1(new_n638), .C2(new_n391), .ZN(new_n642));
  AND4_X1   g0442(.A1(new_n602), .A2(new_n609), .A3(new_n639), .A4(new_n642), .ZN(new_n643));
  AND4_X1   g0443(.A1(new_n461), .A2(new_n509), .A3(new_n560), .A4(new_n643), .ZN(G372));
  INV_X1    g0444(.A(new_n319), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n316), .B1(new_n427), .B2(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n399), .A2(new_n400), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n390), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n455), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n459), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT94), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI211_X1 g0452(.A(KEYINPUT94), .B(new_n459), .C1(new_n648), .C2(new_n649), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n602), .A2(KEYINPUT93), .ZN(new_n655));
  INV_X1    g0455(.A(new_n505), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT89), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n473), .A2(new_n480), .B1(new_n495), .B2(new_n485), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n657), .B1(new_n658), .B2(G169), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n502), .B1(new_n659), .B2(new_n498), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT93), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n661), .B(new_n580), .C1(new_n595), .C2(new_n601), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n655), .A2(new_n656), .A3(new_n660), .A4(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n642), .A2(new_n639), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n594), .A2(new_n408), .A3(new_n479), .ZN(new_n665));
  INV_X1    g0465(.A(new_n599), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n604), .A2(new_n666), .A3(new_n479), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n391), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n580), .B1(new_n665), .B2(new_n668), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n548), .B(new_n553), .C1(new_n544), .C2(new_n391), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n559), .A2(new_n670), .ZN(new_n671));
  NOR3_X1   g0471(.A1(new_n664), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n663), .A2(new_n672), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n636), .A2(new_n382), .A3(new_n479), .ZN(new_n674));
  AOI21_X1  g0474(.A(G169), .B1(new_n636), .B2(new_n479), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n676), .A2(new_n559), .A3(new_n624), .A4(new_n670), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n559), .B1(new_n677), .B2(KEYINPUT26), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n639), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n555), .A2(new_n559), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(KEYINPUT26), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n673), .A2(new_n679), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n461), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n654), .A2(new_n684), .ZN(G369));
  NAND2_X1  g0485(.A1(new_n660), .A2(new_n656), .ZN(new_n686));
  INV_X1    g0486(.A(G13), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(G20), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n474), .A2(new_n688), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n689), .A2(KEYINPUT27), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(KEYINPUT27), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(G213), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(G343), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(new_n496), .ZN(new_n695));
  MUX2_X1   g0495(.A(new_n686), .B(new_n509), .S(new_n695), .Z(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n602), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(new_n669), .ZN(new_n700));
  INV_X1    g0500(.A(new_n694), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n700), .B1(new_n608), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n699), .A2(new_n694), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n698), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n655), .A2(new_n662), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n701), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n694), .B1(new_n660), .B2(new_n656), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n700), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n705), .A2(new_n707), .A3(new_n709), .ZN(G399));
  INV_X1    g0510(.A(new_n209), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(G41), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G1), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n205), .A2(new_n540), .A3(new_n489), .ZN(new_n715));
  OAI22_X1  g0515(.A1(new_n714), .A2(new_n715), .B1(new_n230), .B2(new_n713), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT28), .ZN(new_n717));
  OR2_X1    g0517(.A1(new_n681), .A2(KEYINPUT26), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n672), .B1(new_n686), .B2(new_n699), .ZN(new_n719));
  INV_X1    g0519(.A(new_n559), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n720), .B1(new_n677), .B2(KEYINPUT26), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n718), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n701), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT29), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n678), .B1(new_n663), .B2(new_n672), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n694), .B1(new_n725), .B2(new_n682), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT29), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n604), .A2(new_n666), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n516), .A2(new_n518), .A3(KEYINPUT84), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n524), .B1(new_n520), .B2(new_n523), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n527), .B(new_n547), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT96), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n500), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n588), .A2(new_n599), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT96), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n544), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n734), .A2(new_n735), .A3(new_n638), .A4(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT30), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n733), .A2(KEYINPUT97), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n636), .A2(new_n479), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT97), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n526), .A2(new_n744), .A3(new_n527), .ZN(new_n745));
  AND3_X1   g0545(.A1(new_n742), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n746), .A2(new_n382), .A3(new_n481), .A4(new_n667), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n526), .A2(new_n604), .A3(new_n527), .A4(new_n666), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n500), .B1(new_n748), .B2(KEYINPUT96), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n749), .A2(KEYINPUT30), .A3(new_n638), .A4(new_n738), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n741), .A2(new_n747), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n694), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT31), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g0554(.A(KEYINPUT95), .B(KEYINPUT31), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n751), .A2(new_n694), .A3(new_n755), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n643), .A2(new_n560), .A3(new_n509), .A4(new_n701), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n754), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT98), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n758), .A2(new_n759), .A3(G330), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n759), .B1(new_n758), .B2(G330), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n729), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n717), .B1(new_n763), .B2(G1), .ZN(G364));
  OR2_X1    g0564(.A1(new_n696), .A2(G330), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n714), .B1(G45), .B2(new_n688), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n765), .A2(new_n697), .A3(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT99), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n226), .B1(G20), .B2(new_n283), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n227), .A2(new_n382), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G190), .A2(G200), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G311), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n272), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n393), .A2(new_n391), .A3(new_n773), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n393), .A2(G200), .A3(new_n773), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI22_X1  g0581(.A1(G322), .A2(new_n779), .B1(new_n781), .B2(G326), .ZN(new_n782));
  INV_X1    g0582(.A(G294), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G179), .A2(G200), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n227), .B1(new_n784), .B2(G190), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n227), .A2(G190), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n786), .A2(G179), .A3(G200), .ZN(new_n787));
  XOR2_X1   g0587(.A(KEYINPUT33), .B(G317), .Z(new_n788));
  OAI221_X1 g0588(.A(new_n782), .B1(new_n783), .B2(new_n785), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n786), .A2(new_n784), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n777), .B(new_n789), .C1(G329), .C2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G283), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n391), .A2(G179), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n786), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n794), .A2(G20), .A3(G190), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n792), .B1(new_n793), .B2(new_n795), .C1(new_n466), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n791), .A2(G159), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n798), .A2(KEYINPUT32), .B1(new_n778), .B2(new_n221), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n403), .B1(new_n796), .B2(new_n540), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT101), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n798), .A2(KEYINPUT32), .ZN(new_n802));
  INV_X1    g0602(.A(new_n785), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G97), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n201), .B2(new_n787), .ZN(new_n805));
  OR3_X1    g0605(.A1(new_n801), .A2(new_n802), .A3(new_n805), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n799), .B(new_n806), .C1(G50), .C2(new_n781), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n807), .B1(new_n202), .B2(new_n775), .C1(new_n571), .C2(new_n795), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n772), .B1(new_n797), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(G13), .A2(G33), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(G20), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n771), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n246), .A2(G45), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n711), .A2(new_n403), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n814), .B(new_n815), .C1(G45), .C2(new_n230), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n711), .A2(new_n272), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n817), .A2(G355), .B1(new_n489), .B2(new_n711), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT100), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n809), .B1(new_n813), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n812), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n821), .B(new_n766), .C1(new_n696), .C2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n768), .A2(new_n769), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n770), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT102), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(G396));
  INV_X1    g0627(.A(new_n418), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n416), .B1(new_n415), .B2(new_n417), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n694), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT105), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n424), .A2(KEYINPUT105), .A3(new_n694), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n832), .A2(new_n833), .A3(new_n422), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(new_n427), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n428), .A2(new_n701), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NOR3_X1   g0638(.A1(new_n761), .A2(new_n762), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n758), .A2(G330), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(KEYINPUT98), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n837), .B1(new_n841), .B2(new_n760), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  OR2_X1    g0643(.A1(new_n843), .A2(new_n726), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n726), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n844), .A2(new_n845), .A3(new_n767), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n780), .A2(new_n466), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n804), .B1(new_n489), .B2(new_n775), .C1(new_n776), .C2(new_n790), .ZN(new_n848));
  INV_X1    g0648(.A(new_n796), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n847), .B(new_n848), .C1(G107), .C2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n795), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(G87), .ZN(new_n852));
  INV_X1    g0652(.A(new_n787), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(G283), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n403), .B1(new_n779), .B2(G294), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n850), .A2(new_n852), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  XOR2_X1   g0656(.A(KEYINPUT103), .B(G143), .Z(new_n857));
  AOI22_X1  g0657(.A1(new_n779), .A2(new_n857), .B1(G150), .B2(new_n853), .ZN(new_n858));
  INV_X1    g0658(.A(G137), .ZN(new_n859));
  INV_X1    g0659(.A(G159), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n858), .B1(new_n859), .B2(new_n780), .C1(new_n860), .C2(new_n775), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT34), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n861), .A2(new_n862), .B1(G50), .B2(new_n849), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n863), .B1(new_n221), .B2(new_n785), .C1(new_n201), .C2(new_n795), .ZN(new_n864));
  INV_X1    g0664(.A(G132), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n403), .B1(new_n865), .B2(new_n790), .C1(new_n861), .C2(new_n862), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n856), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  XOR2_X1   g0667(.A(new_n867), .B(KEYINPUT104), .Z(new_n868));
  OAI221_X1 g0668(.A(new_n766), .B1(new_n811), .B2(new_n838), .C1(new_n868), .C2(new_n772), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n771), .A2(new_n810), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n869), .B1(new_n202), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n846), .A2(new_n872), .ZN(G384));
  NAND2_X1  g0673(.A1(new_n315), .A2(new_n694), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n316), .A2(new_n319), .A3(new_n874), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n315), .B(new_n694), .C1(new_n291), .C2(new_n645), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n683), .A2(new_n701), .A3(new_n835), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n878), .B1(new_n879), .B2(new_n836), .ZN(new_n880));
  INV_X1    g0680(.A(new_n692), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n344), .A2(new_n343), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n322), .B1(new_n882), .B2(new_n330), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n883), .A2(new_n301), .A3(new_n345), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n355), .A2(new_n356), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n881), .B(new_n886), .C1(new_n390), .C2(new_n401), .ZN(new_n887));
  INV_X1    g0687(.A(new_n397), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n386), .A2(new_n283), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n384), .B(new_n382), .C1(new_n378), .C2(new_n379), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n891), .A2(new_n692), .B1(new_n885), .B2(new_n884), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT37), .B1(new_n888), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n365), .A2(new_n387), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n365), .A2(new_n881), .ZN(new_n895));
  XOR2_X1   g0695(.A(KEYINPUT106), .B(KEYINPUT37), .Z(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n894), .A2(new_n895), .A3(new_n397), .A4(new_n897), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n893), .A2(new_n898), .A3(KEYINPUT107), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT107), .B1(new_n893), .B2(new_n898), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n887), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT38), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n887), .B(KEYINPUT38), .C1(new_n899), .C2(new_n900), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n880), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT18), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n894), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n365), .A2(new_n387), .A3(KEYINPUT18), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n910), .A2(new_n881), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n906), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT108), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT39), .ZN(new_n915));
  INV_X1    g0715(.A(new_n904), .ZN(new_n916));
  INV_X1    g0716(.A(new_n895), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n399), .A2(KEYINPUT109), .A3(new_n400), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n910), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT109), .B1(new_n399), .B2(new_n400), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n917), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n894), .A2(new_n895), .A3(new_n397), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n896), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n898), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT38), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n915), .B1(new_n916), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n316), .A2(new_n694), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n903), .A2(KEYINPUT39), .A3(new_n904), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT108), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n906), .A2(new_n930), .A3(new_n912), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n914), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT112), .ZN(new_n933));
  INV_X1    g0733(.A(new_n729), .ZN(new_n934));
  INV_X1    g0734(.A(new_n461), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n654), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n933), .B(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n916), .A2(new_n925), .ZN(new_n940));
  INV_X1    g0740(.A(new_n755), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n752), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n751), .A2(KEYINPUT31), .A3(new_n694), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n942), .A2(new_n757), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n837), .B1(new_n875), .B2(new_n876), .ZN(new_n945));
  AOI21_X1  g0745(.A(KEYINPUT110), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT40), .B1(new_n940), .B2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT40), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n903), .A2(new_n948), .A3(new_n904), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n757), .A2(new_n943), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n755), .B1(new_n751), .B2(new_n694), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n945), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT110), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(KEYINPUT40), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n949), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n947), .A2(new_n956), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT111), .Z(new_n958));
  NAND2_X1  g0758(.A1(new_n461), .A2(new_n944), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n958), .B(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(G330), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n939), .B(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n474), .B2(new_n688), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n489), .B1(new_n615), .B2(KEYINPUT35), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n964), .B(new_n229), .C1(KEYINPUT35), .C2(new_n615), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT36), .ZN(new_n966));
  OAI21_X1  g0766(.A(G77), .B1(new_n221), .B2(new_n201), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n967), .A2(new_n230), .B1(G50), .B2(new_n201), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n687), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n963), .B(new_n966), .C1(new_n474), .C2(new_n969), .ZN(G367));
  NAND2_X1  g0770(.A1(new_n851), .A2(G77), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n971), .B1(new_n217), .B2(new_n775), .C1(new_n859), .C2(new_n790), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n272), .B(new_n972), .C1(G159), .C2(new_n853), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n781), .A2(new_n857), .B1(G68), .B2(new_n803), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(G150), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n975), .B1(new_n221), .B2(new_n796), .C1(new_n976), .C2(new_n778), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n853), .A2(G294), .B1(new_n791), .B2(G317), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n978), .B1(new_n487), .B2(new_n795), .C1(new_n793), .C2(new_n775), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n849), .A2(KEYINPUT46), .A3(G116), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n803), .A2(G107), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(KEYINPUT46), .B1(new_n849), .B2(G116), .ZN(new_n983));
  NOR4_X1   g0783(.A1(new_n979), .A2(new_n403), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n984), .B1(new_n466), .B2(new_n778), .C1(new_n776), .C2(new_n780), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n977), .A2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT47), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n771), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n701), .A2(new_n553), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n720), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n671), .B2(new_n989), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n991), .A2(new_n822), .ZN(new_n992));
  INV_X1    g0792(.A(new_n815), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n813), .B1(new_n209), .B2(new_n413), .C1(new_n235), .C2(new_n993), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n988), .A2(new_n766), .A3(new_n992), .A4(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n263), .B1(new_n688), .B2(G45), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n642), .B(new_n639), .C1(new_n640), .C2(new_n701), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n680), .A2(new_n694), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(new_n709), .B2(new_n707), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT44), .Z(new_n1002));
  AOI21_X1  g0802(.A(new_n697), .B1(new_n702), .B2(new_n703), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n709), .A2(new_n707), .A3(new_n1000), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT45), .ZN(new_n1005));
  OR3_X1    g0805(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1003), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n709), .B1(new_n704), .B2(new_n708), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(new_n697), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n763), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n712), .B(KEYINPUT41), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n997), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1000), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n705), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n643), .A2(new_n708), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT42), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n639), .B1(new_n998), .B2(new_n602), .ZN(new_n1019));
  AND2_X1   g0819(.A1(new_n1019), .A2(new_n701), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1016), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1015), .A2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1015), .A2(new_n1021), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  OR3_X1    g0825(.A1(new_n1022), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1025), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n995), .B1(new_n1013), .B2(new_n1028), .ZN(G387));
  INV_X1    g0829(.A(G322), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n780), .A2(new_n1030), .B1(new_n776), .B2(new_n787), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT116), .ZN(new_n1032));
  INV_X1    g0832(.A(G317), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n778), .A2(new_n1033), .B1(new_n466), .B2(new_n775), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT115), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT48), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n803), .A2(G283), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n849), .A2(G294), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT117), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT49), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n1041), .A2(new_n1042), .B1(G326), .B2(new_n791), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n851), .A2(G116), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1043), .A2(new_n1044), .A3(new_n272), .A4(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n795), .A2(new_n487), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n778), .A2(new_n217), .B1(new_n348), .B2(new_n787), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n803), .A2(new_n537), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n849), .A2(G77), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1049), .A2(new_n403), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1047), .B(new_n1052), .C1(G150), .C2(new_n791), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1053), .B1(new_n201), .B2(new_n775), .C1(new_n860), .C2(new_n780), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT114), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n772), .B1(new_n1046), .B2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n348), .A2(G50), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT113), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT50), .ZN(new_n1059));
  NOR4_X1   g0859(.A1(new_n1059), .A2(G45), .A3(new_n241), .A4(new_n715), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n993), .B1(new_n239), .B2(G45), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n715), .B2(new_n817), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n1060), .A2(new_n1062), .B1(G107), .B2(new_n209), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1063), .A2(new_n813), .ZN(new_n1064));
  NOR3_X1   g0864(.A1(new_n1056), .A2(new_n767), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n702), .A2(new_n703), .A3(new_n812), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1010), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1065), .A2(new_n1066), .B1(new_n997), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n763), .A2(new_n1067), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n712), .B1(new_n763), .B2(new_n1067), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1068), .B1(new_n1070), .B2(new_n1071), .ZN(G393));
  NAND3_X1  g0872(.A1(new_n1006), .A2(new_n997), .A3(new_n1007), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n776), .A2(new_n778), .B1(new_n780), .B2(new_n1033), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT52), .Z(new_n1075));
  NOR2_X1   g0875(.A1(new_n795), .A2(new_n571), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n272), .B1(new_n785), .B2(new_n489), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n787), .A2(new_n466), .B1(new_n790), .B2(new_n1030), .ZN(new_n1078));
  NOR4_X1   g0878(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1079), .B1(new_n793), .B2(new_n796), .C1(new_n783), .C2(new_n775), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n217), .A2(new_n787), .B1(new_n775), .B2(new_n348), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT119), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1082), .A2(new_n272), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n1083), .B1(new_n201), .B2(new_n796), .C1(new_n202), .C2(new_n785), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n976), .A2(new_n780), .B1(new_n778), .B2(new_n860), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT118), .Z(new_n1086));
  OR2_X1    g0886(.A1(new_n1086), .A2(KEYINPUT51), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(KEYINPUT51), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n791), .A2(new_n857), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1087), .A2(new_n1088), .A3(new_n852), .A4(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1080), .B1(new_n1084), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n771), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1014), .A2(new_n812), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n813), .B1(new_n487), .B2(new_n209), .C1(new_n249), .C2(new_n993), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1092), .A2(new_n766), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1073), .A2(new_n1095), .ZN(new_n1096));
  OR2_X1    g0896(.A1(new_n1008), .A2(new_n1069), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n713), .B1(new_n1008), .B2(new_n1069), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1096), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(G390));
  NAND2_X1  g0900(.A1(new_n926), .A2(new_n928), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n927), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n836), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n726), .B2(new_n835), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1102), .B1(new_n1104), .B2(new_n878), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT109), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n401), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1108), .A2(new_n910), .A3(new_n918), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1109), .A2(new_n917), .B1(new_n898), .B2(new_n923), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n904), .B1(new_n1110), .B2(KEYINPUT38), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n722), .A2(new_n701), .A3(new_n835), .ZN(new_n1112));
  AND2_X1   g0912(.A1(new_n1112), .A2(new_n836), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1111), .B(new_n1102), .C1(new_n1113), .C2(new_n878), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n838), .B(new_n877), .C1(new_n761), .C2(new_n762), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n1106), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n944), .A2(G330), .A3(new_n945), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n1106), .B2(new_n1114), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n461), .A2(G330), .A3(new_n944), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n654), .B(new_n1120), .C1(new_n934), .C2(new_n935), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1117), .B1(new_n842), .B2(new_n877), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n879), .A2(new_n836), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n944), .A2(G330), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n878), .B1(new_n1125), .B2(new_n837), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1115), .A2(new_n1113), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1121), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT120), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1119), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1117), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n838), .B1(new_n761), .B2(new_n762), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1131), .B1(new_n1132), .B2(new_n878), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1127), .B1(new_n1133), .B2(new_n1104), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1121), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n880), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n1137), .A2(new_n1102), .B1(new_n926), .B2(new_n928), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1111), .A2(new_n1102), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1112), .A2(new_n836), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1139), .B1(new_n877), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1131), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1106), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1136), .A2(KEYINPUT120), .A3(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1130), .A2(new_n1145), .A3(new_n712), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1101), .A2(new_n810), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n870), .A2(new_n348), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n796), .A2(KEYINPUT53), .A3(new_n976), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n272), .B(new_n1149), .C1(G159), .C2(new_n803), .ZN(new_n1150));
  INV_X1    g0950(.A(G128), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n1150), .B1(new_n1151), .B2(new_n780), .C1(new_n865), .C2(new_n778), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n787), .A2(new_n859), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT54), .B(G143), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n775), .A2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(KEYINPUT53), .B1(new_n796), .B2(new_n976), .ZN(new_n1156));
  INV_X1    g0956(.A(G125), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1156), .B1(new_n217), .B2(new_n795), .C1(new_n1157), .C2(new_n790), .ZN(new_n1158));
  NOR4_X1   g0958(.A1(new_n1152), .A2(new_n1153), .A3(new_n1155), .A4(new_n1158), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n781), .A2(G283), .B1(G77), .B2(new_n803), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n1160), .B1(new_n487), .B2(new_n775), .C1(new_n489), .C2(new_n778), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n790), .A2(new_n783), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n787), .A2(new_n571), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n272), .B1(new_n795), .B2(new_n201), .C1(new_n540), .C2(new_n796), .ZN(new_n1164));
  NOR4_X1   g0964(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n771), .B1(new_n1159), .B2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1147), .A2(new_n766), .A3(new_n1148), .A4(new_n1166), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT121), .Z(new_n1168));
  NAND2_X1  g0968(.A1(new_n1119), .A2(new_n997), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1146), .A2(new_n1168), .A3(new_n1169), .ZN(G378));
  INV_X1    g0970(.A(KEYINPUT57), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1121), .B1(new_n1119), .B2(new_n1134), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n930), .B1(new_n906), .B2(new_n912), .ZN(new_n1173));
  AOI211_X1 g0973(.A(KEYINPUT108), .B(new_n911), .C1(new_n880), .C2(new_n905), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n929), .ZN(new_n1175));
  NOR3_X1   g0975(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  AND3_X1   g0976(.A1(new_n949), .A2(new_n953), .A3(new_n955), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n952), .A2(new_n954), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n948), .B1(new_n1178), .B2(new_n1111), .ZN(new_n1179));
  OAI21_X1  g0979(.A(G330), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n456), .A2(new_n881), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT55), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n455), .B2(new_n459), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n459), .ZN(new_n1185));
  AOI211_X1 g0985(.A(KEYINPUT55), .B(new_n1185), .C1(new_n452), .C2(new_n454), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1182), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n448), .B1(new_n447), .B2(new_n451), .ZN(new_n1188));
  NOR3_X1   g0988(.A1(new_n453), .A2(KEYINPUT10), .A3(new_n450), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n459), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(KEYINPUT55), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n455), .A2(new_n1183), .A3(new_n459), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1191), .A2(new_n1192), .A3(new_n1181), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n1187), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1194), .B1(new_n1187), .B2(new_n1193), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1180), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1197), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n957), .A2(G330), .A3(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1176), .A2(new_n1198), .A3(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1199), .B1(new_n957), .B2(G330), .ZN(new_n1202));
  INV_X1    g1002(.A(G330), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1203), .B(new_n1197), .C1(new_n947), .C2(new_n956), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n932), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1201), .A2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1171), .B1(new_n1172), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1125), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n877), .B1(new_n1208), .B2(new_n838), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n842), .B2(new_n877), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1113), .A2(new_n1210), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1135), .B1(new_n1211), .B2(new_n1144), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1212), .A2(KEYINPUT57), .A3(new_n1201), .A4(new_n1205), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1207), .A2(new_n1213), .A3(new_n712), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1201), .A2(new_n1205), .A3(new_n997), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1199), .A2(new_n810), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n217), .B1(new_n270), .B2(G41), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n796), .A2(new_n1154), .B1(new_n775), .B2(new_n859), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n780), .A2(new_n1157), .B1(new_n865), .B2(new_n787), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(G128), .C2(new_n779), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n976), .B2(new_n785), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1221), .A2(KEYINPUT59), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n851), .A2(G159), .ZN(new_n1223));
  AOI21_X1  g1023(.A(G41), .B1(new_n791), .B2(G124), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1222), .A2(new_n258), .A3(new_n1223), .A4(new_n1224), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1221), .A2(KEYINPUT59), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1217), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n252), .B1(new_n487), .B2(new_n787), .C1(new_n778), .C2(new_n571), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1051), .B1(new_n201), .B2(new_n785), .C1(new_n780), .C2(new_n489), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1228), .B(new_n1229), .C1(G283), .C2(new_n791), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n403), .B1(new_n851), .B2(G58), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1230), .B(new_n1231), .C1(new_n413), .C2(new_n775), .ZN(new_n1232));
  XOR2_X1   g1032(.A(new_n1232), .B(KEYINPUT58), .Z(new_n1233));
  OAI21_X1  g1033(.A(new_n771), .B1(new_n1227), .B2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n870), .A2(new_n217), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1216), .A2(new_n766), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1215), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1214), .A2(new_n1237), .ZN(G375));
  OAI211_X1 g1038(.A(new_n1121), .B(new_n1127), .C1(new_n1133), .C2(new_n1104), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT123), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1124), .A2(KEYINPUT123), .A3(new_n1121), .A4(new_n1127), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1243), .A2(new_n1012), .A3(new_n1136), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1244), .B(KEYINPUT124), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n878), .A2(new_n810), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n870), .A2(new_n201), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n779), .A2(G137), .B1(G159), .B2(new_n849), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n1248), .B1(new_n865), .B2(new_n780), .C1(new_n787), .C2(new_n1154), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n785), .A2(new_n217), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n790), .A2(new_n1151), .ZN(new_n1251));
  OAI221_X1 g1051(.A(new_n403), .B1(new_n795), .B2(new_n221), .C1(new_n976), .C2(new_n775), .ZN(new_n1252));
  NOR4_X1   g1052(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .A4(new_n1252), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n849), .A2(G97), .B1(new_n791), .B2(G303), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n403), .B1(new_n1254), .B2(KEYINPUT125), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1255), .B(new_n971), .C1(KEYINPUT125), .C2(new_n1254), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n1050), .B1(new_n489), .B2(new_n787), .C1(new_n778), .C2(new_n793), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n775), .A2(new_n571), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n780), .A2(new_n783), .ZN(new_n1259));
  NOR4_X1   g1059(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .A4(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n771), .B1(new_n1253), .B2(new_n1260), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1246), .A2(new_n766), .A3(new_n1247), .A4(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(new_n1211), .B2(new_n996), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1245), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(G381));
  NOR2_X1   g1065(.A1(G375), .A2(G378), .ZN(new_n1266));
  INV_X1    g1066(.A(G384), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1099), .B(new_n995), .C1(new_n1013), .C2(new_n1028), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n826), .B(new_n1068), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1264), .A2(new_n1266), .A3(new_n1267), .A4(new_n1270), .ZN(G407));
  INV_X1    g1071(.A(G213), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(new_n1266), .B2(new_n693), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(G407), .A2(new_n1273), .ZN(G409));
  INV_X1    g1074(.A(KEYINPUT60), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n712), .B1(new_n1239), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1136), .A2(KEYINPUT60), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1276), .B1(new_n1243), .B2(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1267), .B1(new_n1278), .B2(new_n1263), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1263), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n1241), .A2(new_n1242), .B1(new_n1136), .B2(KEYINPUT60), .ZN(new_n1281));
  OAI211_X1 g1081(.A(G384), .B(new_n1280), .C1(new_n1281), .C2(new_n1276), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1279), .A2(new_n1282), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1272), .A2(G343), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(G2897), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1283), .A2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1279), .A2(new_n1282), .A3(new_n1285), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(G378), .A2(new_n1214), .A3(new_n1237), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1212), .A2(new_n1012), .A3(new_n1201), .A4(new_n1205), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1237), .A2(new_n1291), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1292), .A2(new_n1168), .A3(new_n1169), .A4(new_n1146), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1284), .B1(new_n1290), .B2(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(KEYINPUT63), .B1(new_n1289), .B2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1284), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1279), .A2(new_n1282), .ZN(new_n1297));
  AND3_X1   g1097(.A1(G378), .A2(new_n1214), .A3(new_n1237), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1215), .A2(new_n1236), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1172), .A2(new_n1206), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1299), .B1(new_n1300), .B2(new_n1012), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(G378), .A2(new_n1301), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1296), .B(new_n1297), .C1(new_n1298), .C2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1295), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(G387), .A2(G390), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(G393), .A2(G396), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1269), .ZN(new_n1307));
  AND3_X1   g1107(.A1(new_n1305), .A2(new_n1307), .A3(new_n1268), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1307), .B1(new_n1305), .B2(new_n1268), .ZN(new_n1309));
  OR2_X1    g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1310), .A2(KEYINPUT61), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT63), .ZN(new_n1312));
  OAI21_X1  g1112(.A(KEYINPUT126), .B1(new_n1303), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT126), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1294), .A2(new_n1314), .A3(KEYINPUT63), .A4(new_n1297), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1304), .A2(new_n1311), .A3(new_n1313), .A4(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1303), .A2(KEYINPUT62), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1296), .B1(new_n1298), .B2(new_n1302), .ZN(new_n1318));
  AND3_X1   g1118(.A1(new_n1279), .A2(new_n1282), .A3(new_n1285), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1285), .B1(new_n1279), .B2(new_n1282), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1318), .A2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT61), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT62), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1294), .A2(new_n1324), .A3(new_n1297), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1317), .A2(new_n1322), .A3(new_n1323), .A4(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n1310), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1316), .A2(new_n1327), .ZN(G405));
  INV_X1    g1128(.A(G378), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(G375), .A2(new_n1329), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(new_n1297), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1332), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1298), .A2(KEYINPUT127), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1331), .A2(new_n1297), .ZN(new_n1335));
  NOR3_X1   g1135(.A1(new_n1333), .A2(new_n1334), .A3(new_n1335), .ZN(new_n1336));
  OR2_X1    g1136(.A1(new_n1298), .A2(KEYINPUT127), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1310), .A2(new_n1283), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1337), .B1(new_n1338), .B2(new_n1332), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1330), .B1(new_n1336), .B2(new_n1339), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1334), .B1(new_n1333), .B2(new_n1335), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1338), .A2(new_n1337), .A3(new_n1332), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1341), .A2(new_n1329), .A3(G375), .A4(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1340), .A2(new_n1343), .ZN(G402));
endmodule


