//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n777, new_n778,
    new_n779, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G227), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n193), .B(KEYINPUT78), .ZN(new_n194));
  XNOR2_X1  g008(.A(G110), .B(G140), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n194), .B(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G134), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT11), .B1(new_n198), .B2(G137), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT11), .ZN(new_n200));
  INV_X1    g014(.A(G137), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(G134), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT65), .B1(new_n201), .B2(G134), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(new_n198), .A3(G137), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT66), .A2(G131), .ZN(new_n207));
  AND4_X1   g021(.A1(new_n203), .A2(new_n204), .A3(new_n206), .A4(new_n207), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n204), .A2(new_n206), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n207), .B1(new_n209), .B2(new_n203), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G143), .ZN(new_n213));
  INV_X1    g027(.A(G143), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G146), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT1), .B1(new_n214), .B2(G146), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(G128), .A3(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G128), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n213), .B(new_n215), .C1(KEYINPUT1), .C2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G104), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G107), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT81), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n222), .A2(G107), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(G101), .B1(new_n223), .B2(KEYINPUT81), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G101), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n230));
  AOI22_X1  g044(.A1(KEYINPUT79), .A2(new_n230), .B1(new_n222), .B2(G107), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT79), .ZN(new_n232));
  INV_X1    g046(.A(G107), .ZN(new_n233));
  AND4_X1   g047(.A1(new_n232), .A2(new_n233), .A3(KEYINPUT3), .A4(G104), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n232), .A2(KEYINPUT3), .B1(new_n233), .B2(G104), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n229), .B(new_n231), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT80), .ZN(new_n237));
  OAI22_X1  g051(.A1(KEYINPUT79), .A2(new_n230), .B1(new_n222), .B2(G107), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n232), .A2(new_n233), .A3(KEYINPUT3), .A4(G104), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT80), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n240), .A2(new_n241), .A3(new_n229), .A4(new_n231), .ZN(new_n242));
  AOI211_X1 g056(.A(new_n221), .B(new_n228), .C1(new_n237), .C2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n237), .A2(new_n242), .ZN(new_n244));
  OAI22_X1  g058(.A1(new_n232), .A2(KEYINPUT3), .B1(new_n233), .B2(G104), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n245), .B1(new_n238), .B2(new_n239), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT4), .B1(new_n246), .B2(new_n229), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(KEYINPUT0), .A2(G128), .ZN(new_n250));
  OR2_X1    g064(.A1(KEYINPUT0), .A2(G128), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n216), .A2(KEYINPUT64), .A3(new_n250), .A4(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n250), .ZN(new_n253));
  XNOR2_X1  g067(.A(G143), .B(G146), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT64), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n240), .A2(new_n231), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(new_n259), .A3(G101), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  AOI22_X1  g075(.A1(new_n243), .A2(KEYINPUT10), .B1(new_n249), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT82), .ZN(new_n263));
  NOR3_X1   g077(.A1(new_n243), .A2(new_n263), .A3(KEYINPUT10), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n218), .A2(new_n220), .ZN(new_n265));
  INV_X1    g079(.A(new_n228), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n244), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT10), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT82), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n211), .B(new_n262), .C1(new_n264), .C2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n263), .B1(new_n243), .B2(KEYINPUT10), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n267), .A2(KEYINPUT82), .A3(new_n268), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n211), .B1(new_n274), .B2(new_n262), .ZN(new_n275));
  OAI211_X1 g089(.A(KEYINPUT83), .B(new_n197), .C1(new_n271), .C2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n211), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n228), .B1(new_n237), .B2(new_n242), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n278), .A2(new_n265), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n277), .B1(new_n279), .B2(new_n243), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT12), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT12), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n282), .B(new_n277), .C1(new_n279), .C2(new_n243), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n270), .A2(new_n196), .A3(new_n281), .A4(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n276), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n262), .B1(new_n264), .B2(new_n269), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n277), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n270), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT83), .B1(new_n288), .B2(new_n197), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n190), .B(new_n191), .C1(new_n285), .C2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n281), .A2(new_n283), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n197), .B1(new_n271), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n287), .A2(new_n196), .A3(new_n270), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(G469), .A3(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n190), .A2(new_n191), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n189), .B1(new_n290), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(G214), .B1(G237), .B2(G902), .ZN(new_n299));
  INV_X1    g113(.A(G119), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G116), .ZN(new_n301));
  INV_X1    g115(.A(G116), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G119), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT2), .B(G113), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n304), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT84), .B(KEYINPUT5), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G113), .ZN(new_n310));
  AND2_X1   g124(.A1(KEYINPUT84), .A2(KEYINPUT5), .ZN(new_n311));
  NOR2_X1   g125(.A1(KEYINPUT84), .A2(KEYINPUT5), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n301), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n310), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n306), .B1(new_n309), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n241), .B1(new_n246), .B2(new_n229), .ZN(new_n317));
  AND4_X1   g131(.A1(new_n241), .A2(new_n240), .A3(new_n229), .A4(new_n231), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n316), .B(new_n266), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n247), .B1(new_n242), .B2(new_n237), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n304), .B(new_n305), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n260), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n319), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(G110), .B(G122), .ZN(new_n324));
  OR2_X1    g138(.A1(new_n324), .A2(KEYINPUT85), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(KEYINPUT85), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n319), .B(new_n327), .C1(new_n320), .C2(new_n322), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(KEYINPUT6), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT6), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n323), .A2(new_n332), .A3(new_n328), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n252), .A2(new_n256), .A3(G125), .ZN(new_n334));
  INV_X1    g148(.A(G125), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n218), .A2(new_n335), .A3(new_n220), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n192), .A2(G224), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(KEYINPUT86), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n337), .B(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n331), .A2(new_n333), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(KEYINPUT7), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n334), .A2(new_n336), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n342), .B1(new_n334), .B2(new_n336), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(G113), .B1(new_n308), .B2(new_n301), .ZN(new_n346));
  AND3_X1   g160(.A1(new_n301), .A2(new_n303), .A3(KEYINPUT5), .ZN(new_n347));
  OAI22_X1  g161(.A1(new_n346), .A2(new_n347), .B1(new_n304), .B2(new_n305), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n266), .B(new_n348), .C1(new_n317), .C2(new_n318), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n325), .A2(KEYINPUT8), .A3(new_n326), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT8), .B1(new_n325), .B2(new_n326), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n316), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n278), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n345), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT87), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI211_X1 g172(.A(KEYINPUT87), .B(new_n345), .C1(new_n353), .C2(new_n355), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n330), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n341), .A2(new_n360), .A3(new_n191), .ZN(new_n361));
  OAI21_X1  g175(.A(G210), .B1(G237), .B2(G902), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n341), .A2(new_n360), .A3(new_n191), .A4(new_n362), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n192), .A2(G952), .ZN(new_n367));
  NAND2_X1  g181(.A1(G234), .A2(G237), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(G902), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n371), .A2(new_n192), .ZN(new_n372));
  XNOR2_X1  g186(.A(KEYINPUT21), .B(G898), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n370), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G217), .ZN(new_n376));
  NOR3_X1   g190(.A1(new_n187), .A2(new_n376), .A3(G953), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT13), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT91), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT91), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT13), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n214), .A2(G128), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT92), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n386), .B1(new_n214), .B2(G128), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n219), .A2(KEYINPUT92), .A3(G143), .ZN(new_n388));
  AOI22_X1  g202(.A1(new_n383), .A2(new_n385), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n384), .A2(new_n380), .A3(new_n382), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n198), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n387), .A2(new_n388), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(new_n198), .A3(new_n384), .ZN(new_n393));
  INV_X1    g207(.A(G122), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G116), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n302), .A2(G122), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n233), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n395), .A2(new_n396), .A3(G107), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n393), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n391), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n395), .A2(KEYINPUT14), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n397), .A2(new_n402), .A3(G107), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n395), .B(new_n396), .C1(KEYINPUT14), .C2(new_n233), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n198), .B1(new_n392), .B2(new_n384), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n405), .B1(new_n407), .B2(new_n393), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n378), .B1(new_n401), .B2(new_n408), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n393), .A2(new_n399), .A3(new_n398), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n383), .A2(new_n385), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(new_n390), .A3(new_n392), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G134), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n393), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n404), .B(new_n403), .C1(new_n415), .C2(new_n406), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(new_n416), .A3(new_n377), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n409), .A2(new_n417), .A3(KEYINPUT93), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT94), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT93), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n420), .B(new_n378), .C1(new_n401), .C2(new_n408), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n418), .A2(new_n419), .A3(new_n191), .A4(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G478), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(KEYINPUT15), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n422), .B(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(G140), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G125), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n335), .A2(G140), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT74), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n426), .A2(KEYINPUT74), .A3(G125), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n430), .A2(KEYINPUT16), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT16), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n427), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G146), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n432), .A2(new_n212), .A3(new_n434), .ZN(new_n437));
  NOR2_X1   g251(.A1(G237), .A2(G953), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n438), .A2(G143), .A3(G214), .ZN(new_n439));
  AOI21_X1  g253(.A(G143), .B1(new_n438), .B2(G214), .ZN(new_n440));
  OAI211_X1 g254(.A(KEYINPUT17), .B(G131), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G131), .B1(new_n439), .B2(new_n440), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT17), .ZN(new_n443));
  INV_X1    g257(.A(G237), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(new_n192), .A3(G214), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n214), .ZN(new_n446));
  INV_X1    g260(.A(G131), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n438), .A2(G143), .A3(G214), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n442), .A2(new_n443), .A3(new_n449), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n436), .A2(new_n437), .A3(new_n441), .A4(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(G113), .B(G122), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(new_n222), .ZN(new_n453));
  OAI211_X1 g267(.A(KEYINPUT18), .B(G131), .C1(new_n439), .C2(new_n440), .ZN(new_n454));
  NAND2_X1  g268(.A1(KEYINPUT18), .A2(G131), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n446), .A2(new_n448), .A3(new_n455), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n430), .A2(G146), .A3(new_n431), .ZN(new_n458));
  XNOR2_X1  g272(.A(G125), .B(G140), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n212), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n451), .A2(new_n453), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n453), .B1(new_n451), .B2(new_n462), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n191), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT90), .B(G475), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n451), .A2(new_n453), .A3(new_n462), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n430), .A2(KEYINPUT19), .A3(new_n431), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT88), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT19), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n471), .B1(new_n459), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n430), .A2(new_n471), .A3(KEYINPUT19), .A4(new_n431), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n212), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n435), .A2(G146), .B1(new_n442), .B2(new_n449), .ZN(new_n478));
  AOI22_X1  g292(.A1(new_n477), .A2(new_n478), .B1(new_n461), .B2(new_n457), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n469), .B1(new_n479), .B2(new_n453), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT20), .ZN(new_n481));
  NOR2_X1   g295(.A1(G475), .A2(G902), .ZN(new_n482));
  XOR2_X1   g296(.A(new_n482), .B(KEYINPUT89), .Z(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n480), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n481), .B1(new_n480), .B2(new_n484), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n468), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n425), .A2(new_n487), .ZN(new_n488));
  AND4_X1   g302(.A1(new_n299), .A2(new_n366), .A3(new_n375), .A4(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n257), .B1(new_n210), .B2(new_n208), .ZN(new_n490));
  AOI21_X1  g304(.A(G131), .B1(new_n209), .B2(new_n203), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n198), .A2(G137), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n201), .A2(G134), .ZN(new_n493));
  NOR3_X1   g307(.A1(new_n492), .A2(new_n493), .A3(new_n447), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n265), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n321), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n490), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT28), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(KEYINPUT71), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(KEYINPUT71), .B1(new_n497), .B2(new_n498), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n252), .A2(new_n256), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n200), .B1(G134), .B2(new_n201), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n198), .A2(KEYINPUT11), .A3(G137), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n204), .B(new_n206), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(KEYINPUT66), .A3(G131), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n209), .A2(new_n203), .A3(new_n207), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n503), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n504), .A2(new_n505), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n204), .A2(new_n206), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n447), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n494), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n221), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n509), .A2(new_n514), .A3(new_n321), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n496), .B1(new_n490), .B2(new_n495), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT28), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT70), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT70), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n519), .B(KEYINPUT28), .C1(new_n515), .C2(new_n516), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n438), .A2(G210), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n521), .B(KEYINPUT27), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT26), .B(G101), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n522), .B(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT29), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n502), .A2(new_n518), .A3(new_n520), .A4(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT72), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n497), .A2(new_n498), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT71), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n520), .A2(new_n499), .A3(new_n533), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n534), .A2(KEYINPUT72), .A3(new_n518), .A4(new_n527), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT67), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n537), .B1(new_n491), .B2(new_n494), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n512), .A2(KEYINPUT67), .A3(new_n513), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(new_n539), .A3(new_n265), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n496), .B1(new_n540), .B2(new_n490), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n536), .B1(new_n541), .B2(new_n515), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n542), .A2(new_n524), .A3(new_n531), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT30), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n494), .B1(new_n506), .B2(new_n447), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n265), .B1(new_n545), .B2(KEYINPUT67), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n491), .A2(new_n537), .A3(new_n494), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n544), .B(new_n490), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT30), .B1(new_n509), .B2(new_n514), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n496), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n525), .B1(new_n550), .B2(new_n515), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n543), .A2(new_n551), .A3(new_n526), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n530), .A2(new_n535), .A3(new_n191), .A4(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(G472), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT31), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n548), .A2(new_n549), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n515), .B1(new_n556), .B2(new_n321), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n555), .B1(new_n557), .B2(new_n524), .ZN(new_n558));
  XNOR2_X1  g372(.A(KEYINPUT68), .B(KEYINPUT31), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NOR4_X1   g374(.A1(new_n550), .A2(new_n525), .A3(new_n515), .A4(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n524), .B1(new_n542), .B2(new_n531), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n558), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(G472), .A2(G902), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n563), .A2(KEYINPUT32), .A3(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT32), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n556), .A2(new_n321), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n568), .A2(new_n524), .A3(new_n497), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT31), .ZN(new_n570));
  INV_X1    g384(.A(new_n562), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n568), .A2(new_n524), .A3(new_n497), .A4(new_n559), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n567), .B1(new_n573), .B2(new_n564), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n554), .B1(new_n566), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n192), .A2(G221), .A3(G234), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(KEYINPUT76), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT22), .B(G137), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n300), .A2(G128), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT23), .B1(new_n580), .B2(KEYINPUT73), .ZN(new_n581));
  AOI21_X1  g395(.A(KEYINPUT73), .B1(new_n219), .B2(G119), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT23), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(G110), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n300), .A2(G128), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n581), .A2(new_n584), .A3(new_n585), .A4(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(G119), .B(G128), .ZN(new_n588));
  XOR2_X1   g402(.A(KEYINPUT24), .B(G110), .Z(new_n589));
  OAI21_X1  g403(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n436), .A2(new_n590), .A3(new_n460), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT75), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n460), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n594), .B1(new_n435), .B2(G146), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n595), .A2(KEYINPUT75), .A3(new_n590), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n586), .B1(new_n582), .B2(new_n583), .ZN(new_n598));
  AOI211_X1 g412(.A(KEYINPUT73), .B(KEYINPUT23), .C1(new_n219), .C2(G119), .ZN(new_n599));
  OAI21_X1  g413(.A(G110), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n589), .A2(new_n588), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n602), .B1(new_n436), .B2(new_n437), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n579), .B1(new_n597), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n579), .ZN(new_n606));
  AOI211_X1 g420(.A(new_n606), .B(new_n603), .C1(new_n593), .C2(new_n596), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n376), .B1(G234), .B2(new_n191), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n610), .A2(G902), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n595), .A2(KEYINPUT75), .A3(new_n590), .ZN(new_n613));
  AOI21_X1  g427(.A(KEYINPUT75), .B1(new_n595), .B2(new_n590), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n604), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n606), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n597), .A2(new_n604), .A3(new_n579), .ZN(new_n617));
  AOI21_X1  g431(.A(G902), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(KEYINPUT77), .B1(new_n618), .B2(KEYINPUT25), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n191), .B1(new_n605), .B2(new_n607), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT25), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n620), .A2(new_n621), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n610), .B1(new_n624), .B2(KEYINPUT77), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n612), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n298), .A2(new_n489), .A3(new_n575), .A4(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G101), .ZN(G3));
  NOR3_X1   g443(.A1(new_n550), .A2(new_n525), .A3(new_n515), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n572), .B1(new_n630), .B2(new_n555), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n191), .B1(new_n631), .B2(new_n562), .ZN(new_n632));
  AOI22_X1  g446(.A1(new_n632), .A2(G472), .B1(new_n564), .B2(new_n573), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n298), .A2(new_n627), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT95), .ZN(new_n635));
  INV_X1    g449(.A(new_n299), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n636), .B1(new_n364), .B2(new_n365), .ZN(new_n637));
  INV_X1    g451(.A(new_n487), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT33), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n418), .A2(new_n639), .A3(new_n421), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n409), .A2(new_n417), .A3(KEYINPUT33), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n423), .A2(G902), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n418), .A2(new_n191), .A3(new_n421), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n423), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT96), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n643), .A2(KEYINPUT96), .A3(new_n645), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n638), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AND3_X1   g464(.A1(new_n637), .A2(new_n375), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n635), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT34), .B(G104), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G6));
  AOI211_X1 g468(.A(new_n636), .B(new_n374), .C1(new_n364), .C2(new_n365), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT97), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n656), .B1(new_n485), .B2(new_n486), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n477), .A2(new_n478), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n453), .B1(new_n658), .B2(new_n462), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n484), .B1(new_n659), .B2(new_n463), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(KEYINPUT20), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n480), .A2(new_n481), .A3(new_n484), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n661), .A2(KEYINPUT97), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n657), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n468), .ZN(new_n665));
  OR2_X1    g479(.A1(new_n422), .A2(new_n424), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n422), .A2(new_n424), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(KEYINPUT98), .B1(new_n655), .B2(new_n669), .ZN(new_n670));
  AND4_X1   g484(.A1(KEYINPUT98), .A2(new_n637), .A3(new_n669), .A4(new_n375), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n635), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT35), .B(G107), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G9));
  NOR2_X1   g490(.A1(new_n579), .A2(KEYINPUT36), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n615), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n611), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n679), .B1(new_n623), .B2(new_n625), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n298), .A2(new_n489), .A3(new_n633), .A4(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT37), .B(G110), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G12));
  NOR3_X1   g497(.A1(new_n371), .A2(G900), .A3(new_n192), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n370), .B1(KEYINPUT99), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n685), .B1(KEYINPUT99), .B2(new_n684), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n664), .A2(new_n668), .A3(new_n686), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n687), .A2(new_n637), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n298), .A2(new_n688), .A3(new_n575), .A4(new_n680), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT100), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n610), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n618), .A2(KEYINPUT25), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT77), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n618), .A2(KEYINPUT25), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n624), .A2(new_n696), .A3(KEYINPUT77), .ZN(new_n697));
  AOI22_X1  g511(.A1(new_n695), .A2(new_n697), .B1(new_n611), .B2(new_n678), .ZN(new_n698));
  OAI21_X1  g512(.A(KEYINPUT32), .B1(new_n563), .B2(new_n565), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n573), .A2(new_n567), .A3(new_n564), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n698), .B1(new_n701), .B2(new_n554), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n702), .A2(KEYINPUT100), .A3(new_n298), .A4(new_n688), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n691), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G128), .ZN(G30));
  INV_X1    g519(.A(KEYINPUT38), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n366), .B(new_n706), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n425), .A2(new_n299), .A3(new_n487), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n698), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n557), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n524), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n321), .B1(new_n509), .B2(new_n514), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n497), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n191), .B1(new_n715), .B2(new_n524), .ZN(new_n716));
  OAI21_X1  g530(.A(G472), .B1(new_n713), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n701), .A2(new_n717), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n718), .A2(KEYINPUT101), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n718), .A2(KEYINPUT101), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n710), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT102), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g537(.A(KEYINPUT103), .B(KEYINPUT39), .Z(new_n724));
  XNOR2_X1  g538(.A(new_n686), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n298), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT40), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(new_n728));
  OAI211_X1 g542(.A(KEYINPUT102), .B(new_n710), .C1(new_n719), .C2(new_n720), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n723), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G143), .ZN(G45));
  AND3_X1   g545(.A1(new_n643), .A2(KEYINPUT96), .A3(new_n645), .ZN(new_n732));
  AOI21_X1  g546(.A(KEYINPUT96), .B1(new_n643), .B2(new_n645), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n487), .B(new_n686), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n735), .A2(KEYINPUT104), .A3(new_n637), .ZN(new_n736));
  AOI21_X1  g550(.A(KEYINPUT104), .B1(new_n735), .B2(new_n637), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n702), .B(new_n298), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G146), .ZN(G48));
  INV_X1    g553(.A(new_n290), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n197), .B1(new_n271), .B2(new_n275), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT83), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n284), .A3(new_n276), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n190), .B1(new_n744), .B2(new_n191), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n740), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n626), .B1(new_n701), .B2(new_n554), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n746), .A2(new_n747), .A3(new_n188), .A4(new_n651), .ZN(new_n748));
  XNOR2_X1  g562(.A(KEYINPUT41), .B(G113), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(G15));
  NAND3_X1  g564(.A1(new_n746), .A2(new_n747), .A3(new_n188), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(new_n672), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n302), .ZN(G18));
  NAND4_X1  g567(.A1(new_n575), .A2(new_n375), .A3(new_n488), .A4(new_n680), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n191), .B1(new_n285), .B2(new_n289), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(G469), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n756), .A2(new_n637), .A3(new_n188), .A4(new_n290), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(new_n300), .ZN(G21));
  NAND2_X1  g573(.A1(new_n366), .A2(new_n708), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT105), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT105), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n366), .A2(new_n708), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n632), .A2(G472), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n520), .A2(new_n499), .A3(new_n533), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n519), .B1(new_n715), .B2(KEYINPUT28), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n525), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(new_n570), .A3(new_n572), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n564), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n765), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(new_n626), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n764), .A2(new_n375), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n746), .A2(new_n188), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(new_n394), .ZN(G24));
  AOI22_X1  g590(.A1(new_n632), .A2(G472), .B1(new_n564), .B2(new_n769), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n777), .A2(new_n680), .A3(new_n735), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n746), .A2(new_n778), .A3(new_n637), .A4(new_n188), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G125), .ZN(G27));
  INV_X1    g594(.A(KEYINPUT107), .ZN(new_n781));
  AOI22_X1  g595(.A1(new_n701), .A2(new_n781), .B1(G472), .B2(new_n553), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n699), .A2(KEYINPUT107), .A3(new_n700), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n626), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n292), .A2(new_n293), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT106), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n293), .A2(KEYINPUT106), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n290), .B(new_n296), .C1(new_n789), .C2(new_n190), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n366), .A2(new_n636), .A3(new_n189), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT42), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n734), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n784), .A2(new_n790), .A3(new_n791), .A4(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n747), .A2(new_n790), .A3(new_n791), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n792), .B1(new_n795), .B2(new_n734), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G131), .ZN(G33));
  NAND4_X1  g612(.A1(new_n747), .A2(new_n790), .A3(new_n687), .A4(new_n791), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G134), .ZN(G36));
  NAND3_X1  g614(.A1(new_n787), .A2(KEYINPUT45), .A3(new_n788), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT45), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n190), .B1(new_n785), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n295), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n804), .A2(KEYINPUT46), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(KEYINPUT46), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(new_n290), .A3(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n807), .A2(new_n188), .A3(new_n725), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT108), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n807), .A2(KEYINPUT108), .A3(new_n188), .A4(new_n725), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT44), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n633), .A2(new_n698), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n638), .B1(new_n732), .B2(new_n733), .ZN(new_n814));
  OR2_X1    g628(.A1(new_n814), .A2(KEYINPUT43), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(KEYINPUT43), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n812), .B1(new_n813), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n364), .A2(new_n299), .A3(new_n365), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n813), .A2(new_n817), .A3(new_n812), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n810), .A2(new_n811), .A3(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(G137), .ZN(G39));
  NAND3_X1  g639(.A1(new_n820), .A2(new_n626), .A3(new_n735), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n826), .A2(new_n575), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n807), .A2(KEYINPUT47), .A3(new_n188), .ZN(new_n829));
  INV_X1    g643(.A(new_n806), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n290), .B1(new_n804), .B2(KEYINPUT46), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n188), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT47), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n828), .B1(new_n829), .B2(new_n834), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(new_n426), .ZN(G42));
  XNOR2_X1  g650(.A(new_n746), .B(KEYINPUT110), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  OR2_X1    g652(.A1(new_n838), .A2(KEYINPUT49), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n719), .A2(new_n720), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n838), .A2(KEYINPUT49), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n627), .A2(new_n299), .A3(new_n188), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT109), .ZN(new_n843));
  INV_X1    g657(.A(new_n814), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n843), .A2(new_n707), .A3(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n839), .A2(new_n840), .A3(new_n841), .A4(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n691), .A2(new_n703), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT52), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n686), .A2(new_n188), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n679), .B(new_n850), .C1(new_n623), .C2(new_n625), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n851), .B1(new_n701), .B2(new_n717), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n852), .A2(new_n764), .A3(new_n790), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n779), .A2(new_n738), .A3(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n848), .A2(new_n849), .A3(new_n854), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n779), .A2(new_n738), .A3(new_n853), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT52), .B1(new_n856), .B2(new_n704), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n468), .A2(new_n686), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n664), .A2(new_n666), .A3(new_n667), .A4(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(new_n820), .A3(KEYINPUT112), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT112), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n863), .B1(new_n860), .B2(new_n819), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n702), .A2(new_n298), .A3(new_n862), .A4(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n778), .A2(new_n790), .A3(new_n791), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n865), .A2(new_n799), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n867), .B1(new_n794), .B2(new_n796), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n366), .A2(new_n299), .A3(new_n375), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n648), .A2(new_n487), .A3(new_n649), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n870), .B1(new_n487), .B2(new_n425), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n872), .A2(new_n298), .A3(new_n627), .A4(new_n633), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n873), .A2(new_n628), .A3(new_n681), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT111), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n873), .A2(new_n628), .A3(new_n681), .A4(KEYINPUT111), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI22_X1  g692(.A1(new_n773), .A2(new_n774), .B1(new_n757), .B2(new_n754), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n748), .B1(new_n751), .B2(new_n672), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n868), .A2(new_n878), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n847), .B1(new_n858), .B2(new_n882), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n868), .A2(new_n878), .A3(new_n881), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n849), .B1(new_n848), .B2(new_n854), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n856), .A2(KEYINPUT52), .A3(new_n704), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n884), .A2(KEYINPUT53), .A3(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n883), .A2(KEYINPUT54), .A3(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT54), .B1(new_n883), .B2(new_n888), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n774), .A2(new_n819), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT114), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n894), .B1(new_n817), .B2(new_n369), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n815), .A2(KEYINPUT114), .A3(new_n370), .A4(new_n816), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n893), .A2(new_n897), .A3(new_n784), .ZN(new_n898));
  XNOR2_X1  g712(.A(KEYINPUT117), .B(KEYINPUT48), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n772), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n901), .B1(new_n895), .B2(new_n896), .ZN(new_n902));
  INV_X1    g716(.A(new_n757), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT116), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n900), .A2(new_n904), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n902), .A2(new_n903), .ZN(new_n906));
  AOI22_X1  g720(.A1(new_n906), .A2(KEYINPUT116), .B1(new_n898), .B2(new_n899), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n626), .A2(new_n369), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n893), .A2(new_n840), .A3(new_n650), .A4(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n905), .A2(new_n907), .A3(new_n909), .A4(new_n367), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n829), .A2(new_n834), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n838), .A2(new_n188), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n820), .B(new_n902), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  AND4_X1   g727(.A1(new_n636), .A2(new_n746), .A3(new_n188), .A4(new_n707), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n902), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(KEYINPUT50), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n893), .A2(new_n897), .A3(new_n680), .A4(new_n777), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n732), .A2(new_n733), .A3(new_n487), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n893), .A2(new_n840), .A3(new_n908), .A4(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT50), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n902), .A2(new_n914), .A3(new_n920), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n916), .A2(new_n917), .A3(new_n919), .A4(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT51), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n910), .B1(new_n913), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n922), .A2(KEYINPUT115), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n917), .A2(new_n919), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT115), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n927), .A2(new_n928), .A3(new_n916), .A4(new_n921), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n926), .A2(new_n929), .A3(new_n913), .ZN(new_n930));
  XOR2_X1   g744(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n931));
  OAI21_X1  g745(.A(new_n925), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n892), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(G952), .A2(G953), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n846), .B1(new_n933), .B2(new_n934), .ZN(G75));
  NAND2_X1  g749(.A1(new_n883), .A2(new_n888), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n936), .A2(G210), .A3(G902), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n331), .A2(new_n333), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(new_n340), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT55), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT118), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n941), .A2(KEYINPUT56), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n937), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n940), .B1(new_n937), .B2(new_n942), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n192), .A2(G952), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(G51));
  INV_X1    g760(.A(KEYINPUT54), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n936), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n295), .B(KEYINPUT57), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n948), .A2(new_n889), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n744), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n191), .B1(new_n883), .B2(new_n888), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n952), .A2(new_n801), .A3(new_n803), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n945), .B1(new_n951), .B2(new_n953), .ZN(G54));
  INV_X1    g768(.A(new_n945), .ZN(new_n955));
  NAND2_X1  g769(.A1(KEYINPUT58), .A2(G475), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT119), .Z(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  AOI211_X1 g772(.A(new_n191), .B(new_n958), .C1(new_n883), .C2(new_n888), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n955), .B1(new_n959), .B2(new_n480), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT120), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n959), .A2(new_n961), .A3(new_n480), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n952), .A2(new_n480), .A3(new_n957), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(KEYINPUT120), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n960), .B1(new_n962), .B2(new_n964), .ZN(G60));
  AND2_X1   g779(.A1(new_n640), .A2(new_n641), .ZN(new_n966));
  NAND2_X1  g780(.A1(G478), .A2(G902), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT121), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT59), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n966), .B1(new_n892), .B2(new_n969), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n948), .A2(new_n966), .A3(new_n889), .A4(new_n969), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n955), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n970), .A2(new_n972), .ZN(G63));
  INV_X1    g787(.A(KEYINPUT123), .ZN(new_n974));
  NAND2_X1  g788(.A1(G217), .A2(G902), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT122), .Z(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT60), .Z(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n978), .B1(new_n883), .B2(new_n888), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n974), .B(new_n955), .C1(new_n979), .C2(new_n609), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT61), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n955), .B1(new_n979), .B2(new_n609), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n936), .A2(new_n678), .A3(new_n977), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n980), .B(new_n981), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  NOR3_X1   g798(.A1(new_n858), .A2(new_n847), .A3(new_n882), .ZN(new_n985));
  AOI21_X1  g799(.A(KEYINPUT53), .B1(new_n884), .B2(new_n887), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n977), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n945), .B1(new_n987), .B2(new_n608), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n979), .A2(new_n678), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n988), .B(new_n989), .C1(new_n974), .C2(KEYINPUT61), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n984), .A2(new_n990), .ZN(G66));
  INV_X1    g805(.A(G224), .ZN(new_n992));
  OAI21_X1  g806(.A(G953), .B1(new_n373), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n878), .A2(new_n881), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n993), .B1(new_n995), .B2(G953), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n938), .B1(G898), .B2(new_n192), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n996), .B(new_n997), .ZN(G69));
  AOI21_X1  g812(.A(new_n192), .B1(G227), .B2(G900), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n999), .A2(KEYINPUT124), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n779), .A2(new_n738), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n1001), .A2(new_n704), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(new_n730), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(KEYINPUT62), .ZN(new_n1004));
  INV_X1    g818(.A(new_n747), .ZN(new_n1005));
  NOR4_X1   g819(.A1(new_n1005), .A2(new_n726), .A3(new_n819), .A4(new_n871), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n835), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT62), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1002), .A2(new_n730), .A3(new_n1008), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n1004), .A2(new_n1007), .A3(new_n824), .A4(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n556), .B(new_n476), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n1011), .A2(G953), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1000), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n797), .A2(new_n704), .A3(new_n799), .A4(new_n1001), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n835), .A2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n810), .A2(new_n764), .A3(new_n784), .A4(new_n811), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1015), .A2(new_n824), .A3(new_n1016), .ZN(new_n1017));
  AND2_X1   g831(.A1(new_n1017), .A2(new_n192), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1011), .B1(G900), .B2(new_n192), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1013), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n999), .A2(KEYINPUT124), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1020), .B(new_n1021), .ZN(G72));
  NOR2_X1   g836(.A1(new_n711), .A2(new_n524), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1023), .ZN(new_n1024));
  NAND4_X1  g838(.A1(new_n1015), .A2(new_n824), .A3(new_n995), .A4(new_n1016), .ZN(new_n1025));
  XNOR2_X1  g839(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1026));
  NAND2_X1  g840(.A1(G472), .A2(G902), .ZN(new_n1027));
  XNOR2_X1  g841(.A(new_n1026), .B(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1024), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g843(.A(KEYINPUT126), .ZN(new_n1030));
  OR3_X1    g844(.A1(new_n1029), .A2(new_n1030), .A3(new_n945), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n1030), .B1(new_n1029), .B2(new_n945), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n1028), .B1(new_n1010), .B2(new_n994), .ZN(new_n1033));
  INV_X1    g847(.A(new_n1028), .ZN(new_n1034));
  INV_X1    g848(.A(KEYINPUT127), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n630), .B1(new_n1035), .B2(new_n551), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n711), .A2(KEYINPUT127), .A3(new_n525), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n1034), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  AOI22_X1  g852(.A1(new_n1033), .A2(new_n713), .B1(new_n936), .B2(new_n1038), .ZN(new_n1039));
  AND3_X1   g853(.A1(new_n1031), .A2(new_n1032), .A3(new_n1039), .ZN(G57));
endmodule


