

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736;

  XNOR2_X1 U373 ( .A(n416), .B(n379), .ZN(n432) );
  NOR2_X1 U374 ( .A1(n494), .A2(n491), .ZN(n493) );
  INV_X2 U375 ( .A(G953), .ZN(n724) );
  NOR2_X2 U376 ( .A1(n499), .A2(n498), .ZN(n500) );
  NOR2_X2 U377 ( .A1(n526), .A2(n536), .ZN(n527) );
  NAND2_X1 U378 ( .A1(n656), .A2(n655), .ZN(n653) );
  NOR2_X1 U379 ( .A1(n534), .A2(n563), .ZN(n531) );
  XNOR2_X1 U380 ( .A(n553), .B(n452), .ZN(n545) );
  NAND2_X1 U381 ( .A1(n520), .A2(n668), .ZN(n553) );
  XNOR2_X1 U382 ( .A(n406), .B(n405), .ZN(n703) );
  XNOR2_X2 U383 ( .A(n435), .B(n434), .ZN(n677) );
  NAND2_X1 U384 ( .A1(n367), .A2(n353), .ZN(n359) );
  AND2_X1 U385 ( .A1(n366), .A2(n368), .ZN(n367) );
  INV_X1 U386 ( .A(KEYINPUT70), .ZN(n358) );
  XNOR2_X1 U387 ( .A(n361), .B(KEYINPUT46), .ZN(n360) );
  NOR2_X1 U388 ( .A1(n734), .A2(n735), .ZN(n361) );
  INV_X1 U389 ( .A(KEYINPUT78), .ZN(n379) );
  XNOR2_X1 U390 ( .A(n370), .B(n369), .ZN(n511) );
  INV_X1 U391 ( .A(G478), .ZN(n369) );
  NAND2_X1 U392 ( .A1(n698), .A2(n481), .ZN(n370) );
  XNOR2_X1 U393 ( .A(n364), .B(n363), .ZN(n475) );
  XNOR2_X1 U394 ( .A(G134), .B(G122), .ZN(n363) );
  XNOR2_X1 U395 ( .A(n365), .B(KEYINPUT105), .ZN(n364) );
  XNOR2_X1 U396 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n365) );
  XNOR2_X1 U397 ( .A(KEYINPUT22), .B(KEYINPUT74), .ZN(n486) );
  AND2_X1 U398 ( .A1(n560), .A2(n639), .ZN(n368) );
  OR2_X1 U399 ( .A1(n506), .A2(KEYINPUT34), .ZN(n377) );
  OR2_X2 U400 ( .A1(n620), .A2(G902), .ZN(n362) );
  XNOR2_X1 U401 ( .A(n420), .B(n419), .ZN(n447) );
  XNOR2_X1 U402 ( .A(n720), .B(G146), .ZN(n427) );
  INV_X1 U403 ( .A(KEYINPUT48), .ZN(n355) );
  NAND2_X1 U404 ( .A1(n360), .A2(n357), .ZN(n356) );
  XNOR2_X1 U405 ( .A(n359), .B(n358), .ZN(n357) );
  XNOR2_X1 U406 ( .A(n473), .B(n472), .ZN(n512) );
  INV_X1 U407 ( .A(n511), .ZN(n513) );
  XNOR2_X1 U408 ( .A(n480), .B(n479), .ZN(n698) );
  AND2_X1 U409 ( .A1(n599), .A2(G953), .ZN(n707) );
  BUF_X1 U410 ( .A(n732), .Z(n733) );
  OR2_X1 U411 ( .A1(KEYINPUT86), .A2(n556), .ZN(n353) );
  XNOR2_X1 U412 ( .A(n429), .B(n428), .ZN(n538) );
  XNOR2_X1 U413 ( .A(n378), .B(n483), .ZN(n498) );
  XNOR2_X1 U414 ( .A(n444), .B(n386), .ZN(n720) );
  XNOR2_X1 U415 ( .A(n427), .B(n383), .ZN(n620) );
  OR2_X1 U416 ( .A1(n590), .A2(n589), .ZN(n354) );
  XNOR2_X2 U417 ( .A(n356), .B(n355), .ZN(n586) );
  XNOR2_X2 U418 ( .A(n362), .B(n392), .ZN(n541) );
  NOR2_X1 U419 ( .A1(n649), .A2(n561), .ZN(n366) );
  XNOR2_X2 U420 ( .A(n371), .B(G143), .ZN(n478) );
  XNOR2_X2 U421 ( .A(G128), .B(KEYINPUT64), .ZN(n371) );
  NAND2_X1 U422 ( .A1(n373), .A2(n372), .ZN(n378) );
  NAND2_X1 U423 ( .A1(n677), .A2(KEYINPUT34), .ZN(n372) );
  NOR2_X1 U424 ( .A1(n376), .A2(n374), .ZN(n373) );
  NAND2_X1 U425 ( .A1(n375), .A2(n482), .ZN(n374) );
  NAND2_X1 U426 ( .A1(n506), .A2(KEYINPUT34), .ZN(n375) );
  NOR2_X1 U427 ( .A1(n677), .A2(n377), .ZN(n376) );
  NAND2_X1 U428 ( .A1(n432), .A2(n661), .ZN(n665) );
  NAND2_X1 U429 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U430 ( .A(n519), .B(KEYINPUT45), .ZN(n582) );
  BUF_X1 U431 ( .A(n619), .Z(n702) );
  XNOR2_X2 U432 ( .A(n478), .B(KEYINPUT4), .ZN(n444) );
  INV_X1 U433 ( .A(n721), .ZN(n405) );
  XOR2_X1 U434 ( .A(G110), .B(G137), .Z(n380) );
  AND2_X1 U435 ( .A1(G210), .A2(n451), .ZN(n381) );
  XOR2_X1 U436 ( .A(KEYINPUT17), .B(KEYINPUT92), .Z(n382) );
  XOR2_X1 U437 ( .A(n443), .B(n390), .Z(n383) );
  INV_X1 U438 ( .A(KEYINPUT18), .ZN(n437) );
  XNOR2_X1 U439 ( .A(n438), .B(n437), .ZN(n439) );
  INV_X1 U440 ( .A(KEYINPUT0), .ZN(n460) );
  BUF_X1 U441 ( .A(n677), .Z(n686) );
  XNOR2_X1 U442 ( .A(n541), .B(n393), .ZN(n488) );
  BUF_X1 U443 ( .A(n611), .Z(n613) );
  BUF_X1 U444 ( .A(n520), .Z(n575) );
  XNOR2_X1 U445 ( .A(G137), .B(G134), .ZN(n385) );
  XNOR2_X1 U446 ( .A(G131), .B(KEYINPUT69), .ZN(n384) );
  XNOR2_X1 U447 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U448 ( .A(G104), .B(G110), .ZN(n387) );
  XNOR2_X1 U449 ( .A(n387), .B(G107), .ZN(n714) );
  XNOR2_X1 U450 ( .A(n714), .B(KEYINPUT73), .ZN(n443) );
  XNOR2_X1 U451 ( .A(G140), .B(G101), .ZN(n389) );
  NAND2_X1 U452 ( .A1(n724), .A2(G227), .ZN(n388) );
  XNOR2_X1 U453 ( .A(n389), .B(n388), .ZN(n390) );
  INV_X1 U454 ( .A(KEYINPUT71), .ZN(n391) );
  XNOR2_X1 U455 ( .A(n391), .B(G469), .ZN(n392) );
  XNOR2_X1 U456 ( .A(KEYINPUT65), .B(KEYINPUT1), .ZN(n393) );
  XNOR2_X1 U457 ( .A(G119), .B(G128), .ZN(n394) );
  XNOR2_X1 U458 ( .A(n380), .B(n394), .ZN(n398) );
  XOR2_X1 U459 ( .A(KEYINPUT23), .B(KEYINPUT72), .Z(n396) );
  XNOR2_X1 U460 ( .A(KEYINPUT24), .B(KEYINPUT96), .ZN(n395) );
  XNOR2_X1 U461 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U462 ( .A(n398), .B(n397), .Z(n402) );
  XOR2_X1 U463 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n400) );
  NAND2_X1 U464 ( .A1(G234), .A2(n724), .ZN(n399) );
  XNOR2_X1 U465 ( .A(n400), .B(n399), .ZN(n476) );
  NAND2_X1 U466 ( .A1(G221), .A2(n476), .ZN(n401) );
  XNOR2_X1 U467 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U468 ( .A(G146), .B(G125), .Z(n442) );
  XNOR2_X1 U469 ( .A(n442), .B(G140), .ZN(n404) );
  INV_X1 U470 ( .A(KEYINPUT10), .ZN(n403) );
  XNOR2_X1 U471 ( .A(n404), .B(n403), .ZN(n721) );
  NOR2_X2 U472 ( .A1(G902), .A2(n703), .ZN(n412) );
  XOR2_X1 U473 ( .A(KEYINPUT25), .B(KEYINPUT82), .Z(n409) );
  XNOR2_X1 U474 ( .A(G902), .B(KEYINPUT15), .ZN(n590) );
  NAND2_X1 U475 ( .A1(n590), .A2(G234), .ZN(n407) );
  XNOR2_X1 U476 ( .A(n407), .B(KEYINPUT20), .ZN(n413) );
  NAND2_X1 U477 ( .A1(n413), .A2(G217), .ZN(n408) );
  XNOR2_X1 U478 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U479 ( .A(KEYINPUT97), .B(n410), .ZN(n411) );
  XNOR2_X2 U480 ( .A(n412), .B(n411), .ZN(n656) );
  NAND2_X1 U481 ( .A1(G221), .A2(n413), .ZN(n415) );
  INV_X1 U482 ( .A(KEYINPUT21), .ZN(n414) );
  XNOR2_X1 U483 ( .A(n415), .B(n414), .ZN(n655) );
  OR2_X2 U484 ( .A1(n488), .A2(n653), .ZN(n416) );
  XNOR2_X1 U485 ( .A(G113), .B(G101), .ZN(n418) );
  INV_X1 U486 ( .A(G119), .ZN(n417) );
  XNOR2_X1 U487 ( .A(n418), .B(n417), .ZN(n420) );
  XOR2_X1 U488 ( .A(KEYINPUT3), .B(G116), .Z(n419) );
  XOR2_X1 U489 ( .A(KEYINPUT99), .B(KEYINPUT79), .Z(n422) );
  XNOR2_X1 U490 ( .A(KEYINPUT100), .B(KEYINPUT5), .ZN(n421) );
  XNOR2_X1 U491 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U492 ( .A(n447), .B(n423), .Z(n425) );
  NOR2_X1 U493 ( .A1(G953), .A2(G237), .ZN(n468) );
  NAND2_X1 U494 ( .A1(n468), .A2(G210), .ZN(n424) );
  XNOR2_X1 U495 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U496 ( .A(n427), .B(n426), .ZN(n596) );
  INV_X1 U497 ( .A(G902), .ZN(n481) );
  NAND2_X1 U498 ( .A1(n596), .A2(n481), .ZN(n429) );
  XNOR2_X1 U499 ( .A(G472), .B(KEYINPUT101), .ZN(n428) );
  INV_X1 U500 ( .A(KEYINPUT6), .ZN(n430) );
  XNOR2_X1 U501 ( .A(n538), .B(n430), .ZN(n549) );
  INV_X1 U502 ( .A(n549), .ZN(n431) );
  NAND2_X1 U503 ( .A1(n432), .A2(n431), .ZN(n435) );
  INV_X1 U504 ( .A(KEYINPUT106), .ZN(n433) );
  XNOR2_X1 U505 ( .A(n433), .B(KEYINPUT33), .ZN(n434) );
  XNOR2_X1 U506 ( .A(KEYINPUT90), .B(KEYINPUT83), .ZN(n436) );
  XNOR2_X1 U507 ( .A(n382), .B(n436), .ZN(n440) );
  NAND2_X1 U508 ( .A1(G224), .A2(n724), .ZN(n438) );
  XNOR2_X1 U509 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U510 ( .A(n442), .B(n441), .Z(n446) );
  XNOR2_X1 U511 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U512 ( .A(n446), .B(n445), .ZN(n449) );
  XNOR2_X1 U513 ( .A(n447), .B(KEYINPUT16), .ZN(n448) );
  XNOR2_X1 U514 ( .A(n448), .B(G122), .ZN(n713) );
  XNOR2_X1 U515 ( .A(n449), .B(n713), .ZN(n611) );
  INV_X1 U516 ( .A(n590), .ZN(n581) );
  OR2_X2 U517 ( .A1(n611), .A2(n581), .ZN(n450) );
  OR2_X1 U518 ( .A1(G237), .A2(G902), .ZN(n451) );
  XNOR2_X2 U519 ( .A(n450), .B(n381), .ZN(n520) );
  NAND2_X1 U520 ( .A1(G214), .A2(n451), .ZN(n668) );
  XNOR2_X1 U521 ( .A(KEYINPUT81), .B(KEYINPUT19), .ZN(n452) );
  NAND2_X1 U522 ( .A1(G234), .A2(G237), .ZN(n453) );
  XNOR2_X1 U523 ( .A(n453), .B(KEYINPUT14), .ZN(n454) );
  NAND2_X1 U524 ( .A1(G952), .A2(n454), .ZN(n685) );
  NOR2_X1 U525 ( .A1(G953), .A2(n685), .ZN(n525) );
  NAND2_X1 U526 ( .A1(n454), .A2(G902), .ZN(n455) );
  XNOR2_X1 U527 ( .A(n455), .B(KEYINPUT94), .ZN(n522) );
  NOR2_X1 U528 ( .A1(G898), .A2(n724), .ZN(n456) );
  XNOR2_X1 U529 ( .A(KEYINPUT93), .B(n456), .ZN(n716) );
  NOR2_X1 U530 ( .A1(n522), .A2(n716), .ZN(n457) );
  XOR2_X1 U531 ( .A(KEYINPUT95), .B(n457), .Z(n458) );
  NOR2_X1 U532 ( .A1(n525), .A2(n458), .ZN(n459) );
  NOR2_X2 U533 ( .A1(n545), .A2(n459), .ZN(n461) );
  XNOR2_X2 U534 ( .A(n461), .B(n460), .ZN(n506) );
  XOR2_X1 U535 ( .A(G122), .B(G104), .Z(n463) );
  XNOR2_X1 U536 ( .A(G113), .B(G143), .ZN(n462) );
  XNOR2_X1 U537 ( .A(n463), .B(n462), .ZN(n467) );
  XOR2_X1 U538 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n465) );
  XNOR2_X1 U539 ( .A(G131), .B(KEYINPUT104), .ZN(n464) );
  XNOR2_X1 U540 ( .A(n465), .B(n464), .ZN(n466) );
  XOR2_X1 U541 ( .A(n467), .B(n466), .Z(n470) );
  AND2_X1 U542 ( .A1(G214), .A2(n468), .ZN(n469) );
  XNOR2_X1 U543 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U544 ( .A(n471), .B(n721), .ZN(n604) );
  NAND2_X1 U545 ( .A1(n604), .A2(n481), .ZN(n473) );
  XOR2_X1 U546 ( .A(KEYINPUT13), .B(G475), .Z(n472) );
  XNOR2_X1 U547 ( .A(G116), .B(G107), .ZN(n474) );
  XNOR2_X1 U548 ( .A(n475), .B(n474), .ZN(n480) );
  NAND2_X1 U549 ( .A1(G217), .A2(n476), .ZN(n477) );
  XNOR2_X1 U550 ( .A(n478), .B(n477), .ZN(n479) );
  NAND2_X1 U551 ( .A1(n512), .A2(n513), .ZN(n562) );
  INV_X1 U552 ( .A(n562), .ZN(n482) );
  XNOR2_X1 U553 ( .A(KEYINPUT84), .B(KEYINPUT35), .ZN(n483) );
  XOR2_X1 U554 ( .A(n498), .B(G122), .Z(G24) );
  INV_X1 U555 ( .A(n506), .ZN(n485) );
  NOR2_X1 U556 ( .A1(n512), .A2(n513), .ZN(n533) );
  AND2_X1 U557 ( .A1(n655), .A2(n533), .ZN(n484) );
  NAND2_X1 U558 ( .A1(n485), .A2(n484), .ZN(n487) );
  XNOR2_X1 U559 ( .A(n487), .B(n486), .ZN(n494) );
  BUF_X1 U560 ( .A(n488), .Z(n489) );
  NOR2_X1 U561 ( .A1(n489), .A2(n656), .ZN(n490) );
  NAND2_X1 U562 ( .A1(n490), .A2(n549), .ZN(n491) );
  INV_X1 U563 ( .A(KEYINPUT32), .ZN(n492) );
  XNOR2_X1 U564 ( .A(n493), .B(n492), .ZN(n732) );
  INV_X1 U565 ( .A(n494), .ZN(n503) );
  INV_X1 U566 ( .A(n656), .ZN(n495) );
  AND2_X1 U567 ( .A1(n538), .A2(n495), .ZN(n496) );
  AND2_X1 U568 ( .A1(n489), .A2(n496), .ZN(n497) );
  NAND2_X1 U569 ( .A1(n503), .A2(n497), .ZN(n633) );
  NAND2_X1 U570 ( .A1(n732), .A2(n633), .ZN(n499) );
  XNOR2_X1 U571 ( .A(n500), .B(KEYINPUT44), .ZN(n518) );
  AND2_X1 U572 ( .A1(n489), .A2(n656), .ZN(n501) );
  AND2_X1 U573 ( .A1(n501), .A2(n549), .ZN(n502) );
  NAND2_X1 U574 ( .A1(n503), .A2(n502), .ZN(n626) );
  NOR2_X1 U575 ( .A1(n506), .A2(n665), .ZN(n504) );
  XOR2_X1 U576 ( .A(KEYINPUT103), .B(n504), .Z(n505) );
  XNOR2_X1 U577 ( .A(KEYINPUT31), .B(n505), .ZN(n646) );
  INV_X1 U578 ( .A(n538), .ZN(n661) );
  INV_X1 U579 ( .A(n653), .ZN(n507) );
  NAND2_X1 U580 ( .A1(n507), .A2(n541), .ZN(n508) );
  XNOR2_X1 U581 ( .A(n508), .B(KEYINPUT98), .ZN(n526) );
  NOR2_X1 U582 ( .A1(n661), .A2(n526), .ZN(n509) );
  NAND2_X1 U583 ( .A1(n485), .A2(n509), .ZN(n510) );
  XNOR2_X1 U584 ( .A(KEYINPUT102), .B(n510), .ZN(n630) );
  NAND2_X1 U585 ( .A1(n646), .A2(n630), .ZN(n515) );
  NAND2_X1 U586 ( .A1(n512), .A2(n511), .ZN(n551) );
  INV_X1 U587 ( .A(n512), .ZN(n514) );
  NAND2_X1 U588 ( .A1(n514), .A2(n513), .ZN(n647) );
  NAND2_X1 U589 ( .A1(n551), .A2(n647), .ZN(n557) );
  NAND2_X1 U590 ( .A1(n515), .A2(n557), .ZN(n516) );
  AND2_X1 U591 ( .A1(n626), .A2(n516), .ZN(n517) );
  NAND2_X1 U592 ( .A1(n518), .A2(n517), .ZN(n519) );
  BUF_X1 U593 ( .A(n582), .Z(n708) );
  XNOR2_X1 U594 ( .A(KEYINPUT77), .B(KEYINPUT38), .ZN(n521) );
  XOR2_X1 U595 ( .A(n575), .B(n521), .Z(n534) );
  OR2_X1 U596 ( .A1(n522), .A2(n724), .ZN(n523) );
  NOR2_X1 U597 ( .A1(G900), .A2(n523), .ZN(n524) );
  NOR2_X1 U598 ( .A1(n525), .A2(n524), .ZN(n536) );
  XNOR2_X1 U599 ( .A(n527), .B(KEYINPUT80), .ZN(n530) );
  NAND2_X1 U600 ( .A1(n661), .A2(n668), .ZN(n528) );
  XOR2_X1 U601 ( .A(KEYINPUT30), .B(n528), .Z(n529) );
  NAND2_X1 U602 ( .A1(n530), .A2(n529), .ZN(n563) );
  XNOR2_X1 U603 ( .A(n531), .B(KEYINPUT39), .ZN(n565) );
  NOR2_X1 U604 ( .A1(n565), .A2(n551), .ZN(n532) );
  XNOR2_X1 U605 ( .A(n532), .B(KEYINPUT40), .ZN(n734) );
  INV_X1 U606 ( .A(n533), .ZN(n671) );
  INV_X1 U607 ( .A(n534), .ZN(n669) );
  NAND2_X1 U608 ( .A1(n669), .A2(n668), .ZN(n674) );
  NOR2_X1 U609 ( .A1(n671), .A2(n674), .ZN(n535) );
  XNOR2_X1 U610 ( .A(n535), .B(KEYINPUT41), .ZN(n687) );
  XNOR2_X1 U611 ( .A(KEYINPUT109), .B(KEYINPUT28), .ZN(n540) );
  NOR2_X1 U612 ( .A1(n656), .A2(n536), .ZN(n537) );
  NAND2_X1 U613 ( .A1(n537), .A2(n655), .ZN(n550) );
  NOR2_X1 U614 ( .A1(n550), .A2(n538), .ZN(n539) );
  XOR2_X1 U615 ( .A(n540), .B(n539), .Z(n542) );
  NAND2_X1 U616 ( .A1(n542), .A2(n541), .ZN(n546) );
  NOR2_X1 U617 ( .A1(n687), .A2(n546), .ZN(n543) );
  XNOR2_X1 U618 ( .A(n543), .B(KEYINPUT42), .ZN(n735) );
  INV_X1 U619 ( .A(n557), .ZN(n673) );
  NOR2_X1 U620 ( .A1(n673), .A2(KEYINPUT47), .ZN(n544) );
  XNOR2_X1 U621 ( .A(KEYINPUT76), .B(n544), .ZN(n547) );
  NOR2_X1 U622 ( .A1(n546), .A2(n545), .ZN(n641) );
  NAND2_X1 U623 ( .A1(n547), .A2(n641), .ZN(n548) );
  XNOR2_X1 U624 ( .A(n548), .B(KEYINPUT75), .ZN(n561) );
  NOR2_X1 U625 ( .A1(n550), .A2(n549), .ZN(n552) );
  XOR2_X1 U626 ( .A(KEYINPUT107), .B(n551), .Z(n643) );
  INV_X1 U627 ( .A(n643), .ZN(n640) );
  NAND2_X1 U628 ( .A1(n552), .A2(n640), .ZN(n569) );
  NOR2_X1 U629 ( .A1(n569), .A2(n553), .ZN(n554) );
  XOR2_X1 U630 ( .A(KEYINPUT36), .B(n554), .Z(n555) );
  NOR2_X1 U631 ( .A1(n555), .A2(n489), .ZN(n649) );
  INV_X1 U632 ( .A(n641), .ZN(n634) );
  AND2_X1 U633 ( .A1(n634), .A2(KEYINPUT47), .ZN(n556) );
  NAND2_X1 U634 ( .A1(n634), .A2(KEYINPUT86), .ZN(n558) );
  NAND2_X1 U635 ( .A1(n558), .A2(n557), .ZN(n559) );
  NAND2_X1 U636 ( .A1(n559), .A2(KEYINPUT47), .ZN(n560) );
  NOR2_X1 U637 ( .A1(n563), .A2(n562), .ZN(n564) );
  NAND2_X1 U638 ( .A1(n575), .A2(n564), .ZN(n639) );
  INV_X1 U639 ( .A(n586), .ZN(n579) );
  INV_X1 U640 ( .A(n565), .ZN(n567) );
  INV_X1 U641 ( .A(n647), .ZN(n566) );
  NAND2_X1 U642 ( .A1(n567), .A2(n566), .ZN(n652) );
  NAND2_X1 U643 ( .A1(n652), .A2(KEYINPUT2), .ZN(n568) );
  XNOR2_X1 U644 ( .A(n568), .B(KEYINPUT85), .ZN(n577) );
  INV_X1 U645 ( .A(n569), .ZN(n570) );
  NAND2_X1 U646 ( .A1(n570), .A2(n668), .ZN(n572) );
  INV_X1 U647 ( .A(n489), .ZN(n571) );
  NOR2_X1 U648 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U649 ( .A(n573), .B(KEYINPUT43), .ZN(n574) );
  NOR2_X1 U650 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U651 ( .A(KEYINPUT108), .B(n576), .ZN(n731) );
  INV_X1 U652 ( .A(n731), .ZN(n584) );
  NAND2_X1 U653 ( .A1(n577), .A2(n584), .ZN(n578) );
  NOR2_X1 U654 ( .A1(n579), .A2(n578), .ZN(n580) );
  AND2_X1 U655 ( .A1(n708), .A2(n580), .ZN(n694) );
  INV_X1 U656 ( .A(n694), .ZN(n593) );
  XNOR2_X1 U657 ( .A(n583), .B(KEYINPUT87), .ZN(n588) );
  AND2_X1 U658 ( .A1(n652), .A2(n584), .ZN(n585) );
  NAND2_X1 U659 ( .A1(n586), .A2(n585), .ZN(n719) );
  INV_X1 U660 ( .A(n719), .ZN(n587) );
  NAND2_X1 U661 ( .A1(n588), .A2(n587), .ZN(n591) );
  INV_X1 U662 ( .A(KEYINPUT2), .ZN(n589) );
  NAND2_X1 U663 ( .A1(n591), .A2(n354), .ZN(n592) );
  AND2_X2 U664 ( .A1(n593), .A2(n592), .ZN(n619) );
  NAND2_X1 U665 ( .A1(n619), .A2(G472), .ZN(n598) );
  XNOR2_X1 U666 ( .A(KEYINPUT91), .B(KEYINPUT110), .ZN(n594) );
  XNOR2_X1 U667 ( .A(n594), .B(KEYINPUT62), .ZN(n595) );
  XNOR2_X1 U668 ( .A(n596), .B(n595), .ZN(n597) );
  XNOR2_X1 U669 ( .A(n598), .B(n597), .ZN(n600) );
  INV_X1 U670 ( .A(G952), .ZN(n599) );
  NOR2_X2 U671 ( .A1(n600), .A2(n707), .ZN(n602) );
  XNOR2_X1 U672 ( .A(KEYINPUT89), .B(KEYINPUT63), .ZN(n601) );
  XNOR2_X1 U673 ( .A(n602), .B(n601), .ZN(G57) );
  NAND2_X1 U674 ( .A1(n619), .A2(G475), .ZN(n606) );
  XNOR2_X1 U675 ( .A(KEYINPUT66), .B(KEYINPUT59), .ZN(n603) );
  XNOR2_X1 U676 ( .A(n604), .B(n603), .ZN(n605) );
  XNOR2_X1 U677 ( .A(n606), .B(n605), .ZN(n607) );
  NOR2_X2 U678 ( .A1(n607), .A2(n707), .ZN(n610) );
  XNOR2_X1 U679 ( .A(KEYINPUT122), .B(KEYINPUT60), .ZN(n608) );
  XOR2_X1 U680 ( .A(n608), .B(KEYINPUT67), .Z(n609) );
  XNOR2_X1 U681 ( .A(n610), .B(n609), .ZN(G60) );
  NAND2_X1 U682 ( .A1(n619), .A2(G210), .ZN(n615) );
  XOR2_X1 U683 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n612) );
  XNOR2_X1 U684 ( .A(n613), .B(n612), .ZN(n614) );
  XNOR2_X1 U685 ( .A(n615), .B(n614), .ZN(n616) );
  NOR2_X2 U686 ( .A1(n616), .A2(n707), .ZN(n618) );
  XNOR2_X1 U687 ( .A(KEYINPUT88), .B(KEYINPUT56), .ZN(n617) );
  XNOR2_X1 U688 ( .A(n618), .B(n617), .ZN(G51) );
  NAND2_X1 U689 ( .A1(n702), .A2(G469), .ZN(n623) );
  XOR2_X1 U690 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n621) );
  XNOR2_X1 U691 ( .A(n620), .B(n621), .ZN(n622) );
  XNOR2_X1 U692 ( .A(n623), .B(n622), .ZN(n624) );
  NOR2_X1 U693 ( .A1(n624), .A2(n707), .ZN(G54) );
  XOR2_X1 U694 ( .A(G101), .B(KEYINPUT111), .Z(n625) );
  XNOR2_X1 U695 ( .A(n626), .B(n625), .ZN(G3) );
  NOR2_X1 U696 ( .A1(n630), .A2(n643), .ZN(n627) );
  XOR2_X1 U697 ( .A(G104), .B(n627), .Z(G6) );
  XOR2_X1 U698 ( .A(KEYINPUT26), .B(KEYINPUT112), .Z(n629) );
  XNOR2_X1 U699 ( .A(G107), .B(KEYINPUT27), .ZN(n628) );
  XNOR2_X1 U700 ( .A(n629), .B(n628), .ZN(n632) );
  NOR2_X1 U701 ( .A1(n630), .A2(n647), .ZN(n631) );
  XOR2_X1 U702 ( .A(n632), .B(n631), .Z(G9) );
  XNOR2_X1 U703 ( .A(G110), .B(n633), .ZN(G12) );
  NOR2_X1 U704 ( .A1(n647), .A2(n634), .ZN(n638) );
  XOR2_X1 U705 ( .A(KEYINPUT113), .B(KEYINPUT29), .Z(n636) );
  XNOR2_X1 U706 ( .A(G128), .B(KEYINPUT114), .ZN(n635) );
  XNOR2_X1 U707 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U708 ( .A(n638), .B(n637), .ZN(G30) );
  XNOR2_X1 U709 ( .A(G143), .B(n639), .ZN(G45) );
  NAND2_X1 U710 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U711 ( .A(n642), .B(G146), .ZN(G48) );
  NOR2_X1 U712 ( .A1(n643), .A2(n646), .ZN(n645) );
  XNOR2_X1 U713 ( .A(G113), .B(KEYINPUT115), .ZN(n644) );
  XNOR2_X1 U714 ( .A(n645), .B(n644), .ZN(G15) );
  NOR2_X1 U715 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U716 ( .A(G116), .B(n648), .Z(G18) );
  XNOR2_X1 U717 ( .A(n649), .B(KEYINPUT37), .ZN(n650) );
  XNOR2_X1 U718 ( .A(n650), .B(KEYINPUT116), .ZN(n651) );
  XNOR2_X1 U719 ( .A(G125), .B(n651), .ZN(G27) );
  XNOR2_X1 U720 ( .A(G134), .B(n652), .ZN(G36) );
  NAND2_X1 U721 ( .A1(n489), .A2(n653), .ZN(n654) );
  XNOR2_X1 U722 ( .A(n654), .B(KEYINPUT50), .ZN(n663) );
  NOR2_X1 U723 ( .A1(n656), .A2(n655), .ZN(n658) );
  XNOR2_X1 U724 ( .A(KEYINPUT118), .B(KEYINPUT49), .ZN(n657) );
  XNOR2_X1 U725 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U726 ( .A(KEYINPUT117), .B(n659), .ZN(n660) );
  NOR2_X1 U727 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U728 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U729 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U730 ( .A(KEYINPUT51), .B(n666), .ZN(n667) );
  NOR2_X1 U731 ( .A1(n687), .A2(n667), .ZN(n681) );
  NOR2_X1 U732 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U733 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U734 ( .A(KEYINPUT119), .B(n672), .Z(n676) );
  NOR2_X1 U735 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U736 ( .A1(n676), .A2(n675), .ZN(n678) );
  NOR2_X1 U737 ( .A1(n678), .A2(n686), .ZN(n679) );
  XNOR2_X1 U738 ( .A(n679), .B(KEYINPUT120), .ZN(n680) );
  NOR2_X1 U739 ( .A1(n681), .A2(n680), .ZN(n683) );
  XOR2_X1 U740 ( .A(KEYINPUT52), .B(KEYINPUT121), .Z(n682) );
  XNOR2_X1 U741 ( .A(n683), .B(n682), .ZN(n684) );
  NOR2_X1 U742 ( .A1(n685), .A2(n684), .ZN(n689) );
  NOR2_X1 U743 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U744 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U745 ( .A1(n690), .A2(n724), .ZN(n696) );
  INV_X1 U746 ( .A(n708), .ZN(n691) );
  NOR2_X1 U747 ( .A1(n691), .A2(n719), .ZN(n692) );
  NOR2_X1 U748 ( .A1(n692), .A2(KEYINPUT2), .ZN(n693) );
  NOR2_X1 U749 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U750 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U751 ( .A(n697), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U752 ( .A1(n702), .A2(G478), .ZN(n700) );
  XNOR2_X1 U753 ( .A(n698), .B(KEYINPUT123), .ZN(n699) );
  XNOR2_X1 U754 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U755 ( .A1(n707), .A2(n701), .ZN(G63) );
  NAND2_X1 U756 ( .A1(n702), .A2(G217), .ZN(n705) );
  XNOR2_X1 U757 ( .A(n703), .B(KEYINPUT124), .ZN(n704) );
  XNOR2_X1 U758 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U759 ( .A1(n707), .A2(n706), .ZN(G66) );
  NAND2_X1 U760 ( .A1(n708), .A2(n724), .ZN(n712) );
  NAND2_X1 U761 ( .A1(G953), .A2(G224), .ZN(n709) );
  XNOR2_X1 U762 ( .A(KEYINPUT61), .B(n709), .ZN(n710) );
  NAND2_X1 U763 ( .A1(n710), .A2(G898), .ZN(n711) );
  NAND2_X1 U764 ( .A1(n712), .A2(n711), .ZN(n718) );
  XOR2_X1 U765 ( .A(n714), .B(n713), .Z(n715) );
  NAND2_X1 U766 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U767 ( .A(n718), .B(n717), .Z(G69) );
  XOR2_X1 U768 ( .A(KEYINPUT126), .B(n719), .Z(n723) );
  XNOR2_X1 U769 ( .A(n721), .B(KEYINPUT125), .ZN(n722) );
  XOR2_X1 U770 ( .A(n720), .B(n722), .Z(n726) );
  XOR2_X1 U771 ( .A(n723), .B(n726), .Z(n725) );
  NAND2_X1 U772 ( .A1(n725), .A2(n724), .ZN(n730) );
  XNOR2_X1 U773 ( .A(G227), .B(n726), .ZN(n727) );
  NAND2_X1 U774 ( .A1(n727), .A2(G900), .ZN(n728) );
  NAND2_X1 U775 ( .A1(n728), .A2(G953), .ZN(n729) );
  NAND2_X1 U776 ( .A1(n730), .A2(n729), .ZN(G72) );
  XOR2_X1 U777 ( .A(G140), .B(n731), .Z(G42) );
  XNOR2_X1 U778 ( .A(n733), .B(G119), .ZN(G21) );
  XOR2_X1 U779 ( .A(G131), .B(n734), .Z(G33) );
  XNOR2_X1 U780 ( .A(G137), .B(KEYINPUT127), .ZN(n736) );
  XNOR2_X1 U781 ( .A(n736), .B(n735), .ZN(G39) );
endmodule

