

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771;

  OR2_X1 U369 ( .A1(n741), .A2(G902), .ZN(n393) );
  INV_X2 U370 ( .A(G953), .ZN(n761) );
  AND2_X1 U371 ( .A1(n426), .A2(n422), .ZN(n421) );
  XOR2_X1 U372 ( .A(G140), .B(KEYINPUT10), .Z(n348) );
  NOR2_X1 U373 ( .A1(n698), .A2(n609), .ZN(n610) );
  XNOR2_X2 U374 ( .A(n496), .B(n495), .ZN(n560) );
  NOR2_X2 U375 ( .A1(G902), .A2(n730), .ZN(n496) );
  XNOR2_X1 U376 ( .A(n606), .B(KEYINPUT109), .ZN(n699) );
  INV_X1 U377 ( .A(n667), .ZN(n663) );
  INV_X1 U378 ( .A(n680), .ZN(n349) );
  NOR2_X2 U379 ( .A1(n771), .A2(n770), .ZN(n611) );
  NOR2_X1 U380 ( .A1(n618), .A2(n540), .ZN(n673) );
  INV_X1 U381 ( .A(n677), .ZN(n392) );
  BUF_X1 U382 ( .A(n676), .Z(n677) );
  XNOR2_X1 U383 ( .A(n440), .B(G472), .ZN(n687) );
  XNOR2_X1 U384 ( .A(n759), .B(n512), .ZN(n725) );
  BUF_X1 U385 ( .A(G104), .Z(n362) );
  NAND2_X1 U386 ( .A1(n679), .A2(n625), .ZN(n626) );
  INV_X1 U387 ( .A(n680), .ZN(n350) );
  AND2_X1 U388 ( .A1(n369), .A2(n613), .ZN(n368) );
  NAND2_X1 U389 ( .A1(n385), .A2(n380), .ZN(n578) );
  XNOR2_X1 U390 ( .A(n605), .B(KEYINPUT40), .ZN(n771) );
  AND2_X1 U391 ( .A1(n663), .A2(n620), .ZN(n605) );
  XNOR2_X1 U392 ( .A(n601), .B(KEYINPUT38), .ZN(n702) );
  NAND2_X1 U393 ( .A1(n402), .A2(n399), .ZN(n522) );
  AND2_X1 U394 ( .A1(n560), .A2(n534), .ZN(n704) );
  XNOR2_X1 U395 ( .A(n507), .B(n506), .ZN(n534) );
  XNOR2_X1 U396 ( .A(n725), .B(n724), .ZN(n726) );
  XNOR2_X1 U397 ( .A(n732), .B(n731), .ZN(n733) );
  BUF_X1 U398 ( .A(n511), .Z(n356) );
  XNOR2_X1 U399 ( .A(n511), .B(n467), .ZN(n414) );
  XNOR2_X1 U400 ( .A(n412), .B(n411), .ZN(n468) );
  NAND2_X1 U401 ( .A1(n351), .A2(n354), .ZN(n750) );
  NAND2_X1 U402 ( .A1(n352), .A2(n353), .ZN(n351) );
  NAND2_X1 U403 ( .A1(n420), .A2(n418), .ZN(n417) );
  XNOR2_X1 U404 ( .A(n528), .B(KEYINPUT19), .ZN(n590) );
  NAND2_X1 U405 ( .A1(n590), .A2(n533), .ZN(n410) );
  XNOR2_X1 U406 ( .A(n481), .B(n480), .ZN(n526) );
  NAND2_X1 U407 ( .A1(n414), .A2(n468), .ZN(n354) );
  INV_X1 U408 ( .A(n414), .ZN(n352) );
  INV_X1 U409 ( .A(n468), .ZN(n353) );
  BUF_X1 U410 ( .A(n627), .Z(n355) );
  NAND2_X1 U411 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X2 U412 ( .A(n375), .B(n519), .ZN(n567) );
  XNOR2_X2 U413 ( .A(n608), .B(n607), .ZN(n698) );
  AND2_X1 U414 ( .A1(n379), .A2(n572), .ZN(n389) );
  OR2_X1 U415 ( .A1(n725), .A2(n400), .ZN(n399) );
  AND2_X1 U416 ( .A1(n404), .A2(n403), .ZN(n402) );
  NAND2_X1 U417 ( .A1(G469), .A2(n401), .ZN(n400) );
  XNOR2_X1 U418 ( .A(KEYINPUT3), .B(G119), .ZN(n433) );
  XNOR2_X1 U419 ( .A(G131), .B(G143), .ZN(n482) );
  XOR2_X1 U420 ( .A(KEYINPUT102), .B(KEYINPUT11), .Z(n485) );
  NOR2_X1 U421 ( .A1(n555), .A2(KEYINPUT34), .ZN(n391) );
  NOR2_X1 U422 ( .A1(n384), .A2(n382), .ZN(n381) );
  INV_X1 U423 ( .A(n389), .ZN(n384) );
  XNOR2_X1 U424 ( .A(n522), .B(n374), .ZN(n690) );
  INV_X1 U425 ( .A(KEYINPUT1), .ZN(n374) );
  XNOR2_X1 U426 ( .A(KEYINPUT16), .B(G122), .ZN(n467) );
  XNOR2_X1 U427 ( .A(G128), .B(G137), .ZN(n446) );
  XNOR2_X1 U428 ( .A(G137), .B(G131), .ZN(n437) );
  INV_X1 U429 ( .A(n541), .ZN(n425) );
  XNOR2_X1 U430 ( .A(n461), .B(n395), .ZN(n394) );
  INV_X1 U431 ( .A(KEYINPUT99), .ZN(n395) );
  BUF_X1 U432 ( .A(n687), .Z(n375) );
  BUF_X1 U433 ( .A(n690), .Z(n367) );
  NOR2_X1 U434 ( .A1(n598), .A2(n597), .ZN(n613) );
  XNOR2_X1 U435 ( .A(n571), .B(n570), .ZN(n676) );
  NAND2_X1 U436 ( .A1(n513), .A2(G902), .ZN(n403) );
  XNOR2_X1 U437 ( .A(n583), .B(KEYINPUT64), .ZN(n584) );
  XNOR2_X1 U438 ( .A(KEYINPUT72), .B(G116), .ZN(n411) );
  XNOR2_X1 U439 ( .A(n433), .B(n413), .ZN(n412) );
  INV_X1 U440 ( .A(G113), .ZN(n413) );
  NOR2_X1 U441 ( .A1(G953), .A2(G237), .ZN(n488) );
  XNOR2_X1 U442 ( .A(G122), .B(KEYINPUT12), .ZN(n484) );
  INV_X1 U443 ( .A(KEYINPUT15), .ZN(n455) );
  XNOR2_X1 U444 ( .A(KEYINPUT4), .B(G146), .ZN(n473) );
  XNOR2_X1 U445 ( .A(n553), .B(KEYINPUT76), .ZN(n566) );
  NAND2_X1 U446 ( .A1(n690), .A2(n552), .ZN(n553) );
  BUF_X1 U447 ( .A(n526), .Z(n601) );
  XNOR2_X1 U448 ( .A(n460), .B(n459), .ZN(n461) );
  INV_X1 U449 ( .A(KEYINPUT25), .ZN(n459) );
  INV_X1 U450 ( .A(KEYINPUT0), .ZN(n409) );
  XNOR2_X1 U451 ( .A(G116), .B(G107), .ZN(n500) );
  AND2_X1 U452 ( .A1(n373), .A2(n387), .ZN(n385) );
  XNOR2_X1 U453 ( .A(n494), .B(G475), .ZN(n495) );
  NAND2_X1 U454 ( .A1(n350), .A2(G472), .ZN(n408) );
  XOR2_X1 U455 ( .A(KEYINPUT62), .B(n647), .Z(n648) );
  XNOR2_X1 U456 ( .A(n454), .B(n491), .ZN(n741) );
  NAND2_X1 U457 ( .A1(n350), .A2(G475), .ZN(n407) );
  XNOR2_X1 U458 ( .A(KEYINPUT78), .B(G140), .ZN(n509) );
  NAND2_X1 U459 ( .A1(n349), .A2(G469), .ZN(n406) );
  NAND2_X1 U460 ( .A1(n349), .A2(G210), .ZN(n405) );
  XNOR2_X1 U461 ( .A(n640), .B(n639), .ZN(n641) );
  AND2_X1 U462 ( .A1(n643), .A2(G953), .ZN(n744) );
  NAND2_X1 U463 ( .A1(n423), .A2(n360), .ZN(n422) );
  NAND2_X1 U464 ( .A1(n425), .A2(n424), .ZN(n423) );
  NOR2_X1 U465 ( .A1(n541), .A2(n419), .ZN(n418) );
  OR2_X1 U466 ( .A1(n567), .A2(n360), .ZN(n419) );
  NOR2_X1 U467 ( .A1(n609), .A2(n592), .ZN(n664) );
  INV_X1 U468 ( .A(KEYINPUT85), .ZN(n377) );
  AND2_X1 U469 ( .A1(n371), .A2(n370), .ZN(n722) );
  INV_X1 U470 ( .A(G953), .ZN(n370) );
  XNOR2_X1 U471 ( .A(n721), .B(KEYINPUT119), .ZN(n371) );
  XOR2_X1 U472 ( .A(n446), .B(KEYINPUT97), .Z(n357) );
  XOR2_X1 U473 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n358) );
  AND2_X1 U474 ( .A1(n391), .A2(n573), .ZN(n359) );
  INV_X1 U475 ( .A(G902), .ZN(n401) );
  XOR2_X1 U476 ( .A(n542), .B(KEYINPUT68), .Z(n360) );
  BUF_X1 U477 ( .A(n551), .Z(n361) );
  NOR2_X1 U478 ( .A1(n564), .A2(n565), .ZN(n366) );
  XNOR2_X1 U479 ( .A(n361), .B(KEYINPUT106), .ZN(n363) );
  XNOR2_X1 U480 ( .A(n551), .B(KEYINPUT106), .ZN(n769) );
  NAND2_X1 U481 ( .A1(n421), .A2(n417), .ZN(n364) );
  NAND2_X1 U482 ( .A1(n421), .A2(n417), .ZN(n547) );
  NOR2_X1 U483 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U484 ( .A1(n636), .A2(n680), .ZN(n740) );
  XOR2_X1 U485 ( .A(n362), .B(G113), .Z(n483) );
  NAND2_X1 U486 ( .A1(n366), .A2(n365), .ZN(n397) );
  XNOR2_X1 U487 ( .A(n372), .B(n574), .ZN(n365) );
  XNOR2_X1 U488 ( .A(n750), .B(n476), .ZN(n637) );
  AND2_X2 U489 ( .A1(n612), .A2(n368), .ZN(n619) );
  INV_X1 U490 ( .A(n673), .ZN(n369) );
  NAND2_X1 U491 ( .A1(n578), .A2(KEYINPUT44), .ZN(n372) );
  NAND2_X1 U492 ( .A1(n386), .A2(n573), .ZN(n373) );
  INV_X1 U493 ( .A(n367), .ZN(n540) );
  OR2_X2 U494 ( .A1(n623), .A2(KEYINPUT2), .ZN(n679) );
  NAND2_X1 U495 ( .A1(n637), .A2(n624), .ZN(n481) );
  NAND2_X1 U496 ( .A1(n527), .A2(n701), .ZN(n528) );
  XNOR2_X1 U497 ( .A(n376), .B(n584), .ZN(n627) );
  NAND2_X1 U498 ( .A1(n396), .A2(n582), .ZN(n376) );
  XNOR2_X1 U499 ( .A(n378), .B(n377), .ZN(n550) );
  NOR2_X2 U500 ( .A1(n546), .A2(n567), .ZN(n378) );
  NAND2_X1 U501 ( .A1(n676), .A2(KEYINPUT34), .ZN(n388) );
  NAND2_X1 U502 ( .A1(n392), .A2(n391), .ZN(n390) );
  NAND2_X1 U503 ( .A1(n392), .A2(n359), .ZN(n387) );
  NAND2_X1 U504 ( .A1(n388), .A2(n389), .ZN(n386) );
  NAND2_X1 U505 ( .A1(n555), .A2(KEYINPUT34), .ZN(n379) );
  NAND2_X1 U506 ( .A1(n381), .A2(n390), .ZN(n380) );
  NAND2_X1 U507 ( .A1(n388), .A2(n383), .ZN(n382) );
  INV_X1 U508 ( .A(n573), .ZN(n383) );
  XNOR2_X2 U509 ( .A(n394), .B(n393), .ZN(n543) );
  XNOR2_X1 U510 ( .A(n397), .B(n575), .ZN(n396) );
  XNOR2_X2 U511 ( .A(n398), .B(G143), .ZN(n469) );
  XNOR2_X2 U512 ( .A(G128), .B(KEYINPUT65), .ZN(n398) );
  NAND2_X1 U513 ( .A1(n725), .A2(n513), .ZN(n404) );
  OR2_X1 U514 ( .A1(n636), .A2(n405), .ZN(n642) );
  OR2_X1 U515 ( .A1(n636), .A2(n406), .ZN(n727) );
  OR2_X1 U516 ( .A1(n636), .A2(n407), .ZN(n734) );
  OR2_X1 U517 ( .A1(n636), .A2(n408), .ZN(n649) );
  NAND2_X1 U518 ( .A1(n740), .A2(G478), .ZN(n737) );
  XNOR2_X2 U519 ( .A(n469), .B(G134), .ZN(n504) );
  INV_X1 U520 ( .A(n536), .ZN(n555) );
  XNOR2_X2 U521 ( .A(n410), .B(n409), .ZN(n536) );
  XNOR2_X2 U522 ( .A(n416), .B(n415), .ZN(n511) );
  XNOR2_X2 U523 ( .A(G101), .B(G110), .ZN(n415) );
  XNOR2_X2 U524 ( .A(n466), .B(G107), .ZN(n416) );
  XNOR2_X2 U525 ( .A(n539), .B(n538), .ZN(n546) );
  INV_X1 U526 ( .A(n546), .ZN(n420) );
  INV_X1 U527 ( .A(n567), .ZN(n424) );
  NAND2_X1 U528 ( .A1(n546), .A2(n360), .ZN(n426) );
  AND2_X2 U529 ( .A1(n745), .A2(n635), .ZN(n680) );
  INV_X1 U530 ( .A(KEYINPUT87), .ZN(n574) );
  INV_X1 U531 ( .A(KEYINPUT86), .ZN(n575) );
  NAND2_X1 U532 ( .A1(n568), .A2(n567), .ZN(n571) );
  BUF_X1 U533 ( .A(n677), .Z(n710) );
  AND2_X1 U534 ( .A1(n543), .A2(n682), .ZN(n552) );
  BUF_X1 U535 ( .A(n637), .Z(n640) );
  NAND2_X1 U536 ( .A1(G234), .A2(G237), .ZN(n427) );
  XNOR2_X1 U537 ( .A(n427), .B(KEYINPUT14), .ZN(n429) );
  NAND2_X1 U538 ( .A1(n429), .A2(G952), .ZN(n428) );
  XOR2_X1 U539 ( .A(KEYINPUT95), .B(n428), .Z(n716) );
  NOR2_X1 U540 ( .A1(G953), .A2(n716), .ZN(n531) );
  AND2_X1 U541 ( .A1(G953), .A2(n429), .ZN(n430) );
  NAND2_X1 U542 ( .A1(G902), .A2(n430), .ZN(n529) );
  XOR2_X1 U543 ( .A(n529), .B(KEYINPUT107), .Z(n431) );
  NOR2_X1 U544 ( .A1(G900), .A2(n431), .ZN(n432) );
  NOR2_X1 U545 ( .A1(n531), .A2(n432), .ZN(n517) );
  XOR2_X1 U546 ( .A(KEYINPUT5), .B(G101), .Z(n435) );
  NAND2_X1 U547 ( .A1(n488), .A2(G210), .ZN(n434) );
  XNOR2_X1 U548 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U549 ( .A(n468), .B(n436), .ZN(n439) );
  XNOR2_X1 U550 ( .A(n473), .B(n437), .ZN(n438) );
  XNOR2_X2 U551 ( .A(n504), .B(n438), .ZN(n759) );
  XNOR2_X1 U552 ( .A(n759), .B(n439), .ZN(n647) );
  NAND2_X1 U553 ( .A1(n647), .A2(n401), .ZN(n440) );
  NOR2_X1 U554 ( .A1(G902), .A2(G237), .ZN(n442) );
  INV_X1 U555 ( .A(KEYINPUT77), .ZN(n441) );
  XNOR2_X1 U556 ( .A(n442), .B(n441), .ZN(n477) );
  INV_X1 U557 ( .A(G214), .ZN(n443) );
  OR2_X1 U558 ( .A1(n477), .A2(n443), .ZN(n701) );
  NAND2_X1 U559 ( .A1(n687), .A2(n701), .ZN(n444) );
  XNOR2_X1 U560 ( .A(KEYINPUT30), .B(n444), .ZN(n445) );
  NOR2_X1 U561 ( .A1(n517), .A2(n445), .ZN(n465) );
  XNOR2_X1 U562 ( .A(G119), .B(G110), .ZN(n447) );
  XNOR2_X1 U563 ( .A(n358), .B(n447), .ZN(n448) );
  XNOR2_X1 U564 ( .A(n357), .B(n448), .ZN(n452) );
  XOR2_X1 U565 ( .A(KEYINPUT70), .B(KEYINPUT8), .Z(n450) );
  NAND2_X1 U566 ( .A1(G234), .A2(n761), .ZN(n449) );
  XNOR2_X1 U567 ( .A(n450), .B(n449), .ZN(n497) );
  NAND2_X1 U568 ( .A1(n497), .A2(G221), .ZN(n451) );
  XNOR2_X1 U569 ( .A(n452), .B(n451), .ZN(n454) );
  XNOR2_X1 U570 ( .A(G125), .B(KEYINPUT71), .ZN(n453) );
  XNOR2_X1 U571 ( .A(n348), .B(n453), .ZN(n758) );
  XOR2_X1 U572 ( .A(G146), .B(n758), .Z(n491) );
  XNOR2_X1 U573 ( .A(G902), .B(KEYINPUT93), .ZN(n456) );
  XNOR2_X1 U574 ( .A(n456), .B(n455), .ZN(n624) );
  NAND2_X1 U575 ( .A1(n624), .A2(G234), .ZN(n458) );
  XNOR2_X1 U576 ( .A(KEYINPUT98), .B(KEYINPUT20), .ZN(n457) );
  XNOR2_X1 U577 ( .A(n458), .B(n457), .ZN(n462) );
  NAND2_X1 U578 ( .A1(n462), .A2(G217), .ZN(n460) );
  NAND2_X1 U579 ( .A1(G221), .A2(n462), .ZN(n464) );
  XOR2_X1 U580 ( .A(KEYINPUT100), .B(KEYINPUT21), .Z(n463) );
  XNOR2_X1 U581 ( .A(n464), .B(n463), .ZN(n682) );
  BUF_X1 U582 ( .A(n552), .Z(n689) );
  NAND2_X1 U583 ( .A1(n465), .A2(n689), .ZN(n600) );
  INV_X1 U584 ( .A(n600), .ZN(n516) );
  INV_X2 U585 ( .A(G104), .ZN(n466) );
  NAND2_X1 U586 ( .A1(n761), .A2(G224), .ZN(n470) );
  XNOR2_X1 U587 ( .A(n470), .B(G125), .ZN(n471) );
  XNOR2_X1 U588 ( .A(n469), .B(n471), .ZN(n475) );
  XNOR2_X1 U589 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n472) );
  XNOR2_X1 U590 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U591 ( .A(n475), .B(n474), .ZN(n476) );
  INV_X1 U592 ( .A(n477), .ZN(n478) );
  NAND2_X1 U593 ( .A1(n478), .A2(G210), .ZN(n479) );
  XNOR2_X1 U594 ( .A(n479), .B(KEYINPUT94), .ZN(n480) );
  INV_X1 U595 ( .A(n601), .ZN(n614) );
  XNOR2_X1 U596 ( .A(n483), .B(n482), .ZN(n487) );
  XNOR2_X1 U597 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X1 U598 ( .A(n487), .B(n486), .Z(n490) );
  NAND2_X1 U599 ( .A1(G214), .A2(n488), .ZN(n489) );
  XNOR2_X1 U600 ( .A(n490), .B(n489), .ZN(n493) );
  INV_X1 U601 ( .A(n491), .ZN(n492) );
  XNOR2_X1 U602 ( .A(n493), .B(n492), .ZN(n730) );
  XNOR2_X1 U603 ( .A(KEYINPUT103), .B(KEYINPUT13), .ZN(n494) );
  XOR2_X1 U604 ( .A(KEYINPUT104), .B(KEYINPUT7), .Z(n499) );
  NAND2_X1 U605 ( .A1(G217), .A2(n497), .ZN(n498) );
  XNOR2_X1 U606 ( .A(n499), .B(n498), .ZN(n503) );
  XOR2_X1 U607 ( .A(KEYINPUT9), .B(G122), .Z(n501) );
  XNOR2_X1 U608 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U609 ( .A(n503), .B(n502), .ZN(n505) );
  XNOR2_X1 U610 ( .A(n504), .B(n505), .ZN(n738) );
  NAND2_X1 U611 ( .A1(n738), .A2(n401), .ZN(n507) );
  INV_X1 U612 ( .A(G478), .ZN(n506) );
  NOR2_X1 U613 ( .A1(n560), .A2(n534), .ZN(n572) );
  NAND2_X1 U614 ( .A1(n614), .A2(n572), .ZN(n514) );
  AND2_X1 U615 ( .A1(n761), .A2(G227), .ZN(n508) );
  XNOR2_X1 U616 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U617 ( .A(n356), .B(n510), .ZN(n512) );
  INV_X1 U618 ( .A(G469), .ZN(n513) );
  INV_X1 U619 ( .A(n522), .ZN(n588) );
  INV_X1 U620 ( .A(n588), .ZN(n599) );
  NOR2_X1 U621 ( .A1(n514), .A2(n599), .ZN(n515) );
  NAND2_X1 U622 ( .A1(n516), .A2(n515), .ZN(n593) );
  XNOR2_X1 U623 ( .A(n593), .B(G143), .ZN(G45) );
  NOR2_X1 U624 ( .A1(n517), .A2(n543), .ZN(n518) );
  NAND2_X1 U625 ( .A1(n682), .A2(n518), .ZN(n586) );
  INV_X1 U626 ( .A(n534), .ZN(n561) );
  OR2_X1 U627 ( .A1(n560), .A2(n561), .ZN(n667) );
  INV_X1 U628 ( .A(KEYINPUT6), .ZN(n519) );
  AND2_X1 U629 ( .A1(n663), .A2(n567), .ZN(n520) );
  NAND2_X1 U630 ( .A1(n520), .A2(n701), .ZN(n521) );
  NOR2_X1 U631 ( .A1(n586), .A2(n521), .ZN(n615) );
  NAND2_X1 U632 ( .A1(n615), .A2(n540), .ZN(n524) );
  XOR2_X1 U633 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n523) );
  XNOR2_X1 U634 ( .A(n524), .B(n523), .ZN(n525) );
  NOR2_X1 U635 ( .A1(n525), .A2(n614), .ZN(n630) );
  XOR2_X1 U636 ( .A(G140), .B(n630), .Z(G42) );
  INV_X1 U637 ( .A(n526), .ZN(n527) );
  NOR2_X1 U638 ( .A1(G898), .A2(n529), .ZN(n530) );
  OR2_X1 U639 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U640 ( .A(n532), .B(KEYINPUT96), .ZN(n533) );
  AND2_X1 U641 ( .A1(n704), .A2(n682), .ZN(n535) );
  NAND2_X1 U642 ( .A1(n536), .A2(n535), .ZN(n539) );
  XNOR2_X1 U643 ( .A(KEYINPUT75), .B(KEYINPUT22), .ZN(n537) );
  XNOR2_X1 U644 ( .A(n537), .B(KEYINPUT69), .ZN(n538) );
  XNOR2_X1 U645 ( .A(n543), .B(KEYINPUT105), .ZN(n684) );
  NAND2_X1 U646 ( .A1(n684), .A2(n367), .ZN(n541) );
  XNOR2_X1 U647 ( .A(KEYINPUT79), .B(KEYINPUT32), .ZN(n542) );
  XNOR2_X1 U648 ( .A(n364), .B(G119), .ZN(G21) );
  NOR2_X1 U649 ( .A1(n543), .A2(n375), .ZN(n544) );
  NAND2_X1 U650 ( .A1(n544), .A2(n540), .ZN(n545) );
  OR2_X1 U651 ( .A1(n546), .A2(n545), .ZN(n659) );
  NAND2_X1 U652 ( .A1(n547), .A2(n659), .ZN(n576) );
  NAND2_X1 U653 ( .A1(n576), .A2(KEYINPUT44), .ZN(n548) );
  XNOR2_X1 U654 ( .A(n548), .B(KEYINPUT67), .ZN(n565) );
  NOR2_X1 U655 ( .A1(n684), .A2(n367), .ZN(n549) );
  INV_X1 U656 ( .A(n687), .ZN(n585) );
  NOR2_X1 U657 ( .A1(n566), .A2(n585), .ZN(n554) );
  XNOR2_X1 U658 ( .A(n554), .B(KEYINPUT101), .ZN(n694) );
  NOR2_X1 U659 ( .A1(n694), .A2(n555), .ZN(n556) );
  XNOR2_X1 U660 ( .A(n556), .B(KEYINPUT31), .ZN(n669) );
  INV_X1 U661 ( .A(n555), .ZN(n559) );
  NAND2_X1 U662 ( .A1(n689), .A2(n588), .ZN(n557) );
  NOR2_X1 U663 ( .A1(n557), .A2(n375), .ZN(n558) );
  NAND2_X1 U664 ( .A1(n559), .A2(n558), .ZN(n654) );
  NAND2_X1 U665 ( .A1(n669), .A2(n654), .ZN(n562) );
  NAND2_X1 U666 ( .A1(n561), .A2(n560), .ZN(n670) );
  NAND2_X1 U667 ( .A1(n667), .A2(n670), .ZN(n700) );
  NAND2_X1 U668 ( .A1(n562), .A2(n700), .ZN(n563) );
  NAND2_X1 U669 ( .A1(n769), .A2(n563), .ZN(n564) );
  INV_X1 U670 ( .A(n566), .ZN(n568) );
  XNOR2_X1 U671 ( .A(KEYINPUT90), .B(KEYINPUT33), .ZN(n569) );
  XNOR2_X1 U672 ( .A(n569), .B(KEYINPUT73), .ZN(n570) );
  XNOR2_X1 U673 ( .A(KEYINPUT84), .B(KEYINPUT35), .ZN(n573) );
  BUF_X1 U674 ( .A(n576), .Z(n577) );
  XOR2_X1 U675 ( .A(KEYINPUT88), .B(n577), .Z(n581) );
  BUF_X1 U676 ( .A(n578), .Z(n579) );
  NOR2_X1 U677 ( .A1(n579), .A2(KEYINPUT44), .ZN(n580) );
  NAND2_X1 U678 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U679 ( .A(KEYINPUT83), .B(KEYINPUT45), .ZN(n583) );
  NOR2_X1 U680 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U681 ( .A(KEYINPUT28), .B(n587), .ZN(n589) );
  NAND2_X1 U682 ( .A1(n589), .A2(n588), .ZN(n609) );
  BUF_X1 U683 ( .A(n590), .Z(n591) );
  INV_X1 U684 ( .A(n591), .ZN(n592) );
  NAND2_X1 U685 ( .A1(n664), .A2(n700), .ZN(n596) );
  NAND2_X1 U686 ( .A1(n596), .A2(KEYINPUT47), .ZN(n594) );
  NAND2_X1 U687 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U688 ( .A(n595), .B(KEYINPUT82), .ZN(n598) );
  NOR2_X1 U689 ( .A1(KEYINPUT47), .A2(n596), .ZN(n597) );
  NOR2_X1 U690 ( .A1(n600), .A2(n599), .ZN(n602) );
  NAND2_X1 U691 ( .A1(n602), .A2(n702), .ZN(n604) );
  XNOR2_X1 U692 ( .A(KEYINPUT74), .B(KEYINPUT39), .ZN(n603) );
  XNOR2_X1 U693 ( .A(n604), .B(n603), .ZN(n620) );
  XOR2_X1 U694 ( .A(KEYINPUT41), .B(KEYINPUT110), .Z(n608) );
  NAND2_X1 U695 ( .A1(n702), .A2(n701), .ZN(n606) );
  NAND2_X1 U696 ( .A1(n704), .A2(n699), .ZN(n607) );
  XNOR2_X1 U697 ( .A(KEYINPUT42), .B(n610), .ZN(n770) );
  XNOR2_X1 U698 ( .A(n611), .B(KEYINPUT46), .ZN(n612) );
  NAND2_X1 U699 ( .A1(n615), .A2(n614), .ZN(n617) );
  XOR2_X1 U700 ( .A(KEYINPUT36), .B(KEYINPUT89), .Z(n616) );
  XNOR2_X1 U701 ( .A(n617), .B(n616), .ZN(n618) );
  XNOR2_X1 U702 ( .A(n619), .B(KEYINPUT48), .ZN(n628) );
  INV_X1 U703 ( .A(n670), .ZN(n660) );
  NAND2_X1 U704 ( .A1(n620), .A2(n660), .ZN(n675) );
  INV_X1 U705 ( .A(n675), .ZN(n621) );
  NOR2_X1 U706 ( .A1(n621), .A2(n630), .ZN(n622) );
  NAND2_X1 U707 ( .A1(n628), .A2(n622), .ZN(n760) );
  NOR2_X1 U708 ( .A1(n627), .A2(n760), .ZN(n623) );
  INV_X1 U709 ( .A(n624), .ZN(n625) );
  XNOR2_X2 U710 ( .A(n626), .B(KEYINPUT66), .ZN(n636) );
  INV_X1 U711 ( .A(n355), .ZN(n745) );
  INV_X1 U712 ( .A(n628), .ZN(n634) );
  NAND2_X1 U713 ( .A1(KEYINPUT2), .A2(n675), .ZN(n629) );
  XOR2_X1 U714 ( .A(KEYINPUT80), .B(n629), .Z(n632) );
  INV_X1 U715 ( .A(n630), .ZN(n631) );
  NAND2_X1 U716 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U717 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U718 ( .A(KEYINPUT81), .B(KEYINPUT54), .ZN(n638) );
  XOR2_X1 U719 ( .A(n638), .B(KEYINPUT55), .Z(n639) );
  XNOR2_X1 U720 ( .A(n642), .B(n641), .ZN(n644) );
  INV_X1 U721 ( .A(G952), .ZN(n643) );
  NOR2_X2 U722 ( .A1(n644), .A2(n744), .ZN(n646) );
  XNOR2_X1 U723 ( .A(KEYINPUT120), .B(KEYINPUT56), .ZN(n645) );
  XNOR2_X1 U724 ( .A(n646), .B(n645), .ZN(G51) );
  XNOR2_X1 U725 ( .A(n649), .B(n648), .ZN(n650) );
  NOR2_X2 U726 ( .A1(n650), .A2(n744), .ZN(n652) );
  XOR2_X1 U727 ( .A(KEYINPUT92), .B(KEYINPUT63), .Z(n651) );
  XNOR2_X1 U728 ( .A(n652), .B(n651), .ZN(G57) );
  XOR2_X1 U729 ( .A(n579), .B(G122), .Z(G24) );
  NOR2_X1 U730 ( .A1(n667), .A2(n654), .ZN(n653) );
  XOR2_X1 U731 ( .A(n362), .B(n653), .Z(G6) );
  NOR2_X1 U732 ( .A1(n654), .A2(n670), .ZN(n658) );
  XOR2_X1 U733 ( .A(KEYINPUT27), .B(KEYINPUT111), .Z(n656) );
  XNOR2_X1 U734 ( .A(G107), .B(KEYINPUT26), .ZN(n655) );
  XNOR2_X1 U735 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U736 ( .A(n658), .B(n657), .ZN(G9) );
  XNOR2_X1 U737 ( .A(G110), .B(n659), .ZN(G12) );
  XOR2_X1 U738 ( .A(G128), .B(KEYINPUT29), .Z(n662) );
  NAND2_X1 U739 ( .A1(n664), .A2(n660), .ZN(n661) );
  XNOR2_X1 U740 ( .A(n662), .B(n661), .ZN(G30) );
  XNOR2_X1 U741 ( .A(G146), .B(KEYINPUT112), .ZN(n666) );
  NAND2_X1 U742 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U743 ( .A(n666), .B(n665), .ZN(G48) );
  NOR2_X1 U744 ( .A1(n667), .A2(n669), .ZN(n668) );
  XOR2_X1 U745 ( .A(G113), .B(n668), .Z(G15) );
  NOR2_X1 U746 ( .A1(n670), .A2(n669), .ZN(n672) );
  XNOR2_X1 U747 ( .A(G116), .B(KEYINPUT113), .ZN(n671) );
  XNOR2_X1 U748 ( .A(n672), .B(n671), .ZN(G18) );
  XNOR2_X1 U749 ( .A(n673), .B(G125), .ZN(n674) );
  XNOR2_X1 U750 ( .A(n674), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U751 ( .A(G134), .B(n675), .ZN(G36) );
  NOR2_X1 U752 ( .A1(n698), .A2(n710), .ZN(n678) );
  XOR2_X1 U753 ( .A(KEYINPUT118), .B(n678), .Z(n720) );
  INV_X1 U754 ( .A(n679), .ZN(n681) );
  NOR2_X1 U755 ( .A1(n681), .A2(n680), .ZN(n718) );
  INV_X1 U756 ( .A(n682), .ZN(n683) );
  NAND2_X1 U757 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U758 ( .A(KEYINPUT49), .B(n685), .ZN(n686) );
  NOR2_X1 U759 ( .A1(n375), .A2(n686), .ZN(n688) );
  XNOR2_X1 U760 ( .A(n688), .B(KEYINPUT114), .ZN(n693) );
  NOR2_X1 U761 ( .A1(n367), .A2(n689), .ZN(n691) );
  XOR2_X1 U762 ( .A(KEYINPUT50), .B(n691), .Z(n692) );
  NAND2_X1 U763 ( .A1(n693), .A2(n692), .ZN(n695) );
  NAND2_X1 U764 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U765 ( .A(KEYINPUT51), .B(n696), .ZN(n697) );
  NOR2_X1 U766 ( .A1(n698), .A2(n697), .ZN(n712) );
  NAND2_X1 U767 ( .A1(n700), .A2(n699), .ZN(n708) );
  NOR2_X1 U768 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U769 ( .A(KEYINPUT115), .B(n703), .ZN(n705) );
  NAND2_X1 U770 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U771 ( .A(KEYINPUT116), .B(n706), .ZN(n707) );
  AND2_X1 U772 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U773 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U774 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U775 ( .A(n713), .B(KEYINPUT52), .Z(n714) );
  XNOR2_X1 U776 ( .A(KEYINPUT117), .B(n714), .ZN(n715) );
  NOR2_X1 U777 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U778 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U779 ( .A(KEYINPUT53), .B(n722), .ZN(G75) );
  XNOR2_X1 U780 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n723) );
  XNOR2_X1 U781 ( .A(n723), .B(KEYINPUT57), .ZN(n724) );
  XNOR2_X1 U782 ( .A(n727), .B(n726), .ZN(n728) );
  NOR2_X2 U783 ( .A1(n728), .A2(n744), .ZN(n729) );
  XNOR2_X1 U784 ( .A(n729), .B(KEYINPUT122), .ZN(G54) );
  XOR2_X1 U785 ( .A(KEYINPUT91), .B(KEYINPUT123), .Z(n732) );
  XNOR2_X1 U786 ( .A(n730), .B(KEYINPUT59), .ZN(n731) );
  XNOR2_X1 U787 ( .A(n734), .B(n733), .ZN(n735) );
  NOR2_X2 U788 ( .A1(n735), .A2(n744), .ZN(n736) );
  XNOR2_X1 U789 ( .A(n736), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U790 ( .A(n738), .B(n737), .Z(n739) );
  NOR2_X1 U791 ( .A1(n744), .A2(n739), .ZN(G63) );
  NAND2_X1 U792 ( .A1(n740), .A2(G217), .ZN(n742) );
  XNOR2_X1 U793 ( .A(n742), .B(n741), .ZN(n743) );
  NOR2_X1 U794 ( .A1(n744), .A2(n743), .ZN(G66) );
  NAND2_X1 U795 ( .A1(n745), .A2(n761), .ZN(n749) );
  NAND2_X1 U796 ( .A1(G953), .A2(G224), .ZN(n746) );
  XNOR2_X1 U797 ( .A(KEYINPUT61), .B(n746), .ZN(n747) );
  NAND2_X1 U798 ( .A1(n747), .A2(G898), .ZN(n748) );
  NAND2_X1 U799 ( .A1(n749), .A2(n748), .ZN(n756) );
  NOR2_X1 U800 ( .A1(G898), .A2(n761), .ZN(n753) );
  BUF_X1 U801 ( .A(n750), .Z(n751) );
  XOR2_X1 U802 ( .A(n751), .B(KEYINPUT125), .Z(n752) );
  NOR2_X1 U803 ( .A1(n753), .A2(n752), .ZN(n754) );
  XOR2_X1 U804 ( .A(KEYINPUT124), .B(n754), .Z(n755) );
  XNOR2_X1 U805 ( .A(n756), .B(n755), .ZN(n757) );
  XOR2_X1 U806 ( .A(KEYINPUT126), .B(n757), .Z(G69) );
  XNOR2_X1 U807 ( .A(n759), .B(n758), .ZN(n763) );
  XNOR2_X1 U808 ( .A(n760), .B(n763), .ZN(n762) );
  NAND2_X1 U809 ( .A1(n762), .A2(n761), .ZN(n768) );
  XNOR2_X1 U810 ( .A(n763), .B(G227), .ZN(n764) );
  NAND2_X1 U811 ( .A1(n764), .A2(G900), .ZN(n765) );
  XOR2_X1 U812 ( .A(KEYINPUT127), .B(n765), .Z(n766) );
  NAND2_X1 U813 ( .A1(G953), .A2(n766), .ZN(n767) );
  NAND2_X1 U814 ( .A1(n768), .A2(n767), .ZN(G72) );
  XNOR2_X1 U815 ( .A(n363), .B(G101), .ZN(G3) );
  XOR2_X1 U816 ( .A(G137), .B(n770), .Z(G39) );
  XOR2_X1 U817 ( .A(G131), .B(n771), .Z(G33) );
endmodule

