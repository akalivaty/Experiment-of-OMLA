

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757;

  AND2_X1 U370 ( .A1(n733), .A2(n362), .ZN(n593) );
  XNOR2_X1 U371 ( .A(n655), .B(n471), .ZN(n499) );
  XNOR2_X2 U372 ( .A(n349), .B(n626), .ZN(n683) );
  NAND2_X1 U373 ( .A1(n654), .A2(n415), .ZN(n349) );
  AND2_X1 U374 ( .A1(n652), .A2(n567), .ZN(n423) );
  XNOR2_X1 U375 ( .A(n418), .B(n605), .ZN(n713) );
  XNOR2_X1 U376 ( .A(G131), .B(KEYINPUT73), .ZN(n446) );
  XNOR2_X1 U377 ( .A(n403), .B(KEYINPUT32), .ZN(n579) );
  XNOR2_X1 U378 ( .A(n594), .B(KEYINPUT114), .ZN(n416) );
  XNOR2_X1 U379 ( .A(n419), .B(KEYINPUT112), .ZN(n401) );
  XNOR2_X1 U380 ( .A(n515), .B(n470), .ZN(n655) );
  XNOR2_X1 U381 ( .A(n468), .B(n467), .ZN(n515) );
  XNOR2_X1 U382 ( .A(n446), .B(KEYINPUT72), .ZN(n469) );
  XNOR2_X1 U383 ( .A(n571), .B(n538), .ZN(n350) );
  BUF_X1 U384 ( .A(n675), .Z(n351) );
  NAND2_X1 U385 ( .A1(n501), .A2(n500), .ZN(n354) );
  NAND2_X1 U386 ( .A1(n352), .A2(n353), .ZN(n355) );
  NAND2_X2 U387 ( .A1(n354), .A2(n355), .ZN(n571) );
  INV_X1 U388 ( .A(n501), .ZN(n352) );
  INV_X1 U389 ( .A(n500), .ZN(n353) );
  XNOR2_X1 U390 ( .A(n571), .B(n538), .ZN(n560) );
  NOR2_X2 U391 ( .A1(n618), .A2(n619), .ZN(n369) );
  BUF_X1 U392 ( .A(n630), .Z(n356) );
  XNOR2_X1 U393 ( .A(n499), .B(n498), .ZN(n630) );
  AND2_X1 U394 ( .A1(n675), .A2(G472), .ZN(n632) );
  XNOR2_X1 U395 ( .A(n609), .B(KEYINPUT85), .ZN(n612) );
  INV_X1 U396 ( .A(KEYINPUT47), .ZN(n398) );
  NOR2_X1 U397 ( .A1(n600), .A2(n541), .ZN(n586) );
  XNOR2_X1 U398 ( .A(G113), .B(KEYINPUT75), .ZN(n492) );
  XNOR2_X1 U399 ( .A(n469), .B(G134), .ZN(n470) );
  INV_X1 U400 ( .A(KEYINPUT0), .ZN(n365) );
  NAND2_X1 U401 ( .A1(n401), .A2(n700), .ZN(n418) );
  NOR2_X1 U402 ( .A1(n506), .A2(n551), .ZN(n602) );
  INV_X1 U403 ( .A(n364), .ZN(n549) );
  INV_X1 U404 ( .A(n392), .ZN(n689) );
  NAND2_X1 U405 ( .A1(n375), .A2(n685), .ZN(n596) );
  XNOR2_X1 U406 ( .A(n377), .B(n376), .ZN(n375) );
  INV_X1 U407 ( .A(KEYINPUT36), .ZN(n376) );
  NAND2_X1 U408 ( .A1(n416), .A2(n357), .ZN(n377) );
  XNOR2_X1 U409 ( .A(G113), .B(G143), .ZN(n452) );
  INV_X1 U410 ( .A(KEYINPUT88), .ZN(n367) );
  XNOR2_X1 U411 ( .A(n436), .B(n435), .ZN(n479) );
  XNOR2_X1 U412 ( .A(n512), .B(n458), .ZN(n480) );
  INV_X1 U413 ( .A(KEYINPUT10), .ZN(n458) );
  XOR2_X1 U414 ( .A(KEYINPUT96), .B(KEYINPUT11), .Z(n448) );
  XNOR2_X1 U415 ( .A(KEYINPUT71), .B(G101), .ZN(n509) );
  XNOR2_X1 U416 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n511) );
  XNOR2_X1 U417 ( .A(KEYINPUT66), .B(KEYINPUT4), .ZN(n467) );
  AND2_X1 U418 ( .A1(n543), .A2(n732), .ZN(n594) );
  XNOR2_X1 U419 ( .A(n379), .B(n378), .ZN(n543) );
  INV_X1 U420 ( .A(G902), .ZN(n503) );
  NOR2_X1 U421 ( .A1(G902), .A2(n677), .ZN(n478) );
  XNOR2_X1 U422 ( .A(G128), .B(KEYINPUT23), .ZN(n482) );
  XNOR2_X1 U423 ( .A(n480), .B(n481), .ZN(n656) );
  XNOR2_X1 U424 ( .A(n483), .B(n360), .ZN(n395) );
  XOR2_X1 U425 ( .A(KEYINPUT7), .B(G122), .Z(n441) );
  XNOR2_X1 U426 ( .A(G116), .B(G107), .ZN(n440) );
  XOR2_X1 U427 ( .A(G137), .B(G140), .Z(n481) );
  XNOR2_X1 U428 ( .A(n366), .B(n472), .ZN(n519) );
  INV_X1 U429 ( .A(G104), .ZN(n472) );
  XNOR2_X1 U430 ( .A(G110), .B(G107), .ZN(n366) );
  XNOR2_X1 U431 ( .A(n370), .B(KEYINPUT45), .ZN(n415) );
  NAND2_X1 U432 ( .A1(n381), .A2(n382), .ZN(n370) );
  NOR2_X1 U433 ( .A1(n385), .A2(n386), .ZN(n382) );
  XNOR2_X1 U434 ( .A(n407), .B(n406), .ZN(n622) );
  XNOR2_X1 U435 ( .A(n603), .B(KEYINPUT39), .ZN(n406) );
  NAND2_X1 U436 ( .A1(n602), .A2(n601), .ZN(n407) );
  NAND2_X1 U437 ( .A1(n698), .A2(KEYINPUT19), .ZN(n414) );
  INV_X1 U438 ( .A(KEYINPUT104), .ZN(n569) );
  XNOR2_X1 U439 ( .A(n396), .B(n393), .ZN(n667) );
  XNOR2_X1 U440 ( .A(n395), .B(n394), .ZN(n393) );
  XNOR2_X1 U441 ( .A(n397), .B(n656), .ZN(n396) );
  XNOR2_X1 U442 ( .A(n482), .B(KEYINPUT89), .ZN(n394) );
  INV_X1 U443 ( .A(KEYINPUT68), .ZN(n417) );
  NAND2_X1 U444 ( .A1(n683), .A2(n629), .ZN(n372) );
  XNOR2_X1 U445 ( .A(n607), .B(KEYINPUT42), .ZN(n400) );
  INV_X1 U446 ( .A(KEYINPUT35), .ZN(n368) );
  NOR2_X1 U447 ( .A1(n539), .A2(n540), .ZN(n403) );
  NOR2_X1 U448 ( .A1(n549), .A2(n404), .ZN(n550) );
  AND2_X1 U449 ( .A1(n602), .A2(n383), .ZN(n609) );
  AND2_X1 U450 ( .A1(n507), .A2(n384), .ZN(n383) );
  NOR2_X1 U451 ( .A1(n555), .A2(n599), .ZN(n384) );
  INV_X1 U452 ( .A(KEYINPUT87), .ZN(n408) );
  NOR2_X1 U453 ( .A1(n539), .A2(n685), .ZN(n388) );
  INV_X1 U454 ( .A(n596), .ZN(n741) );
  AND2_X1 U455 ( .A1(n413), .A2(n544), .ZN(n357) );
  XNOR2_X1 U456 ( .A(KEYINPUT25), .B(n486), .ZN(n358) );
  AND2_X1 U457 ( .A1(n700), .A2(n428), .ZN(n359) );
  XOR2_X1 U458 ( .A(G119), .B(G110), .Z(n360) );
  NOR2_X1 U459 ( .A1(n553), .A2(n559), .ZN(n361) );
  AND2_X1 U460 ( .A1(n702), .A2(n398), .ZN(n362) );
  NAND2_X1 U461 ( .A1(n410), .A2(n409), .ZN(n363) );
  NAND2_X1 U462 ( .A1(n410), .A2(n409), .ZN(n420) );
  NAND2_X1 U463 ( .A1(n413), .A2(n412), .ZN(n409) );
  XNOR2_X2 U464 ( .A(n431), .B(G953), .ZN(n508) );
  BUF_X1 U465 ( .A(n508), .Z(n660) );
  NOR2_X1 U466 ( .A1(n423), .A2(n422), .ZN(n421) );
  NAND2_X1 U467 ( .A1(n420), .A2(n533), .ZN(n534) );
  BUF_X1 U468 ( .A(n571), .Z(n553) );
  NAND2_X1 U469 ( .A1(n374), .A2(n361), .ZN(n404) );
  NOR2_X1 U470 ( .A1(n350), .A2(n380), .ZN(n379) );
  XNOR2_X2 U471 ( .A(n534), .B(n365), .ZN(n364) );
  NAND2_X1 U472 ( .A1(n580), .A2(n367), .ZN(n578) );
  OR2_X2 U473 ( .A1(n580), .A2(n367), .ZN(n424) );
  XNOR2_X1 U474 ( .A(n580), .B(G122), .ZN(G24) );
  XNOR2_X2 U475 ( .A(n566), .B(n368), .ZN(n580) );
  XNOR2_X2 U476 ( .A(n592), .B(KEYINPUT111), .ZN(n606) );
  XNOR2_X1 U477 ( .A(n369), .B(KEYINPUT48), .ZN(n625) );
  NOR2_X2 U478 ( .A1(n699), .A2(n698), .ZN(n419) );
  XNOR2_X1 U479 ( .A(n388), .B(n408), .ZN(n371) );
  NAND2_X1 U480 ( .A1(n577), .A2(n578), .ZN(n385) );
  NAND2_X1 U481 ( .A1(n371), .A2(n689), .ZN(n556) );
  INV_X1 U482 ( .A(n595), .ZN(n374) );
  NAND2_X1 U483 ( .A1(n725), .A2(n738), .ZN(n391) );
  NAND2_X1 U484 ( .A1(n387), .A2(n585), .ZN(n381) );
  XNOR2_X2 U485 ( .A(n372), .B(n417), .ZN(n675) );
  INV_X1 U486 ( .A(KEYINPUT107), .ZN(n378) );
  INV_X1 U487 ( .A(n586), .ZN(n380) );
  INV_X1 U488 ( .A(n415), .ZN(n748) );
  XNOR2_X1 U489 ( .A(n558), .B(n557), .ZN(n386) );
  NAND2_X1 U490 ( .A1(n424), .A2(n421), .ZN(n387) );
  NAND2_X1 U491 ( .A1(n389), .A2(n556), .ZN(n558) );
  NAND2_X1 U492 ( .A1(n390), .A2(n702), .ZN(n389) );
  XNOR2_X1 U493 ( .A(n391), .B(KEYINPUT94), .ZN(n390) );
  NAND2_X1 U494 ( .A1(n392), .A2(n428), .ZN(n541) );
  XNOR2_X2 U495 ( .A(n487), .B(n358), .ZN(n392) );
  NAND2_X1 U496 ( .A1(n685), .A2(n392), .ZN(n540) );
  NAND2_X1 U497 ( .A1(n479), .A2(G221), .ZN(n397) );
  XNOR2_X2 U498 ( .A(n399), .B(KEYINPUT83), .ZN(n733) );
  NAND2_X1 U499 ( .A1(n606), .A2(n363), .ZN(n399) );
  NAND2_X1 U500 ( .A1(n400), .A2(n757), .ZN(n608) );
  XNOR2_X1 U501 ( .A(n400), .B(G137), .ZN(G39) );
  NAND2_X1 U502 ( .A1(n401), .A2(n702), .ZN(n703) );
  NAND2_X1 U503 ( .A1(n402), .A2(KEYINPUT44), .ZN(n422) );
  NAND2_X1 U504 ( .A1(n579), .A2(n567), .ZN(n402) );
  NAND2_X1 U505 ( .A1(n693), .A2(n404), .ZN(n694) );
  NOR2_X1 U506 ( .A1(n405), .A2(n595), .ZN(n561) );
  XNOR2_X2 U507 ( .A(n589), .B(n527), .ZN(n595) );
  XNOR2_X2 U508 ( .A(n478), .B(n477), .ZN(n589) );
  OR2_X2 U509 ( .A1(n560), .A2(n559), .ZN(n405) );
  AND2_X2 U510 ( .A1(n411), .A2(n414), .ZN(n410) );
  INV_X1 U511 ( .A(n528), .ZN(n413) );
  NAND2_X1 U512 ( .A1(n528), .A2(KEYINPUT19), .ZN(n411) );
  NOR2_X1 U513 ( .A1(n698), .A2(KEYINPUT19), .ZN(n412) );
  XNOR2_X2 U514 ( .A(n526), .B(n525), .ZN(n528) );
  AND2_X2 U515 ( .A1(n625), .A2(n426), .ZN(n654) );
  AND2_X1 U516 ( .A1(n675), .A2(G475), .ZN(n641) );
  AND2_X1 U517 ( .A1(n675), .A2(G210), .ZN(n649) );
  AND2_X1 U518 ( .A1(n351), .A2(G217), .ZN(n668) );
  AND2_X1 U519 ( .A1(n351), .A2(G478), .ZN(n673) );
  NOR2_X1 U520 ( .A1(n652), .A2(n579), .ZN(n584) );
  XNOR2_X2 U521 ( .A(n599), .B(n598), .ZN(n699) );
  AND2_X1 U522 ( .A1(n616), .A2(n615), .ZN(n425) );
  AND2_X1 U523 ( .A1(n624), .A2(n623), .ZN(n426) );
  XNOR2_X1 U524 ( .A(KEYINPUT65), .B(KEYINPUT46), .ZN(n427) );
  XOR2_X1 U525 ( .A(n490), .B(n489), .Z(n428) );
  INV_X1 U526 ( .A(KEYINPUT103), .ZN(n557) );
  XNOR2_X1 U527 ( .A(n608), .B(n427), .ZN(n617) );
  INV_X1 U528 ( .A(G469), .ZN(n476) );
  XNOR2_X1 U529 ( .A(n476), .B(KEYINPUT74), .ZN(n477) );
  XNOR2_X1 U530 ( .A(n505), .B(KEYINPUT30), .ZN(n506) );
  XNOR2_X1 U531 ( .A(KEYINPUT86), .B(KEYINPUT76), .ZN(n603) );
  XNOR2_X1 U532 ( .A(n604), .B(KEYINPUT40), .ZN(n757) );
  NAND2_X1 U533 ( .A1(G234), .A2(G237), .ZN(n429) );
  XNOR2_X1 U534 ( .A(n429), .B(KEYINPUT14), .ZN(n430) );
  NAND2_X1 U535 ( .A1(G952), .A2(n430), .ZN(n710) );
  NOR2_X1 U536 ( .A1(n710), .A2(G953), .ZN(n532) );
  NAND2_X1 U537 ( .A1(G902), .A2(n430), .ZN(n530) );
  NOR2_X1 U538 ( .A1(G900), .A2(n530), .ZN(n432) );
  INV_X2 U539 ( .A(KEYINPUT64), .ZN(n431) );
  INV_X1 U540 ( .A(n660), .ZN(n634) );
  NAND2_X1 U541 ( .A1(n432), .A2(n634), .ZN(n433) );
  XOR2_X1 U542 ( .A(KEYINPUT106), .B(n433), .Z(n434) );
  NOR2_X1 U543 ( .A1(n532), .A2(n434), .ZN(n600) );
  XOR2_X1 U544 ( .A(G134), .B(KEYINPUT9), .Z(n438) );
  NAND2_X1 U545 ( .A1(n508), .A2(G234), .ZN(n436) );
  INV_X1 U546 ( .A(KEYINPUT8), .ZN(n435) );
  NAND2_X1 U547 ( .A1(G217), .A2(n479), .ZN(n437) );
  XNOR2_X1 U548 ( .A(n438), .B(n437), .ZN(n444) );
  XNOR2_X2 U549 ( .A(G128), .B(KEYINPUT67), .ZN(n439) );
  XNOR2_X2 U550 ( .A(n439), .B(G143), .ZN(n468) );
  XNOR2_X1 U551 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U552 ( .A(n468), .B(n442), .ZN(n443) );
  XNOR2_X1 U553 ( .A(n444), .B(n443), .ZN(n671) );
  NAND2_X1 U554 ( .A1(n671), .A2(n503), .ZN(n445) );
  INV_X1 U555 ( .A(G478), .ZN(n670) );
  XNOR2_X1 U556 ( .A(n445), .B(n670), .ZN(n620) );
  NOR2_X1 U557 ( .A1(n600), .A2(n620), .ZN(n507) );
  XNOR2_X1 U558 ( .A(KEYINPUT97), .B(KEYINPUT99), .ZN(n447) );
  XNOR2_X1 U559 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U560 ( .A(n469), .B(n449), .Z(n451) );
  NOR2_X1 U561 ( .A1(G953), .A2(G237), .ZN(n494) );
  NAND2_X1 U562 ( .A1(G214), .A2(n494), .ZN(n450) );
  XNOR2_X1 U563 ( .A(n451), .B(n450), .ZN(n462) );
  XOR2_X1 U564 ( .A(G122), .B(G104), .Z(n453) );
  XNOR2_X1 U565 ( .A(n453), .B(n452), .ZN(n457) );
  XOR2_X1 U566 ( .A(KEYINPUT95), .B(KEYINPUT98), .Z(n455) );
  XNOR2_X1 U567 ( .A(G140), .B(KEYINPUT12), .ZN(n454) );
  XNOR2_X1 U568 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U569 ( .A(n457), .B(n456), .ZN(n460) );
  XNOR2_X2 U570 ( .A(G146), .B(G125), .ZN(n512) );
  INV_X1 U571 ( .A(n480), .ZN(n459) );
  XNOR2_X1 U572 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U573 ( .A(n462), .B(n461), .ZN(n639) );
  NAND2_X1 U574 ( .A1(n639), .A2(n503), .ZN(n466) );
  XOR2_X1 U575 ( .A(KEYINPUT13), .B(KEYINPUT101), .Z(n464) );
  XNOR2_X1 U576 ( .A(KEYINPUT100), .B(G475), .ZN(n463) );
  XNOR2_X1 U577 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U578 ( .A(n466), .B(n465), .ZN(n555) );
  INV_X1 U579 ( .A(n555), .ZN(n621) );
  XNOR2_X1 U580 ( .A(n509), .B(G146), .ZN(n471) );
  NAND2_X1 U581 ( .A1(n660), .A2(G227), .ZN(n473) );
  XNOR2_X1 U582 ( .A(n519), .B(n473), .ZN(n474) );
  XNOR2_X1 U583 ( .A(n481), .B(n474), .ZN(n475) );
  XNOR2_X1 U584 ( .A(n499), .B(n475), .ZN(n677) );
  XOR2_X1 U585 ( .A(KEYINPUT90), .B(KEYINPUT24), .Z(n483) );
  NAND2_X1 U586 ( .A1(n667), .A2(n503), .ZN(n487) );
  XOR2_X1 U587 ( .A(KEYINPUT20), .B(KEYINPUT91), .Z(n485) );
  XNOR2_X1 U588 ( .A(KEYINPUT15), .B(G902), .ZN(n523) );
  NAND2_X1 U589 ( .A1(G234), .A2(n523), .ZN(n484) );
  XNOR2_X1 U590 ( .A(n485), .B(n484), .ZN(n488) );
  NAND2_X1 U591 ( .A1(G217), .A2(n488), .ZN(n486) );
  AND2_X1 U592 ( .A1(n488), .A2(G221), .ZN(n490) );
  INV_X1 U593 ( .A(KEYINPUT21), .ZN(n489) );
  NAND2_X1 U594 ( .A1(n689), .A2(n428), .ZN(n559) );
  INV_X1 U595 ( .A(n559), .ZN(n684) );
  NAND2_X1 U596 ( .A1(n589), .A2(n684), .ZN(n551) );
  XNOR2_X1 U597 ( .A(G119), .B(G116), .ZN(n491) );
  XNOR2_X1 U598 ( .A(n491), .B(KEYINPUT3), .ZN(n493) );
  XNOR2_X1 U599 ( .A(n493), .B(n492), .ZN(n521) );
  XOR2_X1 U600 ( .A(G137), .B(KEYINPUT5), .Z(n496) );
  NAND2_X1 U601 ( .A1(n494), .A2(G210), .ZN(n495) );
  XNOR2_X1 U602 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U603 ( .A(n521), .B(n497), .ZN(n498) );
  NAND2_X1 U604 ( .A1(n630), .A2(n503), .ZN(n501) );
  XNOR2_X1 U605 ( .A(G472), .B(KEYINPUT93), .ZN(n500) );
  INV_X1 U606 ( .A(n571), .ZN(n504) );
  INV_X1 U607 ( .A(G237), .ZN(n502) );
  NAND2_X1 U608 ( .A1(n503), .A2(n502), .ZN(n524) );
  NAND2_X1 U609 ( .A1(n524), .A2(G214), .ZN(n544) );
  NAND2_X1 U610 ( .A1(n504), .A2(n544), .ZN(n505) );
  NAND2_X1 U611 ( .A1(n508), .A2(G224), .ZN(n510) );
  XNOR2_X1 U612 ( .A(n510), .B(n509), .ZN(n514) );
  XNOR2_X1 U613 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U614 ( .A(n514), .B(n513), .ZN(n516) );
  XNOR2_X1 U615 ( .A(n516), .B(n515), .ZN(n522) );
  XNOR2_X1 U616 ( .A(KEYINPUT78), .B(KEYINPUT16), .ZN(n517) );
  XNOR2_X1 U617 ( .A(n517), .B(G122), .ZN(n518) );
  XNOR2_X1 U618 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U619 ( .A(n521), .B(n520), .ZN(n745) );
  XNOR2_X1 U620 ( .A(n522), .B(n745), .ZN(n645) );
  INV_X1 U621 ( .A(n523), .ZN(n628) );
  OR2_X2 U622 ( .A1(n645), .A2(n628), .ZN(n526) );
  NAND2_X1 U623 ( .A1(n524), .A2(G210), .ZN(n525) );
  BUF_X2 U624 ( .A(n528), .Z(n599) );
  XOR2_X1 U625 ( .A(G143), .B(n609), .Z(G45) );
  INV_X1 U626 ( .A(KEYINPUT1), .ZN(n527) );
  INV_X1 U627 ( .A(n595), .ZN(n685) );
  INV_X1 U628 ( .A(n544), .ZN(n698) );
  INV_X1 U629 ( .A(G898), .ZN(n529) );
  NAND2_X1 U630 ( .A1(G953), .A2(n529), .ZN(n746) );
  NOR2_X1 U631 ( .A1(n530), .A2(n746), .ZN(n531) );
  OR2_X1 U632 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U633 ( .A1(n620), .A2(n555), .ZN(n700) );
  NAND2_X1 U634 ( .A1(n364), .A2(n359), .ZN(n536) );
  XNOR2_X1 U635 ( .A(KEYINPUT77), .B(KEYINPUT22), .ZN(n535) );
  XNOR2_X1 U636 ( .A(n536), .B(n535), .ZN(n568) );
  INV_X1 U637 ( .A(KEYINPUT102), .ZN(n537) );
  XNOR2_X1 U638 ( .A(n537), .B(KEYINPUT6), .ZN(n538) );
  NAND2_X1 U639 ( .A1(n568), .A2(n350), .ZN(n539) );
  XNOR2_X1 U640 ( .A(n556), .B(G101), .ZN(G3) );
  XOR2_X1 U641 ( .A(G119), .B(n579), .Z(G21) );
  INV_X1 U642 ( .A(n620), .ZN(n542) );
  NOR2_X1 U643 ( .A1(n542), .A2(n555), .ZN(n732) );
  NAND2_X1 U644 ( .A1(n594), .A2(n544), .ZN(n545) );
  XOR2_X1 U645 ( .A(KEYINPUT108), .B(n545), .Z(n546) );
  NAND2_X1 U646 ( .A1(n546), .A2(n595), .ZN(n547) );
  XNOR2_X1 U647 ( .A(n547), .B(KEYINPUT43), .ZN(n548) );
  NAND2_X1 U648 ( .A1(n548), .A2(n599), .ZN(n623) );
  XNOR2_X1 U649 ( .A(n623), .B(G140), .ZN(G42) );
  XNOR2_X1 U650 ( .A(n550), .B(KEYINPUT31), .ZN(n738) );
  NOR2_X1 U651 ( .A1(n549), .A2(n551), .ZN(n552) );
  XNOR2_X1 U652 ( .A(KEYINPUT92), .B(n552), .ZN(n554) );
  NAND2_X1 U653 ( .A1(n554), .A2(n553), .ZN(n725) );
  NOR2_X1 U654 ( .A1(n555), .A2(n620), .ZN(n563) );
  OR2_X1 U655 ( .A1(n563), .A2(n700), .ZN(n610) );
  INV_X1 U656 ( .A(n610), .ZN(n702) );
  XNOR2_X1 U657 ( .A(n561), .B(KEYINPUT33), .ZN(n697) );
  NOR2_X1 U658 ( .A1(n697), .A2(n549), .ZN(n562) );
  XNOR2_X1 U659 ( .A(n562), .B(KEYINPUT34), .ZN(n565) );
  XNOR2_X1 U660 ( .A(KEYINPUT82), .B(n563), .ZN(n564) );
  NAND2_X1 U661 ( .A1(n565), .A2(n564), .ZN(n566) );
  INV_X1 U662 ( .A(KEYINPUT69), .ZN(n567) );
  NOR2_X1 U663 ( .A1(n579), .A2(n567), .ZN(n576) );
  NAND2_X1 U664 ( .A1(n568), .A2(n595), .ZN(n570) );
  XNOR2_X1 U665 ( .A(n570), .B(n569), .ZN(n573) );
  INV_X1 U666 ( .A(n571), .ZN(n688) );
  NOR2_X1 U667 ( .A1(n504), .A2(n689), .ZN(n572) );
  NAND2_X1 U668 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X2 U669 ( .A(n574), .B(KEYINPUT105), .ZN(n652) );
  INV_X1 U670 ( .A(n652), .ZN(n575) );
  NAND2_X1 U671 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U672 ( .A1(n580), .A2(n584), .ZN(n583) );
  NOR2_X1 U673 ( .A1(KEYINPUT69), .A2(KEYINPUT44), .ZN(n581) );
  AND2_X1 U674 ( .A1(n581), .A2(KEYINPUT88), .ZN(n582) );
  NAND2_X1 U675 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U676 ( .A1(n688), .A2(n586), .ZN(n588) );
  XOR2_X1 U677 ( .A(KEYINPUT110), .B(KEYINPUT28), .Z(n587) );
  XNOR2_X1 U678 ( .A(n588), .B(n587), .ZN(n591) );
  XOR2_X1 U679 ( .A(n589), .B(KEYINPUT109), .Z(n590) );
  NAND2_X1 U680 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U681 ( .A(n593), .B(KEYINPUT79), .ZN(n597) );
  NAND2_X1 U682 ( .A1(n597), .A2(n596), .ZN(n619) );
  XOR2_X1 U683 ( .A(KEYINPUT80), .B(KEYINPUT38), .Z(n598) );
  NOR2_X1 U684 ( .A1(n600), .A2(n699), .ZN(n601) );
  NAND2_X1 U685 ( .A1(n622), .A2(n732), .ZN(n604) );
  XOR2_X1 U686 ( .A(KEYINPUT113), .B(KEYINPUT41), .Z(n605) );
  NAND2_X1 U687 ( .A1(n713), .A2(n606), .ZN(n607) );
  NAND2_X1 U688 ( .A1(n610), .A2(KEYINPUT47), .ZN(n611) );
  NAND2_X1 U689 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U690 ( .A(KEYINPUT84), .B(n613), .Z(n616) );
  INV_X1 U691 ( .A(n733), .ZN(n614) );
  NAND2_X1 U692 ( .A1(KEYINPUT47), .A2(n614), .ZN(n615) );
  NAND2_X1 U693 ( .A1(n617), .A2(n425), .ZN(n618) );
  OR2_X1 U694 ( .A1(n621), .A2(n620), .ZN(n739) );
  INV_X1 U695 ( .A(n739), .ZN(n729) );
  AND2_X1 U696 ( .A1(n729), .A2(n622), .ZN(n743) );
  INV_X1 U697 ( .A(n743), .ZN(n624) );
  INV_X1 U698 ( .A(KEYINPUT2), .ZN(n627) );
  NOR2_X1 U699 ( .A1(n627), .A2(KEYINPUT81), .ZN(n626) );
  NAND2_X1 U700 ( .A1(n627), .A2(KEYINPUT81), .ZN(n682) );
  AND2_X1 U701 ( .A1(n682), .A2(n628), .ZN(n629) );
  XOR2_X1 U702 ( .A(KEYINPUT62), .B(n356), .Z(n631) );
  XNOR2_X1 U703 ( .A(n632), .B(n631), .ZN(n636) );
  INV_X1 U704 ( .A(G952), .ZN(n633) );
  AND2_X1 U705 ( .A1(n634), .A2(n633), .ZN(n680) );
  INV_X1 U706 ( .A(n680), .ZN(n635) );
  NAND2_X1 U707 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U708 ( .A(n637), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U709 ( .A(KEYINPUT122), .B(KEYINPUT59), .Z(n638) );
  XNOR2_X1 U710 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U711 ( .A(n641), .B(n640), .ZN(n642) );
  NOR2_X1 U712 ( .A1(n642), .A2(n680), .ZN(n644) );
  XNOR2_X1 U713 ( .A(KEYINPUT70), .B(KEYINPUT60), .ZN(n643) );
  XNOR2_X1 U714 ( .A(n644), .B(n643), .ZN(G60) );
  BUF_X1 U715 ( .A(n645), .Z(n646) );
  XNOR2_X1 U716 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n647) );
  XNOR2_X1 U717 ( .A(n646), .B(n647), .ZN(n648) );
  XNOR2_X1 U718 ( .A(n649), .B(n648), .ZN(n650) );
  NOR2_X1 U719 ( .A1(n650), .A2(n680), .ZN(n651) );
  XNOR2_X1 U720 ( .A(n651), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U721 ( .A(G110), .B(KEYINPUT116), .ZN(n653) );
  XOR2_X1 U722 ( .A(n653), .B(n652), .Z(G12) );
  INV_X1 U723 ( .A(n654), .ZN(n659) );
  BUF_X1 U724 ( .A(n655), .Z(n657) );
  XNOR2_X1 U725 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U726 ( .A(n658), .B(KEYINPUT127), .ZN(n662) );
  XNOR2_X1 U727 ( .A(n659), .B(n662), .ZN(n661) );
  NAND2_X1 U728 ( .A1(n661), .A2(n660), .ZN(n666) );
  XNOR2_X1 U729 ( .A(G227), .B(n662), .ZN(n663) );
  NAND2_X1 U730 ( .A1(n663), .A2(G900), .ZN(n664) );
  NAND2_X1 U731 ( .A1(n664), .A2(G953), .ZN(n665) );
  NAND2_X1 U732 ( .A1(n666), .A2(n665), .ZN(G72) );
  XNOR2_X1 U733 ( .A(n668), .B(n667), .ZN(n669) );
  NOR2_X1 U734 ( .A1(n669), .A2(n680), .ZN(G66) );
  XOR2_X1 U735 ( .A(KEYINPUT123), .B(n671), .Z(n672) );
  XNOR2_X1 U736 ( .A(n673), .B(n672), .ZN(n674) );
  NOR2_X1 U737 ( .A1(n674), .A2(n680), .ZN(G63) );
  NAND2_X1 U738 ( .A1(n351), .A2(G469), .ZN(n679) );
  XOR2_X1 U739 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n676) );
  XNOR2_X1 U740 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U741 ( .A(n679), .B(n678), .ZN(n681) );
  NOR2_X1 U742 ( .A1(n681), .A2(n680), .ZN(G54) );
  AND2_X1 U743 ( .A1(n683), .A2(n682), .ZN(n720) );
  XOR2_X1 U744 ( .A(KEYINPUT51), .B(KEYINPUT118), .Z(n695) );
  NOR2_X1 U745 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U746 ( .A(n686), .B(KEYINPUT50), .ZN(n687) );
  NOR2_X1 U747 ( .A1(n688), .A2(n687), .ZN(n692) );
  NOR2_X1 U748 ( .A1(n428), .A2(n689), .ZN(n690) );
  XNOR2_X1 U749 ( .A(n690), .B(KEYINPUT49), .ZN(n691) );
  NAND2_X1 U750 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U751 ( .A(n695), .B(n694), .ZN(n696) );
  NAND2_X1 U752 ( .A1(n713), .A2(n696), .ZN(n707) );
  INV_X1 U753 ( .A(n697), .ZN(n712) );
  NAND2_X1 U754 ( .A1(n699), .A2(n698), .ZN(n701) );
  NAND2_X1 U755 ( .A1(n701), .A2(n700), .ZN(n704) );
  NAND2_X1 U756 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U757 ( .A1(n712), .A2(n705), .ZN(n706) );
  NAND2_X1 U758 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U759 ( .A(KEYINPUT52), .B(n708), .Z(n709) );
  NOR2_X1 U760 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U761 ( .A(KEYINPUT119), .B(n711), .Z(n715) );
  AND2_X1 U762 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U763 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U764 ( .A(n716), .B(KEYINPUT120), .ZN(n718) );
  INV_X1 U765 ( .A(G953), .ZN(n717) );
  NAND2_X1 U766 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U767 ( .A1(n720), .A2(n719), .ZN(n722) );
  XOR2_X1 U768 ( .A(KEYINPUT121), .B(KEYINPUT53), .Z(n721) );
  XNOR2_X1 U769 ( .A(n722), .B(n721), .ZN(G75) );
  INV_X1 U770 ( .A(n732), .ZN(n736) );
  NOR2_X1 U771 ( .A1(n736), .A2(n725), .ZN(n724) );
  XNOR2_X1 U772 ( .A(G104), .B(KEYINPUT115), .ZN(n723) );
  XNOR2_X1 U773 ( .A(n724), .B(n723), .ZN(G6) );
  NOR2_X1 U774 ( .A1(n739), .A2(n725), .ZN(n727) );
  XNOR2_X1 U775 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n726) );
  XNOR2_X1 U776 ( .A(n727), .B(n726), .ZN(n728) );
  XNOR2_X1 U777 ( .A(G107), .B(n728), .ZN(G9) );
  XOR2_X1 U778 ( .A(G128), .B(KEYINPUT29), .Z(n731) );
  NAND2_X1 U779 ( .A1(n733), .A2(n729), .ZN(n730) );
  XNOR2_X1 U780 ( .A(n731), .B(n730), .ZN(G30) );
  XOR2_X1 U781 ( .A(G146), .B(KEYINPUT117), .Z(n735) );
  NAND2_X1 U782 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U783 ( .A(n735), .B(n734), .ZN(G48) );
  NOR2_X1 U784 ( .A1(n736), .A2(n738), .ZN(n737) );
  XOR2_X1 U785 ( .A(G113), .B(n737), .Z(G15) );
  NOR2_X1 U786 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U787 ( .A(G116), .B(n740), .Z(G18) );
  XNOR2_X1 U788 ( .A(G125), .B(n741), .ZN(n742) );
  XNOR2_X1 U789 ( .A(n742), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U790 ( .A(G134), .B(n743), .Z(G36) );
  XNOR2_X1 U791 ( .A(G101), .B(KEYINPUT125), .ZN(n744) );
  XNOR2_X1 U792 ( .A(n745), .B(n744), .ZN(n747) );
  NAND2_X1 U793 ( .A1(n747), .A2(n746), .ZN(n755) );
  NOR2_X1 U794 ( .A1(n748), .A2(G953), .ZN(n749) );
  XOR2_X1 U795 ( .A(n749), .B(KEYINPUT124), .Z(n753) );
  NAND2_X1 U796 ( .A1(G953), .A2(G224), .ZN(n750) );
  XNOR2_X1 U797 ( .A(KEYINPUT61), .B(n750), .ZN(n751) );
  NAND2_X1 U798 ( .A1(n751), .A2(G898), .ZN(n752) );
  NAND2_X1 U799 ( .A1(n753), .A2(n752), .ZN(n754) );
  XOR2_X1 U800 ( .A(n755), .B(n754), .Z(n756) );
  XNOR2_X1 U801 ( .A(KEYINPUT126), .B(n756), .ZN(G69) );
  XNOR2_X1 U802 ( .A(n757), .B(G131), .ZN(G33) );
endmodule

