//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1 1 1 0 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n566, new_n567,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n631, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1271;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT65), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n453), .A2(new_n457), .B1(new_n448), .B2(new_n454), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT66), .Z(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G137), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AND3_X1   g041(.A1(new_n460), .A2(G101), .A3(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT67), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n463), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n471));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n470), .B(new_n471), .C1(new_n474), .C2(new_n461), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n468), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n477), .B1(new_n464), .B2(new_n465), .ZN(new_n478));
  AND2_X1   g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  OAI21_X1  g054(.A(G2105), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n484));
  OR2_X1    g059(.A1(new_n484), .A2(KEYINPUT69), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(KEYINPUT69), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n460), .B1(new_n464), .B2(new_n465), .ZN(new_n487));
  AOI22_X1  g062(.A1(new_n485), .A2(new_n486), .B1(G124), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(KEYINPUT68), .B1(new_n474), .B2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n464), .A2(new_n465), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n490), .A2(new_n491), .A3(new_n460), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G136), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n488), .A2(new_n494), .ZN(G162));
  OAI211_X1 g070(.A(G126), .B(G2105), .C1(new_n472), .C2(new_n473), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n502), .B1(new_n472), .B2(new_n473), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT4), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n490), .A2(new_n505), .A3(new_n502), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n500), .B1(new_n504), .B2(new_n506), .ZN(G164));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT70), .B1(new_n508), .B2(G651), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT6), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n513), .B1(new_n511), .B2(KEYINPUT6), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n508), .A2(KEYINPUT71), .A3(G651), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n509), .A2(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n516), .A2(G50), .A3(G543), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n522), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n509), .A2(new_n512), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n514), .A2(new_n515), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n525), .A2(new_n526), .A3(new_n522), .ZN(new_n527));
  OAI221_X1 g102(.A(new_n517), .B1(new_n523), .B2(new_n511), .C1(new_n524), .C2(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  XNOR2_X1  g104(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n530), .B(new_n531), .ZN(new_n532));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n532), .B1(new_n522), .B2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n527), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G89), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n525), .A2(new_n526), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n519), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G51), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n534), .A2(new_n536), .A3(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  NAND2_X1  g116(.A1(new_n538), .A2(G52), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n535), .A2(G90), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n522), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(new_n511), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n542), .A2(new_n543), .A3(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  NAND4_X1  g122(.A1(new_n525), .A2(new_n526), .A3(G43), .A4(G543), .ZN(new_n548));
  NAND4_X1  g123(.A1(new_n525), .A2(new_n526), .A3(G81), .A4(new_n522), .ZN(new_n549));
  AND2_X1   g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT73), .ZN(new_n551));
  INV_X1    g126(.A(G56), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n552), .B1(new_n520), .B2(new_n521), .ZN(new_n553));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n551), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  AND2_X1   g131(.A1(KEYINPUT5), .A2(G543), .ZN(new_n557));
  NOR2_X1   g132(.A1(KEYINPUT5), .A2(G543), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g134(.A(KEYINPUT73), .B(new_n554), .C1(new_n559), .C2(new_n552), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n556), .A2(new_n560), .A3(G651), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n550), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  NAND2_X1  g143(.A1(new_n527), .A2(KEYINPUT74), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT74), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n525), .A2(new_n526), .A3(new_n570), .A4(new_n522), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(G91), .A3(new_n571), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n525), .A2(new_n526), .A3(G53), .A4(G543), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(KEYINPUT9), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n516), .A2(new_n575), .A3(G53), .A4(G543), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(G65), .ZN(new_n578));
  OAI21_X1  g153(.A(KEYINPUT75), .B1(new_n557), .B2(new_n558), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT75), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n520), .A2(new_n580), .A3(new_n521), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n578), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  AND2_X1   g157(.A1(G78), .A2(G543), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n572), .A2(new_n577), .A3(new_n584), .ZN(G299));
  OR2_X1    g160(.A1(new_n522), .A2(G74), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n538), .A2(G49), .B1(G651), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n569), .A2(G87), .A3(new_n571), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(G288));
  NAND3_X1  g164(.A1(new_n569), .A2(G86), .A3(new_n571), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n525), .A2(new_n526), .A3(G48), .A4(G543), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n520), .B2(new_n521), .ZN(new_n593));
  AND2_X1   g168(.A1(G73), .A2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n590), .A2(new_n597), .ZN(G305));
  AOI22_X1  g173(.A1(new_n522), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n599), .A2(new_n511), .ZN(new_n600));
  XOR2_X1   g175(.A(KEYINPUT76), .B(G47), .Z(new_n601));
  NAND4_X1  g176(.A1(new_n525), .A2(new_n601), .A3(new_n526), .A4(G543), .ZN(new_n602));
  INV_X1    g177(.A(G85), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n527), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n604), .A2(KEYINPUT77), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT77), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n516), .A2(G85), .A3(new_n522), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(new_n602), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n600), .B1(new_n605), .B2(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n569), .A2(G92), .A3(new_n571), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g188(.A1(new_n569), .A2(KEYINPUT10), .A3(G92), .A4(new_n571), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AND3_X1   g190(.A1(new_n516), .A2(G54), .A3(G543), .ZN(new_n616));
  AND2_X1   g191(.A1(G79), .A2(G543), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n579), .A2(new_n581), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G66), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT78), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n511), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(G66), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n622), .B1(new_n579), .B2(new_n581), .ZN(new_n623));
  OAI21_X1  g198(.A(KEYINPUT78), .B1(new_n623), .B2(new_n617), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n616), .B1(new_n621), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n615), .A2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n610), .B1(new_n627), .B2(G868), .ZN(G284));
  OAI21_X1  g203(.A(new_n610), .B1(new_n627), .B2(G868), .ZN(G321));
  INV_X1    g204(.A(G868), .ZN(new_n630));
  NAND2_X1  g205(.A1(G299), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(G168), .B2(new_n630), .ZN(G297));
  OAI21_X1  g207(.A(new_n631), .B1(G168), .B2(new_n630), .ZN(G280));
  INV_X1    g208(.A(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n627), .B1(new_n634), .B2(G860), .ZN(G148));
  OAI21_X1  g210(.A(KEYINPUT79), .B1(new_n626), .B2(G559), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT79), .ZN(new_n637));
  NAND4_X1  g212(.A1(new_n615), .A2(new_n625), .A3(new_n637), .A4(new_n634), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n636), .A2(G868), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n563), .A2(new_n630), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(KEYINPUT80), .B(KEYINPUT11), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(G282));
  INV_X1    g218(.A(new_n641), .ZN(G323));
  NAND2_X1  g219(.A1(new_n490), .A2(new_n469), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT12), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT13), .ZN(new_n647));
  INV_X1    g222(.A(G2100), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n493), .A2(G135), .ZN(new_n650));
  INV_X1    g225(.A(G2096), .ZN(new_n651));
  OAI21_X1  g226(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n652));
  INV_X1    g227(.A(G111), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n652), .B1(new_n653), .B2(G2105), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n654), .B1(G123), .B2(new_n487), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n650), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n647), .A2(new_n648), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n650), .A2(new_n655), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(G2096), .ZN(new_n659));
  NAND4_X1  g234(.A1(new_n649), .A2(new_n656), .A3(new_n657), .A4(new_n659), .ZN(G156));
  XNOR2_X1  g235(.A(KEYINPUT15), .B(G2435), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT83), .B(G2438), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2427), .B(G2430), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n665), .A2(KEYINPUT14), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT84), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G1341), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(G1348), .ZN(new_n670));
  XOR2_X1   g245(.A(G2443), .B(G2446), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT82), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G2451), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(G2454), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n673), .B(new_n675), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n668), .A2(G1341), .ZN(new_n677));
  INV_X1    g252(.A(G1348), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n668), .A2(G1341), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n670), .A2(new_n676), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G14), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n676), .B1(new_n670), .B2(new_n680), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT85), .Z(G401));
  INV_X1    g260(.A(KEYINPUT18), .ZN(new_n686));
  XOR2_X1   g261(.A(G2084), .B(G2090), .Z(new_n687));
  XNOR2_X1  g262(.A(G2067), .B(G2678), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(KEYINPUT17), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n687), .A2(new_n688), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n686), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(new_n648), .ZN(new_n693));
  XOR2_X1   g268(.A(G2072), .B(G2078), .Z(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n689), .B2(KEYINPUT18), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(new_n651), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n693), .B(new_n696), .ZN(G227));
  XNOR2_X1  g272(.A(G1971), .B(G1976), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT19), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(G1956), .B(G2474), .Z(new_n701));
  XOR2_X1   g276(.A(G1961), .B(G1966), .Z(new_n702));
  AND2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT20), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n701), .A2(new_n702), .ZN(new_n706));
  NOR3_X1   g281(.A1(new_n700), .A2(new_n703), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(new_n700), .B2(new_n706), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(G1991), .B(G1996), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT86), .Z(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n709), .A2(new_n710), .ZN(new_n715));
  INV_X1    g290(.A(new_n713), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n709), .A2(new_n710), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(G1981), .B(G1986), .ZN(new_n719));
  AND3_X1   g294(.A1(new_n714), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n719), .B1(new_n714), .B2(new_n718), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(G229));
  NAND2_X1  g298(.A1(G162), .A2(G29), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G29), .B2(G35), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n725), .A2(new_n727), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G2090), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(KEYINPUT99), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G29), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G26), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT28), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n489), .A2(G140), .A3(new_n492), .ZN(new_n738));
  OAI21_X1  g313(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n739));
  INV_X1    g314(.A(G116), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n739), .B1(new_n740), .B2(G2105), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G128), .B2(new_n487), .ZN(new_n742));
  AND3_X1   g317(.A1(new_n738), .A2(KEYINPUT92), .A3(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(KEYINPUT92), .B1(new_n738), .B2(new_n742), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n737), .B1(new_n745), .B2(new_n735), .ZN(new_n746));
  INV_X1    g321(.A(G2067), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n732), .B2(KEYINPUT99), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n735), .A2(G32), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n490), .A2(G129), .A3(G2105), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(KEYINPUT94), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT94), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n487), .A2(new_n753), .A3(G129), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n489), .A2(G141), .A3(new_n492), .ZN(new_n756));
  NAND3_X1  g331(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT26), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g334(.A1(KEYINPUT26), .A2(G117), .A3(G2104), .A4(G2105), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n469), .A2(G105), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  AND4_X1   g339(.A1(KEYINPUT95), .A2(new_n755), .A3(new_n756), .A4(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n763), .B1(new_n752), .B2(new_n754), .ZN(new_n766));
  AOI21_X1  g341(.A(KEYINPUT95), .B1(new_n766), .B2(new_n756), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n750), .B1(new_n768), .B2(new_n735), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT27), .B(G1996), .Z(new_n770));
  NOR2_X1   g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR3_X1   g346(.A1(new_n734), .A2(new_n749), .A3(new_n771), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT25), .Z(new_n774));
  AOI22_X1  g349(.A1(new_n490), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(new_n460), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G139), .B2(new_n493), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n777), .A2(new_n735), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n735), .B2(G33), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT93), .Z(new_n780));
  NAND2_X1  g355(.A1(new_n780), .A2(G2072), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n779), .B(KEYINPUT93), .ZN(new_n782));
  INV_X1    g357(.A(G2072), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(G16), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(G19), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n563), .B2(new_n785), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT90), .B(G1341), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT91), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n787), .B(new_n789), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n781), .A2(new_n784), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n730), .A2(new_n731), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n785), .A2(G21), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G168), .B2(new_n785), .ZN(new_n794));
  INV_X1    g369(.A(G1966), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n735), .B1(KEYINPUT24), .B2(G34), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(KEYINPUT24), .B2(G34), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(new_n481), .B2(G29), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G2084), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT31), .B(G11), .Z(new_n802));
  INV_X1    g377(.A(G28), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n803), .A2(KEYINPUT30), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT96), .ZN(new_n805));
  AOI21_X1  g380(.A(G29), .B1(new_n803), .B2(KEYINPUT30), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n802), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n658), .B2(new_n735), .ZN(new_n808));
  NOR2_X1   g383(.A1(G27), .A2(G29), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G164), .B2(G29), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n810), .A2(G2078), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n810), .A2(G2078), .ZN(new_n812));
  NOR3_X1   g387(.A1(new_n808), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n785), .A2(G5), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(G171), .B2(new_n785), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n801), .B(new_n813), .C1(G1961), .C2(new_n815), .ZN(new_n816));
  NOR3_X1   g391(.A1(new_n791), .A2(new_n797), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n769), .A2(new_n770), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n785), .A2(G20), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT23), .ZN(new_n820));
  AND3_X1   g395(.A1(new_n572), .A2(new_n577), .A3(new_n584), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n821), .B2(new_n785), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n818), .B1(G1956), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n815), .A2(G1961), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT97), .Z(new_n825));
  AOI211_X1 g400(.A(new_n823), .B(new_n825), .C1(G1956), .C2(new_n822), .ZN(new_n826));
  NOR2_X1   g401(.A1(G4), .A2(G16), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT89), .Z(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n626), .B2(new_n785), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(G1348), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n772), .A2(new_n817), .A3(new_n826), .A4(new_n830), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n785), .A2(G22), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(G303), .B2(G16), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(G1971), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT32), .B(G1981), .Z(new_n835));
  AND2_X1   g410(.A1(new_n785), .A2(G6), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(G305), .B2(G16), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n834), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(G16), .A2(G23), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT87), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(G288), .B2(new_n785), .ZN(new_n841));
  XNOR2_X1  g416(.A(KEYINPUT33), .B(G1976), .ZN(new_n842));
  AOI22_X1  g417(.A1(new_n841), .A2(new_n842), .B1(new_n837), .B2(new_n835), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n842), .B2(new_n841), .ZN(new_n844));
  OR3_X1    g419(.A1(new_n838), .A2(new_n844), .A3(KEYINPUT34), .ZN(new_n845));
  MUX2_X1   g420(.A(G24), .B(G290), .S(G16), .Z(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(G1986), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n735), .A2(G25), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n493), .A2(G131), .ZN(new_n849));
  OAI21_X1  g424(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n850));
  INV_X1    g425(.A(G107), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n850), .B1(new_n851), .B2(G2105), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n852), .B1(G119), .B2(new_n487), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n848), .B1(new_n855), .B2(new_n735), .ZN(new_n856));
  XOR2_X1   g431(.A(KEYINPUT35), .B(G1991), .Z(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n856), .B(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n847), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n845), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT88), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n845), .A2(new_n860), .A3(KEYINPUT88), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(KEYINPUT34), .B1(new_n838), .B2(new_n844), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(KEYINPUT36), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT36), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n865), .A2(new_n869), .A3(new_n866), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n831), .B1(new_n868), .B2(new_n870), .ZN(G311));
  AND4_X1   g446(.A1(new_n826), .A2(new_n772), .A3(new_n817), .A4(new_n830), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n869), .B1(new_n865), .B2(new_n866), .ZN(new_n873));
  AND3_X1   g448(.A1(new_n865), .A2(new_n869), .A3(new_n866), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(G150));
  NAND4_X1  g450(.A1(new_n525), .A2(new_n526), .A3(G55), .A4(G543), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n525), .A2(new_n526), .A3(G93), .A4(new_n522), .ZN(new_n877));
  INV_X1    g452(.A(G67), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n878), .B1(new_n520), .B2(new_n521), .ZN(new_n879));
  AND2_X1   g454(.A1(G80), .A2(G543), .ZN(new_n880));
  OAI21_X1  g455(.A(G651), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n876), .A2(new_n877), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(G860), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(KEYINPUT37), .Z(new_n884));
  NOR2_X1   g459(.A1(new_n626), .A2(new_n634), .ZN(new_n885));
  XNOR2_X1  g460(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n556), .A2(new_n560), .A3(G651), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n548), .A2(new_n549), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n882), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n876), .A2(new_n877), .A3(new_n881), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n891), .A2(new_n561), .A3(new_n550), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n887), .B(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(KEYINPUT39), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT101), .ZN(new_n896));
  INV_X1    g471(.A(G860), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(new_n894), .B2(KEYINPUT39), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n884), .B1(new_n896), .B2(new_n898), .ZN(G145));
  XNOR2_X1  g474(.A(KEYINPUT105), .B(G37), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(G162), .B(G160), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(new_n658), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n777), .ZN(new_n905));
  OAI21_X1  g480(.A(G164), .B1(new_n743), .B2(new_n744), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n738), .A2(new_n742), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT92), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n504), .A2(new_n506), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n496), .A2(new_n499), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n738), .A2(KEYINPUT92), .A3(new_n742), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n909), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n755), .A2(new_n756), .A3(new_n764), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n906), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n915), .B1(new_n906), .B2(new_n914), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n905), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT103), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI211_X1 g495(.A(KEYINPUT103), .B(new_n905), .C1(new_n916), .C2(new_n917), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n743), .A2(new_n744), .A3(G164), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n912), .B1(new_n909), .B2(new_n913), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n768), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n906), .B(new_n914), .C1(new_n767), .C2(new_n765), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n925), .A2(new_n777), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT102), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n906), .A2(new_n914), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n905), .B1(new_n930), .B2(new_n768), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n931), .A2(KEYINPUT102), .A3(new_n926), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n493), .A2(G142), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n934), .B(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n937));
  INV_X1    g512(.A(G118), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n937), .B1(new_n938), .B2(G2105), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n939), .B1(G130), .B2(new_n487), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n936), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n854), .B(new_n646), .ZN(new_n942));
  XOR2_X1   g517(.A(new_n941), .B(new_n942), .Z(new_n943));
  AND3_X1   g518(.A1(new_n922), .A2(new_n933), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n943), .B1(new_n922), .B2(new_n933), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n904), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n915), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n930), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n906), .A2(new_n914), .A3(new_n915), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT103), .B1(new_n950), .B2(new_n905), .ZN(new_n951));
  INV_X1    g526(.A(new_n921), .ZN(new_n952));
  AND4_X1   g527(.A1(KEYINPUT102), .A2(new_n925), .A3(new_n777), .A4(new_n926), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT102), .B1(new_n931), .B2(new_n926), .ZN(new_n954));
  OAI22_X1  g529(.A1(new_n951), .A2(new_n952), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n943), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n922), .A2(new_n933), .A3(new_n943), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n957), .A2(new_n903), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n901), .B1(new_n946), .B2(new_n959), .ZN(new_n960));
  XOR2_X1   g535(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n961));
  XNOR2_X1  g536(.A(new_n960), .B(new_n961), .ZN(G395));
  NAND2_X1  g537(.A1(new_n636), .A2(new_n638), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n893), .ZN(new_n964));
  INV_X1    g539(.A(new_n893), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n636), .A2(new_n638), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n572), .A2(new_n584), .ZN(new_n968));
  AOI22_X1  g543(.A1(new_n615), .A2(new_n625), .B1(new_n968), .B2(new_n577), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n615), .A2(new_n821), .A3(new_n625), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n967), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n966), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n965), .B1(new_n636), .B2(new_n638), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT41), .B1(new_n970), .B2(new_n969), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n626), .A2(G299), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT41), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n615), .A2(new_n821), .A3(new_n625), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT107), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n975), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n970), .A2(new_n969), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n982), .A2(KEYINPUT107), .A3(new_n977), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n974), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT42), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n971), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n986), .B1(new_n971), .B2(new_n985), .ZN(new_n989));
  INV_X1    g564(.A(G305), .ZN(new_n990));
  NAND2_X1  g565(.A1(G290), .A2(new_n990), .ZN(new_n991));
  OAI211_X1 g566(.A(G305), .B(new_n600), .C1(new_n605), .C2(new_n608), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G288), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(G303), .ZN(new_n995));
  NAND2_X1  g570(.A1(G166), .A2(G288), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n993), .A2(new_n997), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n991), .A2(new_n995), .A3(new_n996), .A4(new_n992), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(KEYINPUT108), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n988), .A2(new_n989), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n971), .A2(new_n985), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT42), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1001), .B1(new_n1005), .B2(new_n987), .ZN(new_n1006));
  OAI21_X1  g581(.A(G868), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n882), .A2(new_n630), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(G295));
  NAND2_X1  g584(.A1(new_n1007), .A2(new_n1008), .ZN(G331));
  AND3_X1   g585(.A1(new_n890), .A2(new_n892), .A3(G301), .ZN(new_n1011));
  AOI21_X1  g586(.A(G301), .B1(new_n890), .B2(new_n892), .ZN(new_n1012));
  OAI21_X1  g587(.A(G286), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n893), .A2(G171), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n890), .A2(new_n892), .A3(G301), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1014), .A2(G168), .A3(new_n1015), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n981), .A2(new_n983), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1019));
  AOI22_X1  g594(.A1(new_n1019), .A2(new_n982), .B1(new_n998), .B2(new_n999), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT110), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1018), .A2(KEYINPUT110), .A3(new_n1020), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1019), .A2(new_n982), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1018), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT109), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1000), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n998), .A2(new_n999), .A3(KEYINPUT109), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(G37), .B1(new_n1027), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT43), .B1(new_n1025), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n975), .A2(new_n979), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n1017), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n1026), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n901), .B1(new_n1036), .B2(new_n1031), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1018), .A2(KEYINPUT110), .A3(new_n1020), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT110), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1037), .B(KEYINPUT43), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT44), .B1(new_n1033), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT44), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT43), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1044), .B1(new_n1025), .B2(new_n1032), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1037), .B(new_n1044), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1043), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1042), .A2(new_n1048), .ZN(G397));
  INV_X1    g624(.A(KEYINPUT45), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1050), .B1(G164), .B2(G1384), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n468), .A2(new_n480), .A3(G40), .A4(new_n475), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n1051), .A2(G1996), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n768), .A2(new_n1053), .ZN(new_n1054));
  XOR2_X1   g629(.A(new_n1054), .B(KEYINPUT111), .Z(new_n1055));
  XNOR2_X1  g630(.A(new_n745), .B(G2067), .ZN(new_n1056));
  INV_X1    g631(.A(G1996), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1056), .B1(new_n1057), .B2(new_n947), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n855), .A2(new_n857), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n854), .A2(new_n858), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1059), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1055), .A2(new_n1060), .A3(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g639(.A(G290), .B(G1986), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1064), .B1(new_n1059), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G1981), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n590), .A2(new_n597), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G86), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n527), .A2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(G1981), .B1(new_n596), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1068), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT49), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1068), .A2(KEYINPUT49), .A3(new_n1071), .ZN(new_n1075));
  INV_X1    g650(.A(G8), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1052), .ZN(new_n1077));
  AOI21_X1  g652(.A(G1384), .B1(new_n910), .B2(new_n911), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1074), .A2(new_n1075), .A3(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n587), .A2(G1976), .A3(new_n588), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT52), .ZN(new_n1083));
  INV_X1    g658(.A(G1976), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT52), .B1(G288), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1085), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1080), .A2(new_n1083), .A3(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT50), .ZN(new_n1089));
  INV_X1    g664(.A(G1384), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n912), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  XOR2_X1   g666(.A(KEYINPUT116), .B(G2084), .Z(new_n1092));
  NAND4_X1  g667(.A1(new_n1088), .A2(new_n1091), .A3(new_n1077), .A4(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1050), .A2(G1384), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1096), .B1(new_n910), .B2(new_n911), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1097), .A2(new_n1052), .ZN(new_n1098));
  AOI21_X1  g673(.A(G1966), .B1(new_n1098), .B2(new_n1051), .ZN(new_n1099));
  OAI211_X1 g674(.A(G8), .B(G168), .C1(new_n1094), .C2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(KEYINPUT117), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n480), .A2(G40), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n476), .B(new_n1102), .C1(G164), .C2(new_n1096), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1078), .A2(KEYINPUT45), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n795), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n1093), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT117), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1106), .A2(new_n1107), .A3(G8), .A4(G168), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1101), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1052), .B1(new_n1097), .B2(KEYINPUT112), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT112), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(G164), .B2(new_n1096), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1114), .A2(new_n1051), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(G1971), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n912), .A2(new_n1090), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1052), .B1(new_n1120), .B2(KEYINPUT50), .ZN(new_n1121));
  AOI211_X1 g696(.A(KEYINPUT50), .B(G1384), .C1(new_n910), .C2(new_n911), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT115), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT115), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1091), .A2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1121), .A2(new_n1123), .A3(new_n1125), .A4(new_n731), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1119), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1113), .B1(new_n1127), .B2(new_n1076), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT63), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1109), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1088), .A2(new_n1077), .A3(new_n1091), .ZN(new_n1131));
  OAI21_X1  g706(.A(KEYINPUT113), .B1(new_n1131), .B2(G2090), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT113), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1121), .A2(new_n1133), .A3(new_n731), .A4(new_n1091), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1119), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT114), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1112), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1138), .A2(KEYINPUT114), .A3(new_n1110), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1135), .A2(G8), .A3(new_n1137), .A4(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1087), .B1(new_n1130), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1079), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1080), .A2(new_n1084), .A3(new_n994), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1142), .B1(new_n1143), .B2(new_n1068), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1087), .B1(new_n1108), .B2(new_n1101), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1135), .A2(G8), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n1113), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1129), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  NOR3_X1   g723(.A1(new_n1141), .A2(new_n1144), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT120), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT119), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1151), .B1(new_n1094), .B2(new_n1099), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1105), .A2(KEYINPUT119), .A3(new_n1093), .ZN(new_n1153));
  AOI21_X1  g728(.A(G286), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT51), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1155), .A2(new_n1076), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1150), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1105), .A2(KEYINPUT119), .A3(new_n1093), .ZN(new_n1159));
  AOI21_X1  g734(.A(KEYINPUT119), .B1(new_n1105), .B2(new_n1093), .ZN(new_n1160));
  OAI21_X1  g735(.A(G168), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1161), .A2(KEYINPUT120), .A3(new_n1156), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1106), .A2(G8), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1163), .B(new_n1155), .C1(new_n1076), .C2(G168), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1158), .A2(new_n1162), .A3(new_n1164), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1152), .A2(G8), .A3(G286), .A4(new_n1153), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT53), .ZN(new_n1168));
  OR4_X1    g743(.A1(new_n1168), .A2(new_n1103), .A3(new_n1104), .A4(G2078), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT118), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1131), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(G1961), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1088), .A2(new_n1091), .A3(KEYINPUT118), .A4(new_n1077), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1168), .B1(new_n1117), .B2(G2078), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1169), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  OR2_X1    g751(.A1(new_n1176), .A2(G171), .ZN(new_n1177));
  XOR2_X1   g752(.A(KEYINPUT121), .B(G2078), .Z(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(KEYINPUT53), .ZN(new_n1179));
  OR2_X1    g754(.A1(new_n1117), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1174), .A2(new_n1180), .A3(new_n1175), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(KEYINPUT122), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(G171), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1181), .A2(KEYINPUT122), .ZN(new_n1184));
  OAI211_X1 g759(.A(KEYINPUT54), .B(new_n1177), .C1(new_n1183), .C2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1176), .A2(G171), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1174), .A2(new_n1180), .A3(G301), .A4(new_n1175), .ZN(new_n1187));
  AOI21_X1  g762(.A(KEYINPUT54), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1087), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1128), .A2(new_n1140), .A3(new_n1189), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1167), .A2(new_n1185), .A3(new_n1191), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1121), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1193));
  INV_X1    g768(.A(G1956), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT57), .ZN(new_n1196));
  XNOR2_X1  g771(.A(G299), .B(new_n1196), .ZN(new_n1197));
  XNOR2_X1  g772(.A(KEYINPUT56), .B(G2072), .ZN(new_n1198));
  NAND4_X1  g773(.A1(new_n1114), .A2(new_n1051), .A3(new_n1116), .A4(new_n1198), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1195), .A2(new_n1197), .A3(new_n1199), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1171), .A2(new_n678), .A3(new_n1173), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1077), .A2(new_n747), .A3(new_n1078), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1200), .A2(new_n1203), .A3(new_n627), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1195), .A2(new_n1199), .ZN(new_n1205));
  INV_X1    g780(.A(new_n1197), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1204), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g783(.A(KEYINPUT61), .ZN(new_n1209));
  AND3_X1   g784(.A1(new_n1195), .A2(new_n1197), .A3(new_n1199), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1197), .B1(new_n1195), .B2(new_n1199), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1209), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1207), .A2(KEYINPUT61), .A3(new_n1200), .ZN(new_n1213));
  NAND4_X1  g788(.A1(new_n1114), .A2(new_n1057), .A3(new_n1051), .A4(new_n1116), .ZN(new_n1214));
  XOR2_X1   g789(.A(KEYINPUT58), .B(G1341), .Z(new_n1215));
  OAI21_X1  g790(.A(new_n1215), .B1(new_n1120), .B2(new_n1052), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n562), .B1(new_n1214), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g792(.A(KEYINPUT59), .ZN(new_n1218));
  XNOR2_X1  g793(.A(new_n1217), .B(new_n1218), .ZN(new_n1219));
  AND3_X1   g794(.A1(new_n1212), .A2(new_n1213), .A3(new_n1219), .ZN(new_n1220));
  NAND3_X1  g795(.A1(new_n1201), .A2(KEYINPUT60), .A3(new_n1202), .ZN(new_n1221));
  XNOR2_X1  g796(.A(new_n1221), .B(new_n627), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT60), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1203), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g800(.A(new_n1208), .B1(new_n1220), .B2(new_n1225), .ZN(new_n1226));
  OAI21_X1  g801(.A(new_n1149), .B1(new_n1192), .B2(new_n1226), .ZN(new_n1227));
  INV_X1    g802(.A(KEYINPUT62), .ZN(new_n1228));
  AND3_X1   g803(.A1(new_n1165), .A2(new_n1228), .A3(new_n1166), .ZN(new_n1229));
  AOI21_X1  g804(.A(new_n1228), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1230));
  OR2_X1    g805(.A1(new_n1190), .A2(new_n1186), .ZN(new_n1231));
  NOR3_X1   g806(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  OAI21_X1  g807(.A(new_n1066), .B1(new_n1227), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g808(.A1(new_n745), .A2(new_n747), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1055), .A2(new_n1060), .ZN(new_n1235));
  XNOR2_X1  g810(.A(new_n1062), .B(KEYINPUT123), .ZN(new_n1236));
  OAI21_X1  g811(.A(new_n1234), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g812(.A1(new_n1237), .A2(new_n1059), .ZN(new_n1238));
  INV_X1    g813(.A(KEYINPUT127), .ZN(new_n1239));
  NAND2_X1  g814(.A1(new_n1064), .A2(new_n1239), .ZN(new_n1240));
  NOR4_X1   g815(.A1(G290), .A2(G1986), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1241));
  XOR2_X1   g816(.A(new_n1241), .B(KEYINPUT48), .Z(new_n1242));
  NAND2_X1  g817(.A1(new_n1240), .A2(new_n1242), .ZN(new_n1243));
  NOR2_X1   g818(.A1(new_n1064), .A2(new_n1239), .ZN(new_n1244));
  OAI21_X1  g819(.A(new_n1238), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g820(.A(KEYINPUT124), .ZN(new_n1246));
  INV_X1    g821(.A(KEYINPUT46), .ZN(new_n1247));
  OR3_X1    g822(.A1(new_n1053), .A2(new_n1246), .A3(new_n1247), .ZN(new_n1248));
  OAI21_X1  g823(.A(new_n1053), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1249));
  AOI22_X1  g824(.A1(new_n1248), .A2(new_n1249), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1250));
  NAND2_X1  g825(.A1(new_n1056), .A2(new_n947), .ZN(new_n1251));
  AND3_X1   g826(.A1(new_n1251), .A2(KEYINPUT125), .A3(new_n1059), .ZN(new_n1252));
  AOI21_X1  g827(.A(KEYINPUT125), .B1(new_n1251), .B2(new_n1059), .ZN(new_n1253));
  OAI21_X1  g828(.A(new_n1250), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  INV_X1    g829(.A(KEYINPUT126), .ZN(new_n1255));
  OR2_X1    g830(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g831(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1257));
  NAND2_X1  g832(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g833(.A1(new_n1258), .A2(KEYINPUT47), .ZN(new_n1259));
  INV_X1    g834(.A(KEYINPUT47), .ZN(new_n1260));
  NAND3_X1  g835(.A1(new_n1256), .A2(new_n1260), .A3(new_n1257), .ZN(new_n1261));
  AOI21_X1  g836(.A(new_n1245), .B1(new_n1259), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g837(.A1(new_n1233), .A2(new_n1262), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g838(.A(G319), .ZN(new_n1265));
  NOR2_X1   g839(.A1(new_n1265), .A2(G227), .ZN(new_n1266));
  OAI211_X1 g840(.A(new_n722), .B(new_n1266), .C1(new_n682), .C2(new_n683), .ZN(new_n1267));
  OAI21_X1  g841(.A(new_n1032), .B1(new_n1039), .B2(new_n1038), .ZN(new_n1268));
  NAND2_X1  g842(.A1(new_n1268), .A2(KEYINPUT43), .ZN(new_n1269));
  AOI211_X1 g843(.A(new_n1267), .B(new_n960), .C1(new_n1269), .C2(new_n1046), .ZN(G308));
  NOR2_X1   g844(.A1(new_n960), .A2(new_n1267), .ZN(new_n1271));
  OAI21_X1  g845(.A(new_n1271), .B1(new_n1045), .B2(new_n1047), .ZN(G225));
endmodule


