//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 1 0 0 1 1 1 1 1 1 0 0 1 0 1 1 0 1 1 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 0 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032;
  NOR2_X1   g000(.A1(G475), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G140), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G125), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(KEYINPUT16), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G140), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n192), .A3(KEYINPUT16), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT77), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n190), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n189), .A2(new_n192), .A3(KEYINPUT77), .A4(KEYINPUT16), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n195), .A2(G146), .A3(new_n196), .ZN(new_n200));
  NOR2_X1   g014(.A1(G237), .A2(G953), .ZN(new_n201));
  AOI21_X1  g015(.A(G143), .B1(new_n201), .B2(G214), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n201), .A2(G143), .A3(G214), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(KEYINPUT17), .A3(G131), .ZN(new_n206));
  INV_X1    g020(.A(new_n204), .ZN(new_n207));
  OAI21_X1  g021(.A(G131), .B1(new_n207), .B2(new_n202), .ZN(new_n208));
  INV_X1    g022(.A(G131), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n203), .A2(new_n209), .A3(new_n204), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT17), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n208), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n199), .A2(new_n200), .A3(new_n206), .A4(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(G113), .B(G122), .ZN(new_n214));
  INV_X1    g028(.A(G104), .ZN(new_n215));
  XNOR2_X1  g029(.A(new_n214), .B(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n189), .A2(new_n192), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT90), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n189), .A2(new_n192), .A3(KEYINPUT90), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(G146), .A3(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n189), .A2(new_n192), .A3(new_n198), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n205), .A2(KEYINPUT18), .A3(G131), .ZN(new_n224));
  NAND2_X1  g038(.A1(KEYINPUT18), .A2(G131), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n203), .A2(new_n204), .A3(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n223), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n213), .A2(new_n216), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n208), .A2(new_n210), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n219), .A2(KEYINPUT19), .A3(new_n220), .ZN(new_n230));
  OR2_X1    g044(.A1(new_n217), .A2(KEYINPUT19), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n200), .B(new_n229), .C1(new_n232), .C2(G146), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n216), .B1(new_n233), .B2(new_n227), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n187), .B1(new_n228), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT20), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT20), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n237), .B(new_n187), .C1(new_n228), .C2(new_n234), .ZN(new_n238));
  INV_X1    g052(.A(G902), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n216), .B1(new_n213), .B2(new_n227), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n239), .B1(new_n228), .B2(new_n240), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n236), .A2(new_n238), .B1(G475), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G953), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G952), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n244), .B1(G234), .B2(G237), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT21), .B(G898), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(G234), .A2(G237), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(G902), .A3(G953), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n246), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G116), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G122), .ZN(new_n253));
  INV_X1    g067(.A(G122), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G116), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G107), .ZN(new_n257));
  INV_X1    g071(.A(G107), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n253), .A2(new_n255), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT91), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT13), .ZN(new_n263));
  INV_X1    g077(.A(G128), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n263), .B1(new_n264), .B2(G143), .ZN(new_n265));
  INV_X1    g079(.A(G143), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(KEYINPUT13), .A3(G128), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n265), .B(new_n267), .C1(G128), .C2(new_n266), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT66), .B(G134), .ZN(new_n269));
  XNOR2_X1  g083(.A(G128), .B(G143), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n268), .A2(G134), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n257), .A2(KEYINPUT91), .A3(new_n259), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n262), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n253), .A2(KEYINPUT14), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n255), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n253), .A2(KEYINPUT14), .ZN(new_n276));
  OAI21_X1  g090(.A(G107), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n270), .A2(new_n269), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n270), .A2(new_n269), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n277), .B(new_n259), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n273), .A2(new_n280), .ZN(new_n281));
  XOR2_X1   g095(.A(KEYINPUT75), .B(G217), .Z(new_n282));
  XOR2_X1   g096(.A(KEYINPUT9), .B(G234), .Z(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n283), .A3(new_n243), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n284), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n273), .A2(new_n280), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(G902), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G478), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n289), .A2(KEYINPUT15), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT92), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n287), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n286), .B1(new_n273), .B2(new_n280), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n239), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT92), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(new_n296), .A3(new_n290), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n239), .B(new_n291), .C1(new_n293), .C2(new_n294), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT93), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n285), .A2(new_n287), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT93), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n300), .A2(new_n301), .A3(new_n239), .A4(new_n291), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n292), .A2(new_n297), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n242), .A2(new_n251), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT94), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n242), .A2(new_n303), .A3(KEYINPUT94), .A4(new_n251), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(G214), .B1(G237), .B2(G902), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(G210), .B1(G237), .B2(G902), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT6), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT81), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n258), .A2(G104), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT80), .ZN(new_n316));
  OAI22_X1  g130(.A1(new_n316), .A2(KEYINPUT3), .B1(new_n215), .B2(G107), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT80), .B(KEYINPUT3), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n258), .A2(G104), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n315), .B(new_n317), .C1(new_n318), .C2(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n313), .B1(new_n320), .B2(G101), .ZN(new_n321));
  INV_X1    g135(.A(new_n319), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT3), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT80), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n323), .A2(KEYINPUT80), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n322), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n314), .B1(new_n319), .B2(new_n324), .ZN(new_n328));
  INV_X1    g142(.A(G101), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n327), .A2(new_n328), .A3(KEYINPUT81), .A4(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n321), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n329), .B1(new_n327), .B2(new_n328), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT4), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT68), .ZN(new_n336));
  XOR2_X1   g150(.A(KEYINPUT2), .B(G113), .Z(new_n337));
  XNOR2_X1  g151(.A(G116), .B(G119), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G119), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G116), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n252), .A2(G119), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT2), .B(G113), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n344), .A3(KEYINPUT68), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n339), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT69), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n337), .A2(new_n347), .A3(new_n338), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT69), .B1(new_n343), .B2(new_n344), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n346), .A2(new_n350), .B1(new_n332), .B2(new_n333), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT82), .B1(new_n258), .B2(G104), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT82), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(new_n215), .A3(G107), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n352), .A2(new_n354), .A3(new_n319), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G101), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n357), .B1(new_n321), .B2(new_n330), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n338), .A2(KEYINPUT5), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT5), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n360), .A2(new_n340), .A3(G116), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n359), .A2(KEYINPUT86), .A3(G113), .A4(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT86), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n341), .A2(new_n342), .A3(KEYINPUT5), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n361), .A2(G113), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n350), .A2(new_n362), .A3(new_n366), .ZN(new_n367));
  AOI22_X1  g181(.A1(new_n335), .A2(new_n351), .B1(new_n358), .B2(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(G110), .B(G122), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n312), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n369), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n335), .A2(new_n351), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n331), .A2(new_n356), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n350), .A2(new_n362), .A3(new_n366), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n371), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n370), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n198), .A2(G143), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n266), .A2(G146), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(KEYINPUT0), .A2(G128), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT64), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n382), .B1(KEYINPUT0), .B2(G128), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT0), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(new_n264), .A3(KEYINPUT64), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n380), .A2(new_n381), .A3(new_n383), .A4(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(G143), .B(G146), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(KEYINPUT0), .A3(G128), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G125), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT1), .B1(new_n266), .B2(G146), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G128), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n380), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n387), .A2(G128), .A3(new_n391), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(new_n394), .A3(new_n191), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n243), .A2(G224), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n397), .B(KEYINPUT87), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n396), .B(new_n398), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n312), .B(new_n371), .C1(new_n372), .C2(new_n375), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n377), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n395), .A2(KEYINPUT88), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT88), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n393), .A2(new_n394), .A3(new_n403), .A4(new_n191), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n402), .A2(new_n390), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n397), .A2(KEYINPUT7), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n406), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n390), .A2(new_n395), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT89), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n390), .A2(KEYINPUT89), .A3(new_n395), .A4(new_n408), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n407), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n413), .B1(new_n369), .B2(new_n368), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n350), .B1(new_n364), .B2(new_n365), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n358), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n369), .B(KEYINPUT8), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n416), .B(new_n417), .C1(new_n358), .C2(new_n374), .ZN(new_n418));
  AOI21_X1  g232(.A(G902), .B1(new_n414), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n311), .B1(new_n401), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n401), .A2(new_n419), .A3(new_n311), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n310), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n308), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G469), .ZN(new_n425));
  INV_X1    g239(.A(G137), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n426), .A2(KEYINPUT11), .A3(G134), .ZN(new_n427));
  INV_X1    g241(.A(G134), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(KEYINPUT66), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT66), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G134), .ZN(new_n431));
  AOI21_X1  g245(.A(G137), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(KEYINPUT65), .B(KEYINPUT11), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n427), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n429), .A2(new_n431), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n435), .A2(new_n426), .ZN(new_n436));
  OAI21_X1  g250(.A(G131), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(G131), .B1(new_n269), .B2(G137), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n438), .B(new_n427), .C1(new_n432), .C2(new_n433), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT12), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT84), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT1), .ZN(new_n443));
  AND4_X1   g257(.A1(new_n443), .A2(new_n378), .A3(new_n379), .A4(G128), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n391), .A2(G128), .B1(new_n378), .B2(new_n379), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n358), .A2(new_n447), .ZN(new_n448));
  AOI211_X1 g262(.A(new_n357), .B(new_n446), .C1(new_n321), .C2(new_n330), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n440), .B(new_n442), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n440), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n373), .A2(new_n446), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n331), .A2(new_n447), .A3(new_n356), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n450), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n389), .B1(new_n332), .B2(new_n333), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n449), .A2(KEYINPUT10), .B1(new_n335), .B2(new_n457), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n449), .A2(KEYINPUT83), .A3(KEYINPUT10), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT83), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT10), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n460), .B1(new_n453), .B2(new_n461), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n458), .B(new_n451), .C1(new_n459), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n456), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(G110), .B(G140), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n243), .A2(G227), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n465), .B(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n458), .B1(new_n459), .B2(new_n462), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n440), .ZN(new_n470));
  INV_X1    g284(.A(new_n467), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(new_n463), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n425), .B1(new_n473), .B2(new_n239), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n471), .B1(new_n470), .B2(new_n463), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n456), .A2(new_n463), .A3(new_n471), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n425), .B(new_n239), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT85), .ZN(new_n478));
  INV_X1    g292(.A(new_n463), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT83), .B1(new_n449), .B2(KEYINPUT10), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n453), .A2(new_n460), .A3(new_n461), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n451), .B1(new_n482), .B2(new_n458), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n467), .B1(new_n479), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n456), .A2(new_n463), .A3(new_n471), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT85), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n486), .A2(new_n487), .A3(new_n425), .A4(new_n239), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n474), .B1(new_n478), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(G221), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n490), .B1(new_n283), .B2(new_n239), .ZN(new_n491));
  NOR3_X1   g305(.A1(new_n424), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(G472), .A2(G902), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT32), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n201), .A2(G210), .ZN(new_n497));
  XOR2_X1   g311(.A(new_n497), .B(KEYINPUT27), .Z(new_n498));
  XNOR2_X1  g312(.A(KEYINPUT26), .B(G101), .ZN(new_n499));
  XOR2_X1   g313(.A(new_n498), .B(new_n499), .Z(new_n500));
  NOR2_X1   g314(.A1(new_n426), .A2(G134), .ZN(new_n501));
  OAI21_X1  g315(.A(G131), .B1(new_n432), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n209), .B1(new_n435), .B2(new_n426), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n502), .B1(new_n434), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT70), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT70), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n439), .A2(new_n506), .A3(new_n502), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n505), .A2(new_n507), .A3(new_n447), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n346), .A2(new_n350), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n389), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n440), .A2(new_n511), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n508), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT67), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n504), .A2(new_n514), .ZN(new_n515));
  OAI211_X1 g329(.A(KEYINPUT67), .B(new_n502), .C1(new_n434), .C2(new_n503), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n447), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n510), .B1(new_n517), .B2(new_n512), .ZN(new_n518));
  OAI21_X1  g332(.A(KEYINPUT28), .B1(new_n513), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT28), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n508), .A2(new_n510), .A3(new_n512), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n519), .A2(KEYINPUT72), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT72), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n523), .B(KEYINPUT28), .C1(new_n513), .C2(new_n518), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n500), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT73), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n508), .A2(KEYINPUT30), .A3(new_n512), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n446), .B1(new_n504), .B2(new_n514), .ZN(new_n528));
  AOI22_X1  g342(.A1(new_n528), .A2(new_n516), .B1(new_n440), .B2(new_n511), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n527), .B(new_n509), .C1(KEYINPUT30), .C2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT31), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n530), .A2(new_n531), .A3(new_n521), .A4(new_n500), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT71), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n532), .A2(new_n533), .ZN(new_n536));
  OAI22_X1  g350(.A1(new_n525), .A2(new_n526), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n500), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n521), .A2(new_n520), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n517), .A2(new_n512), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n509), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n520), .B1(new_n541), .B2(new_n521), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n539), .B1(new_n542), .B2(new_n523), .ZN(new_n543));
  INV_X1    g357(.A(new_n524), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n526), .B(new_n538), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n530), .A2(new_n521), .A3(new_n500), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT31), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n496), .B1(new_n537), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(G472), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n519), .A2(KEYINPUT72), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT29), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n551), .A2(new_n552), .A3(new_n524), .A4(new_n539), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT74), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n510), .B1(new_n508), .B2(new_n512), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n554), .B(KEYINPUT28), .C1(new_n513), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n508), .A2(new_n512), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n509), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n520), .B1(new_n558), .B2(new_n521), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n539), .A2(KEYINPUT74), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n556), .B(KEYINPUT29), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n553), .A2(new_n500), .A3(new_n561), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n530), .A2(new_n552), .A3(new_n521), .A4(new_n538), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n563), .A2(new_n239), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n550), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n538), .B1(new_n543), .B2(new_n544), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n530), .A2(new_n521), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n568), .A2(KEYINPUT71), .A3(new_n531), .A4(new_n500), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n567), .A2(KEYINPUT73), .B1(new_n569), .B2(new_n534), .ZN(new_n570));
  INV_X1    g384(.A(new_n547), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n571), .B1(new_n525), .B2(new_n526), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n494), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n549), .B(new_n566), .C1(new_n573), .C2(KEYINPUT32), .ZN(new_n574));
  INV_X1    g388(.A(new_n282), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n575), .B1(G234), .B2(new_n239), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n199), .A2(new_n200), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT23), .B1(new_n264), .B2(G119), .ZN(new_n578));
  OAI21_X1  g392(.A(KEYINPUT76), .B1(new_n340), .B2(G128), .ZN(new_n579));
  XOR2_X1   g393(.A(new_n578), .B(new_n579), .Z(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(G110), .ZN(new_n581));
  XOR2_X1   g395(.A(G119), .B(G128), .Z(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT24), .B(G110), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n577), .B(new_n581), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n583), .ZN(new_n585));
  OR2_X1    g399(.A1(new_n585), .A2(KEYINPUT78), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(KEYINPUT78), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n586), .B(new_n587), .C1(G110), .C2(new_n580), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(new_n200), .A3(new_n222), .ZN(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT22), .B(G137), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n243), .A2(G221), .A3(G234), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n584), .A2(new_n589), .A3(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n592), .B1(new_n584), .B2(new_n589), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(KEYINPUT25), .B1(new_n596), .B2(new_n239), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT25), .ZN(new_n598));
  NOR4_X1   g412(.A1(new_n594), .A2(new_n595), .A3(new_n598), .A4(G902), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n576), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n576), .A2(G902), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(KEYINPUT79), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n596), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n492), .A2(new_n574), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G101), .ZN(G3));
  NAND2_X1  g421(.A1(new_n567), .A2(KEYINPUT73), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n569), .A2(new_n534), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n608), .A2(new_n547), .A3(new_n545), .A4(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n550), .B1(new_n610), .B2(new_n239), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT95), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n573), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n605), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n614), .A2(new_n489), .A3(new_n491), .ZN(new_n615));
  AOI21_X1  g429(.A(G902), .B1(new_n570), .B2(new_n572), .ZN(new_n616));
  OAI21_X1  g430(.A(KEYINPUT95), .B1(new_n616), .B2(new_n550), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n401), .A2(new_n311), .A3(new_n419), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n309), .B(new_n251), .C1(new_n618), .C2(new_n420), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n236), .A2(new_n238), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n241), .A2(G475), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n300), .A2(KEYINPUT33), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT33), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n285), .A2(new_n624), .A3(new_n287), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n623), .A2(new_n625), .A3(G478), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n288), .A2(new_n289), .ZN(new_n627));
  NAND2_X1  g441(.A1(G478), .A2(G902), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n622), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n619), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n613), .A2(new_n615), .A3(new_n617), .A4(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT34), .B(G104), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  INV_X1    g448(.A(new_n303), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n242), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n619), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n613), .A2(new_n615), .A3(new_n617), .A4(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT35), .B(G107), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  NAND2_X1  g454(.A1(new_n584), .A2(new_n589), .ZN(new_n641));
  INV_X1    g455(.A(new_n592), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n641), .B1(KEYINPUT36), .B2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n642), .A2(KEYINPUT36), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n584), .A2(new_n589), .A3(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n643), .A2(new_n603), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT96), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n600), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n613), .A2(new_n492), .A3(new_n617), .A4(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT37), .B(G110), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G12));
  NOR2_X1   g466(.A1(new_n489), .A2(new_n491), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n574), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n246), .B1(G900), .B2(new_n250), .ZN(new_n655));
  XOR2_X1   g469(.A(new_n655), .B(KEYINPUT97), .Z(new_n656));
  NOR2_X1   g470(.A1(new_n636), .A2(new_n656), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n423), .A2(new_n649), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G128), .ZN(G30));
  NAND2_X1  g474(.A1(new_n421), .A2(new_n422), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n635), .A2(new_n622), .ZN(new_n664));
  INV_X1    g478(.A(new_n649), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n309), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n663), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(KEYINPUT32), .B1(new_n610), .B2(new_n493), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n568), .A2(new_n538), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n558), .A2(new_n521), .A3(new_n538), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n239), .ZN(new_n671));
  OAI21_X1  g485(.A(G472), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n549), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n667), .B1(new_n668), .B2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT40), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n478), .A2(new_n488), .ZN(new_n676));
  INV_X1    g490(.A(new_n474), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT99), .ZN(new_n679));
  XOR2_X1   g493(.A(new_n656), .B(KEYINPUT39), .Z(new_n680));
  INV_X1    g494(.A(new_n491), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n678), .A2(new_n679), .A3(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n679), .B1(new_n678), .B2(new_n682), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n675), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n685), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n687), .A2(KEYINPUT40), .A3(new_n683), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n674), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(new_n266), .ZN(G45));
  NOR2_X1   g504(.A1(new_n630), .A2(new_n656), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n309), .B1(new_n618), .B2(new_n420), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n692), .A2(new_n665), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n654), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G146), .ZN(G48));
  NAND2_X1  g510(.A1(new_n486), .A2(new_n239), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(G469), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n676), .A2(new_n681), .A3(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n574), .A2(new_n605), .A3(new_n699), .A4(new_n631), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT41), .B(G113), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT100), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n700), .B(new_n702), .ZN(G15));
  INV_X1    g517(.A(KEYINPUT101), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n549), .A2(new_n566), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n605), .B1(new_n705), .B2(new_n668), .ZN(new_n706));
  AOI22_X1  g520(.A1(new_n478), .A2(new_n488), .B1(G469), .B2(new_n697), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(new_n637), .A3(new_n681), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n704), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n493), .B1(new_n537), .B2(new_n548), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n495), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n565), .B1(new_n610), .B2(new_n496), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n614), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n707), .A2(new_n681), .A3(new_n637), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n713), .A2(KEYINPUT101), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n709), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G116), .ZN(G18));
  NAND3_X1  g531(.A1(new_n676), .A2(new_n681), .A3(new_n698), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n308), .A2(new_n423), .A3(new_n649), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n574), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G119), .ZN(G21));
  OAI21_X1  g536(.A(new_n239), .B1(new_n537), .B2(new_n548), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(G472), .ZN(new_n724));
  OAI211_X1 g538(.A(new_n556), .B(new_n538), .C1(new_n559), .C2(new_n560), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n547), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(KEYINPUT102), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT102), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n725), .A2(new_n547), .A3(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n727), .A2(new_n609), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n493), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT103), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n730), .A2(KEYINPUT103), .A3(new_n493), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n724), .A2(new_n733), .A3(new_n605), .A4(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT104), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n664), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n635), .A2(new_n622), .A3(KEYINPUT104), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n739), .A2(new_n619), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n681), .A3(new_n707), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n735), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(new_n254), .ZN(G24));
  AOI21_X1  g557(.A(KEYINPUT103), .B1(new_n730), .B2(new_n493), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n611), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n745), .A2(new_n694), .A3(new_n699), .A4(new_n734), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G125), .ZN(G27));
  INV_X1    g561(.A(KEYINPUT42), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n421), .A2(new_n309), .A3(new_n422), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n678), .A2(new_n681), .A3(new_n691), .A4(new_n750), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n748), .B1(new_n706), .B2(new_n751), .ZN(new_n752));
  NOR4_X1   g566(.A1(new_n489), .A2(new_n692), .A3(new_n491), .A4(new_n749), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n713), .A2(KEYINPUT42), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G131), .ZN(G33));
  AND3_X1   g570(.A1(new_n653), .A2(new_n657), .A3(new_n750), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n713), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G134), .ZN(G36));
  NAND2_X1  g573(.A1(new_n613), .A2(new_n617), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n629), .A2(new_n242), .ZN(new_n761));
  NOR2_X1   g575(.A1(KEYINPUT107), .A2(KEYINPUT43), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(KEYINPUT107), .A2(KEYINPUT43), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n762), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n766), .A2(KEYINPUT108), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(KEYINPUT108), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n665), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n760), .A2(new_n769), .A3(KEYINPUT44), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n750), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT109), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT105), .B1(new_n473), .B2(new_n773), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n425), .B1(new_n473), .B2(new_n773), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT105), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n468), .A2(new_n472), .A3(new_n776), .A4(KEYINPUT45), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n774), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(KEYINPUT106), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT106), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n774), .A2(new_n775), .A3(new_n780), .A4(new_n777), .ZN(new_n781));
  AOI22_X1  g595(.A1(new_n779), .A2(new_n781), .B1(G469), .B2(G902), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT46), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n676), .B1(new_n782), .B2(KEYINPUT46), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n681), .B(new_n680), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT109), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n770), .A2(new_n788), .A3(new_n750), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n760), .A2(new_n769), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT44), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n772), .A2(new_n787), .A3(new_n789), .A4(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G137), .ZN(G39));
  OAI21_X1  g608(.A(new_n681), .B1(new_n784), .B2(new_n785), .ZN(new_n795));
  NOR2_X1   g609(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n796));
  NAND2_X1  g610(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n795), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n681), .B(new_n797), .C1(new_n784), .C2(new_n785), .ZN(new_n800));
  NOR4_X1   g614(.A1(new_n574), .A2(new_n605), .A3(new_n692), .A4(new_n749), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G140), .ZN(G42));
  NOR3_X1   g617(.A1(new_n489), .A2(new_n491), .A3(new_n749), .ZN(new_n804));
  NOR4_X1   g618(.A1(new_n665), .A2(new_n622), .A3(new_n635), .A4(new_n656), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n574), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n706), .A2(new_n748), .A3(new_n751), .ZN(new_n808));
  AOI21_X1  g622(.A(KEYINPUT42), .B1(new_n713), .B2(new_n753), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n807), .B(new_n758), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n730), .A2(KEYINPUT103), .A3(new_n493), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n611), .A2(new_n811), .A3(new_n744), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n812), .A2(KEYINPUT111), .A3(new_n649), .A4(new_n753), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT111), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n724), .A2(new_n733), .A3(new_n649), .A4(new_n734), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n814), .B1(new_n815), .B2(new_n751), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n810), .A2(new_n817), .ZN(new_n818));
  AND4_X1   g632(.A1(KEYINPUT101), .A2(new_n714), .A3(new_n574), .A4(new_n605), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT101), .B1(new_n713), .B2(new_n714), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n632), .B(new_n638), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  AOI22_X1  g635(.A1(new_n713), .A2(new_n492), .B1(new_n720), .B2(new_n574), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n718), .A2(new_n619), .A3(new_n739), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n812), .A2(new_n605), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n822), .A2(new_n824), .A3(new_n650), .A4(new_n700), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n821), .A2(new_n825), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n574), .B(new_n653), .C1(new_n658), .C2(new_n694), .ZN(new_n827));
  NOR4_X1   g641(.A1(new_n739), .A2(new_n693), .A3(new_n649), .A4(new_n656), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n828), .B(new_n653), .C1(new_n668), .C2(new_n673), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n746), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n746), .A2(new_n827), .A3(KEYINPUT52), .A4(new_n829), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n818), .A2(new_n826), .A3(KEYINPUT53), .A4(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT113), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n838));
  AOI221_X4 g652(.A(new_n806), .B1(new_n713), .B2(new_n757), .C1(new_n752), .C2(new_n754), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n723), .A2(new_n612), .A3(G472), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n617), .A2(new_n710), .A3(new_n840), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n841), .B(new_n615), .C1(new_n631), .C2(new_n637), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n716), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n825), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n813), .A2(new_n816), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n839), .A2(new_n843), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT112), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n832), .A2(new_n847), .A3(new_n833), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n830), .A2(KEYINPUT112), .A3(new_n831), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n838), .B1(new_n846), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n617), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n840), .A2(new_n710), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n693), .B1(new_n306), .B2(new_n307), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n678), .A2(new_n854), .A3(new_n681), .A4(new_n649), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n852), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(new_n742), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n606), .A2(new_n700), .A3(new_n721), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n857), .A2(new_n716), .A3(new_n858), .A4(new_n842), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n845), .A2(new_n755), .A3(new_n758), .A4(new_n807), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(KEYINPUT113), .A3(KEYINPUT53), .A4(new_n834), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n837), .A2(new_n851), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT54), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n861), .A2(KEYINPUT53), .A3(new_n849), .A4(new_n848), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n818), .A2(new_n826), .A3(new_n834), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n838), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n865), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT114), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n865), .A2(new_n867), .A3(KEYINPUT114), .A4(new_n868), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n718), .A2(new_n246), .A3(new_n749), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n873), .B1(new_n763), .B2(new_n765), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n874), .A2(new_n706), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT48), .Z(new_n876));
  NOR3_X1   g690(.A1(new_n735), .A2(new_n246), .A3(new_n766), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(new_n423), .A3(new_n699), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n673), .A2(new_n668), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n873), .A2(new_n605), .A3(new_n879), .ZN(new_n880));
  OR2_X1    g694(.A1(new_n880), .A2(new_n630), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n244), .B(KEYINPUT116), .Z(new_n882));
  NAND4_X1  g696(.A1(new_n876), .A2(new_n878), .A3(new_n881), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n877), .A2(new_n750), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n779), .A2(new_n781), .ZN(new_n885));
  NAND2_X1  g699(.A1(G469), .A2(G902), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT46), .ZN(new_n888));
  AOI22_X1  g702(.A1(new_n887), .A2(new_n888), .B1(new_n488), .B2(new_n478), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n491), .B1(new_n889), .B2(new_n783), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n798), .A2(new_n796), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n800), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n707), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n893), .A2(new_n681), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n884), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n622), .A2(new_n629), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  OAI22_X1  g712(.A1(new_n874), .A2(new_n815), .B1(new_n880), .B2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n699), .A2(new_n310), .A3(new_n663), .ZN(new_n901));
  NOR4_X1   g715(.A1(new_n901), .A2(new_n735), .A3(new_n246), .A4(new_n766), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n902), .A2(KEYINPUT115), .A3(KEYINPUT50), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT50), .ZN(new_n904));
  INV_X1    g718(.A(new_n901), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n877), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT115), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n900), .B1(new_n903), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT51), .B1(new_n896), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT51), .ZN(new_n911));
  OAI21_X1  g725(.A(KEYINPUT50), .B1(new_n902), .B2(KEYINPUT115), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n906), .A2(new_n907), .A3(new_n904), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n899), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n894), .B1(new_n799), .B2(new_n800), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n911), .B(new_n914), .C1(new_n915), .C2(new_n884), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n883), .B1(new_n910), .B2(new_n916), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n864), .A2(new_n871), .A3(new_n872), .A4(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(G952), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n243), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n707), .B(KEYINPUT49), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n605), .A2(new_n681), .A3(new_n309), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n923), .A2(new_n761), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n922), .A2(new_n879), .A3(new_n663), .A4(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n921), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(KEYINPUT117), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT117), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n921), .A2(new_n928), .A3(new_n925), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n927), .A2(new_n929), .ZN(G75));
  AND2_X1   g744(.A1(new_n865), .A2(new_n867), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n931), .A2(new_n239), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(G210), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT56), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n377), .A2(new_n400), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(new_n399), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT55), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n933), .A2(new_n934), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n937), .B1(new_n933), .B2(new_n934), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n919), .A2(G953), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT118), .Z(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n938), .A2(new_n939), .A3(new_n942), .ZN(G51));
  NAND2_X1  g757(.A1(new_n865), .A2(new_n867), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(KEYINPUT54), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n869), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n886), .B(KEYINPUT57), .Z(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(new_n486), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n932), .A2(new_n781), .A3(new_n779), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n942), .B1(new_n949), .B2(new_n950), .ZN(G54));
  NAND3_X1  g765(.A1(new_n932), .A2(KEYINPUT58), .A3(G475), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n228), .A2(new_n234), .ZN(new_n953));
  OR2_X1    g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n952), .A2(new_n953), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n942), .B1(new_n954), .B2(new_n955), .ZN(G60));
  AND2_X1   g770(.A1(new_n623), .A2(new_n625), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n628), .B(KEYINPUT59), .Z(new_n958));
  AOI211_X1 g772(.A(new_n957), .B(new_n958), .C1(new_n945), .C2(new_n869), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n864), .A2(new_n871), .A3(new_n872), .ZN(new_n960));
  INV_X1    g774(.A(new_n958), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI211_X1 g776(.A(new_n942), .B(new_n959), .C1(new_n962), .C2(new_n957), .ZN(G63));
  INV_X1    g777(.A(KEYINPUT61), .ZN(new_n964));
  NAND2_X1  g778(.A1(G217), .A2(G902), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT60), .ZN(new_n966));
  OAI21_X1  g780(.A(KEYINPUT119), .B1(new_n931), .B2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n596), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT119), .ZN(new_n969));
  INV_X1    g783(.A(new_n966), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n944), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n967), .A2(new_n968), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n941), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n643), .A2(new_n645), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n975), .B1(new_n967), .B2(new_n971), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n964), .B1(new_n973), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n976), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n978), .A2(KEYINPUT61), .A3(new_n941), .A4(new_n972), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n977), .A2(new_n979), .ZN(G66));
  NAND3_X1  g794(.A1(new_n248), .A2(G224), .A3(G953), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n981), .B1(new_n859), .B2(G953), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n935), .B1(G898), .B2(new_n243), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT120), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n982), .B(new_n984), .ZN(G69));
  OAI21_X1  g799(.A(new_n527), .B1(KEYINPUT30), .B2(new_n529), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(new_n232), .ZN(new_n987));
  XNOR2_X1  g801(.A(KEYINPUT121), .B(KEYINPUT122), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT123), .Z(new_n990));
  NAND2_X1  g804(.A1(new_n746), .A2(new_n827), .ZN(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n686), .A2(new_n688), .ZN(new_n993));
  OAI211_X1 g807(.A(KEYINPUT62), .B(new_n992), .C1(new_n993), .C2(new_n674), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT62), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n995), .B1(new_n689), .B2(new_n991), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n749), .B1(new_n630), .B2(new_n636), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n687), .A2(new_n713), .A3(new_n683), .A4(new_n998), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n997), .A2(new_n793), .A3(new_n802), .A4(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n990), .B1(new_n1000), .B2(new_n243), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n992), .A2(new_n755), .A3(new_n758), .ZN(new_n1002));
  NOR3_X1   g816(.A1(new_n706), .A2(new_n693), .A3(new_n739), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1002), .B1(new_n787), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n1004), .A2(new_n793), .A3(new_n802), .ZN(new_n1005));
  OR2_X1    g819(.A1(new_n1005), .A2(G953), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n989), .B1(G900), .B2(G953), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1001), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n243), .B1(G227), .B2(G900), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1008), .B(new_n1009), .Z(G72));
  INV_X1    g824(.A(KEYINPUT127), .ZN(new_n1011));
  INV_X1    g825(.A(new_n568), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n1012), .A2(new_n500), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(new_n669), .ZN(new_n1015));
  NAND2_X1  g829(.A1(G472), .A2(G902), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n1016), .B(KEYINPUT63), .Z(new_n1017));
  NAND3_X1  g831(.A1(new_n1014), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  XOR2_X1   g832(.A(new_n1018), .B(KEYINPUT125), .Z(new_n1019));
  NAND2_X1  g833(.A1(new_n863), .A2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1020), .B(KEYINPUT126), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1017), .B1(new_n1005), .B2(new_n859), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n942), .B1(new_n1022), .B2(new_n1013), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1017), .B1(new_n1000), .B2(new_n859), .ZN(new_n1024));
  AND3_X1   g838(.A1(new_n1024), .A2(KEYINPUT124), .A3(new_n669), .ZN(new_n1025));
  AOI21_X1  g839(.A(KEYINPUT124), .B1(new_n1024), .B2(new_n669), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1023), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1011), .B1(new_n1021), .B2(new_n1027), .ZN(new_n1028));
  OR2_X1    g842(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1029));
  INV_X1    g843(.A(KEYINPUT126), .ZN(new_n1030));
  XNOR2_X1  g844(.A(new_n1020), .B(new_n1030), .ZN(new_n1031));
  NAND4_X1  g845(.A1(new_n1029), .A2(new_n1031), .A3(KEYINPUT127), .A4(new_n1023), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1028), .A2(new_n1032), .ZN(G57));
endmodule


