

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U547 ( .A(n542), .B(n541), .ZN(G160) );
  NOR2_X1 U548 ( .A1(G651), .A2(G543), .ZN(n789) );
  NOR2_X1 U549 ( .A1(n511), .A2(n730), .ZN(n731) );
  AND2_X1 U550 ( .A1(n747), .A2(n717), .ZN(n511) );
  AND2_X1 U551 ( .A1(n634), .A2(G1996), .ZN(n612) );
  NOR2_X1 U552 ( .A1(n1006), .A2(n615), .ZN(n621) );
  NOR2_X1 U553 ( .A1(n645), .A2(n644), .ZN(n647) );
  AND2_X1 U554 ( .A1(n657), .A2(n656), .ZN(n658) );
  INV_X1 U555 ( .A(n634), .ZN(n650) );
  NAND2_X1 U556 ( .A1(G8), .A2(n650), .ZN(n682) );
  NOR2_X1 U557 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U558 ( .A1(G164), .A2(G1384), .ZN(n695) );
  AND2_X1 U559 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U560 ( .A1(G2105), .A2(G2104), .ZN(n512) );
  NOR2_X1 U561 ( .A1(G651), .A2(n581), .ZN(n786) );
  NOR2_X1 U562 ( .A1(n520), .A2(n519), .ZN(G164) );
  INV_X1 U563 ( .A(G2104), .ZN(n516) );
  NOR2_X2 U564 ( .A1(G2105), .A2(n516), .ZN(n989) );
  NAND2_X1 U565 ( .A1(n989), .A2(G102), .ZN(n515) );
  XOR2_X2 U566 ( .A(KEYINPUT17), .B(n512), .Z(n988) );
  NAND2_X1 U567 ( .A1(n988), .A2(G138), .ZN(n513) );
  XOR2_X1 U568 ( .A(KEYINPUT85), .B(n513), .Z(n514) );
  NAND2_X1 U569 ( .A1(n515), .A2(n514), .ZN(n520) );
  AND2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n984) );
  NAND2_X1 U571 ( .A1(G114), .A2(n984), .ZN(n518) );
  AND2_X1 U572 ( .A1(n516), .A2(G2105), .ZN(n985) );
  NAND2_X1 U573 ( .A1(G126), .A2(n985), .ZN(n517) );
  NAND2_X1 U574 ( .A1(n518), .A2(n517), .ZN(n519) );
  XOR2_X1 U575 ( .A(KEYINPUT0), .B(G543), .Z(n581) );
  NAND2_X1 U576 ( .A1(G48), .A2(n786), .ZN(n521) );
  XNOR2_X1 U577 ( .A(n521), .B(KEYINPUT80), .ZN(n531) );
  INV_X1 U578 ( .A(G651), .ZN(n525) );
  NOR2_X1 U579 ( .A1(G543), .A2(n525), .ZN(n522) );
  XOR2_X1 U580 ( .A(KEYINPUT1), .B(n522), .Z(n785) );
  NAND2_X1 U581 ( .A1(G61), .A2(n785), .ZN(n524) );
  NAND2_X1 U582 ( .A1(G86), .A2(n789), .ZN(n523) );
  NAND2_X1 U583 ( .A1(n524), .A2(n523), .ZN(n529) );
  OR2_X1 U584 ( .A1(n525), .A2(n581), .ZN(n526) );
  XOR2_X1 U585 ( .A(KEYINPUT68), .B(n526), .Z(n790) );
  NAND2_X1 U586 ( .A1(n790), .A2(G73), .ZN(n527) );
  XOR2_X1 U587 ( .A(KEYINPUT2), .B(n527), .Z(n528) );
  NOR2_X1 U588 ( .A1(n529), .A2(n528), .ZN(n530) );
  NAND2_X1 U589 ( .A1(n531), .A2(n530), .ZN(G305) );
  NAND2_X1 U590 ( .A1(G137), .A2(n988), .ZN(n532) );
  XNOR2_X1 U591 ( .A(n532), .B(KEYINPUT66), .ZN(n540) );
  XOR2_X1 U592 ( .A(KEYINPUT23), .B(KEYINPUT65), .Z(n534) );
  NAND2_X1 U593 ( .A1(G101), .A2(n989), .ZN(n533) );
  XNOR2_X1 U594 ( .A(n534), .B(n533), .ZN(n538) );
  NAND2_X1 U595 ( .A1(G113), .A2(n984), .ZN(n536) );
  NAND2_X1 U596 ( .A1(G125), .A2(n985), .ZN(n535) );
  NAND2_X1 U597 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U598 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U599 ( .A1(n540), .A2(n539), .ZN(n542) );
  INV_X1 U600 ( .A(KEYINPUT64), .ZN(n541) );
  NAND2_X1 U601 ( .A1(G91), .A2(n789), .ZN(n544) );
  NAND2_X1 U602 ( .A1(G78), .A2(n790), .ZN(n543) );
  NAND2_X1 U603 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U604 ( .A(KEYINPUT72), .B(n545), .Z(n549) );
  NAND2_X1 U605 ( .A1(G65), .A2(n785), .ZN(n547) );
  NAND2_X1 U606 ( .A1(G53), .A2(n786), .ZN(n546) );
  AND2_X1 U607 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U608 ( .A1(n549), .A2(n548), .ZN(G299) );
  NAND2_X1 U609 ( .A1(G90), .A2(n789), .ZN(n551) );
  NAND2_X1 U610 ( .A1(G77), .A2(n790), .ZN(n550) );
  NAND2_X1 U611 ( .A1(n551), .A2(n550), .ZN(n553) );
  XOR2_X1 U612 ( .A(KEYINPUT71), .B(KEYINPUT9), .Z(n552) );
  XNOR2_X1 U613 ( .A(n553), .B(n552), .ZN(n558) );
  NAND2_X1 U614 ( .A1(G64), .A2(n785), .ZN(n555) );
  NAND2_X1 U615 ( .A1(G52), .A2(n786), .ZN(n554) );
  NAND2_X1 U616 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U617 ( .A(KEYINPUT70), .B(n556), .Z(n557) );
  NAND2_X1 U618 ( .A1(n558), .A2(n557), .ZN(G301) );
  INV_X1 U619 ( .A(G301), .ZN(G171) );
  NAND2_X1 U620 ( .A1(G89), .A2(n789), .ZN(n559) );
  XNOR2_X1 U621 ( .A(n559), .B(KEYINPUT76), .ZN(n560) );
  XNOR2_X1 U622 ( .A(KEYINPUT4), .B(n560), .ZN(n563) );
  NAND2_X1 U623 ( .A1(G76), .A2(n790), .ZN(n561) );
  XOR2_X1 U624 ( .A(KEYINPUT77), .B(n561), .Z(n562) );
  NAND2_X1 U625 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U626 ( .A(KEYINPUT5), .B(n564), .ZN(n570) );
  NAND2_X1 U627 ( .A1(n786), .A2(G51), .ZN(n565) );
  XNOR2_X1 U628 ( .A(n565), .B(KEYINPUT78), .ZN(n567) );
  NAND2_X1 U629 ( .A1(G63), .A2(n785), .ZN(n566) );
  NAND2_X1 U630 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U631 ( .A(KEYINPUT6), .B(n568), .Z(n569) );
  NAND2_X1 U632 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U633 ( .A(KEYINPUT7), .B(n571), .ZN(G168) );
  XOR2_X1 U634 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U635 ( .A1(G88), .A2(n789), .ZN(n573) );
  NAND2_X1 U636 ( .A1(G75), .A2(n790), .ZN(n572) );
  NAND2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n577) );
  NAND2_X1 U638 ( .A1(G62), .A2(n785), .ZN(n575) );
  NAND2_X1 U639 ( .A1(G50), .A2(n786), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U641 ( .A1(n577), .A2(n576), .ZN(G166) );
  INV_X1 U642 ( .A(G166), .ZN(G303) );
  NAND2_X1 U643 ( .A1(G49), .A2(n786), .ZN(n579) );
  NAND2_X1 U644 ( .A1(G74), .A2(G651), .ZN(n578) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U646 ( .A1(n785), .A2(n580), .ZN(n583) );
  NAND2_X1 U647 ( .A1(n581), .A2(G87), .ZN(n582) );
  NAND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(G288) );
  NAND2_X1 U649 ( .A1(G60), .A2(n785), .ZN(n585) );
  NAND2_X1 U650 ( .A1(G47), .A2(n786), .ZN(n584) );
  NAND2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U652 ( .A(KEYINPUT69), .B(n586), .Z(n589) );
  NAND2_X1 U653 ( .A1(G85), .A2(n789), .ZN(n587) );
  XNOR2_X1 U654 ( .A(KEYINPUT67), .B(n587), .ZN(n588) );
  NOR2_X1 U655 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U656 ( .A1(G72), .A2(n790), .ZN(n590) );
  NAND2_X1 U657 ( .A1(n591), .A2(n590), .ZN(G290) );
  XOR2_X1 U658 ( .A(G1981), .B(G305), .Z(n849) );
  NAND2_X1 U659 ( .A1(G66), .A2(n785), .ZN(n593) );
  NAND2_X1 U660 ( .A1(G92), .A2(n789), .ZN(n592) );
  NAND2_X1 U661 ( .A1(n593), .A2(n592), .ZN(n597) );
  NAND2_X1 U662 ( .A1(G54), .A2(n786), .ZN(n595) );
  NAND2_X1 U663 ( .A1(G79), .A2(n790), .ZN(n594) );
  NAND2_X1 U664 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U665 ( .A1(n597), .A2(n596), .ZN(n599) );
  XNOR2_X1 U666 ( .A(KEYINPUT74), .B(KEYINPUT75), .ZN(n598) );
  XNOR2_X1 U667 ( .A(n599), .B(n598), .ZN(n600) );
  XOR2_X1 U668 ( .A(KEYINPUT15), .B(n600), .Z(n763) );
  INV_X1 U669 ( .A(n763), .ZN(n1003) );
  NAND2_X1 U670 ( .A1(G56), .A2(n785), .ZN(n601) );
  XOR2_X1 U671 ( .A(KEYINPUT14), .B(n601), .Z(n607) );
  NAND2_X1 U672 ( .A1(n789), .A2(G81), .ZN(n602) );
  XNOR2_X1 U673 ( .A(n602), .B(KEYINPUT12), .ZN(n604) );
  NAND2_X1 U674 ( .A1(G68), .A2(n790), .ZN(n603) );
  NAND2_X1 U675 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U676 ( .A(KEYINPUT13), .B(n605), .Z(n606) );
  NOR2_X1 U677 ( .A1(n607), .A2(n606), .ZN(n609) );
  NAND2_X1 U678 ( .A1(n786), .A2(G43), .ZN(n608) );
  NAND2_X1 U679 ( .A1(n609), .A2(n608), .ZN(n1006) );
  INV_X1 U680 ( .A(n695), .ZN(n610) );
  NAND2_X1 U681 ( .A1(G40), .A2(G160), .ZN(n696) );
  NOR2_X4 U682 ( .A1(n610), .A2(n696), .ZN(n634) );
  INV_X1 U683 ( .A(KEYINPUT26), .ZN(n611) );
  XNOR2_X1 U684 ( .A(n612), .B(n611), .ZN(n614) );
  NAND2_X1 U685 ( .A1(n650), .A2(G1341), .ZN(n613) );
  NAND2_X1 U686 ( .A1(n614), .A2(n613), .ZN(n615) );
  NAND2_X1 U687 ( .A1(n1003), .A2(n621), .ZN(n620) );
  INV_X1 U688 ( .A(G1348), .ZN(n835) );
  NOR2_X1 U689 ( .A1(n634), .A2(n835), .ZN(n616) );
  XNOR2_X1 U690 ( .A(n616), .B(KEYINPUT97), .ZN(n618) );
  NAND2_X1 U691 ( .A1(n634), .A2(G2067), .ZN(n617) );
  NAND2_X1 U692 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U693 ( .A1(n620), .A2(n619), .ZN(n623) );
  OR2_X1 U694 ( .A1(n1003), .A2(n621), .ZN(n622) );
  NAND2_X1 U695 ( .A1(n623), .A2(n622), .ZN(n628) );
  INV_X1 U696 ( .A(G299), .ZN(n803) );
  NAND2_X1 U697 ( .A1(n634), .A2(G2072), .ZN(n624) );
  XNOR2_X1 U698 ( .A(n624), .B(KEYINPUT27), .ZN(n626) );
  INV_X1 U699 ( .A(G1956), .ZN(n962) );
  NOR2_X1 U700 ( .A1(n962), .A2(n634), .ZN(n625) );
  NOR2_X1 U701 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U702 ( .A1(n803), .A2(n629), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n628), .A2(n627), .ZN(n632) );
  NOR2_X1 U704 ( .A1(n803), .A2(n629), .ZN(n630) );
  XOR2_X1 U705 ( .A(n630), .B(KEYINPUT28), .Z(n631) );
  NAND2_X1 U706 ( .A1(n632), .A2(n631), .ZN(n633) );
  XOR2_X1 U707 ( .A(KEYINPUT29), .B(n633), .Z(n639) );
  INV_X1 U708 ( .A(G1961), .ZN(n963) );
  NAND2_X1 U709 ( .A1(n650), .A2(n963), .ZN(n636) );
  XNOR2_X1 U710 ( .A(G2078), .B(KEYINPUT25), .ZN(n923) );
  NAND2_X1 U711 ( .A1(n634), .A2(n923), .ZN(n635) );
  NAND2_X1 U712 ( .A1(n636), .A2(n635), .ZN(n640) );
  AND2_X1 U713 ( .A1(n640), .A2(G171), .ZN(n637) );
  XOR2_X1 U714 ( .A(KEYINPUT96), .B(n637), .Z(n638) );
  NAND2_X1 U715 ( .A1(n639), .A2(n638), .ZN(n649) );
  NOR2_X1 U716 ( .A1(G171), .A2(n640), .ZN(n645) );
  NOR2_X1 U717 ( .A1(G1966), .A2(n682), .ZN(n662) );
  NOR2_X1 U718 ( .A1(G2084), .A2(n650), .ZN(n659) );
  NOR2_X1 U719 ( .A1(n662), .A2(n659), .ZN(n641) );
  NAND2_X1 U720 ( .A1(G8), .A2(n641), .ZN(n642) );
  XNOR2_X1 U721 ( .A(KEYINPUT30), .B(n642), .ZN(n643) );
  NOR2_X1 U722 ( .A1(G168), .A2(n643), .ZN(n644) );
  XOR2_X1 U723 ( .A(KEYINPUT31), .B(KEYINPUT98), .Z(n646) );
  XNOR2_X1 U724 ( .A(n647), .B(n646), .ZN(n648) );
  NAND2_X1 U725 ( .A1(n649), .A2(n648), .ZN(n660) );
  NAND2_X1 U726 ( .A1(n660), .A2(G286), .ZN(n657) );
  INV_X1 U727 ( .A(G8), .ZN(n655) );
  NOR2_X1 U728 ( .A1(G1971), .A2(n682), .ZN(n652) );
  NOR2_X1 U729 ( .A1(G2090), .A2(n650), .ZN(n651) );
  NOR2_X1 U730 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U731 ( .A1(n653), .A2(G303), .ZN(n654) );
  OR2_X1 U732 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U733 ( .A(n658), .B(KEYINPUT32), .ZN(n666) );
  NAND2_X1 U734 ( .A1(G8), .A2(n659), .ZN(n664) );
  INV_X1 U735 ( .A(n660), .ZN(n661) );
  NOR2_X1 U736 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U737 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U738 ( .A1(n666), .A2(n665), .ZN(n686) );
  NOR2_X1 U739 ( .A1(G1976), .A2(G288), .ZN(n675) );
  NOR2_X1 U740 ( .A1(G1971), .A2(G303), .ZN(n667) );
  NOR2_X1 U741 ( .A1(n675), .A2(n667), .ZN(n841) );
  XOR2_X1 U742 ( .A(n841), .B(KEYINPUT99), .Z(n669) );
  INV_X1 U743 ( .A(KEYINPUT33), .ZN(n668) );
  AND2_X1 U744 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U745 ( .A1(n686), .A2(n670), .ZN(n674) );
  NAND2_X1 U746 ( .A1(G1976), .A2(G288), .ZN(n840) );
  INV_X1 U747 ( .A(n840), .ZN(n671) );
  NOR2_X1 U748 ( .A1(n682), .A2(n671), .ZN(n672) );
  OR2_X1 U749 ( .A1(KEYINPUT33), .A2(n672), .ZN(n673) );
  NAND2_X1 U750 ( .A1(n674), .A2(n673), .ZN(n678) );
  NAND2_X1 U751 ( .A1(n675), .A2(KEYINPUT33), .ZN(n676) );
  NOR2_X1 U752 ( .A1(n676), .A2(n682), .ZN(n677) );
  NAND2_X1 U753 ( .A1(n849), .A2(n679), .ZN(n694) );
  NOR2_X1 U754 ( .A1(G1981), .A2(G305), .ZN(n680) );
  XOR2_X1 U755 ( .A(n680), .B(KEYINPUT24), .Z(n681) );
  NOR2_X1 U756 ( .A1(n682), .A2(n681), .ZN(n692) );
  INV_X1 U757 ( .A(n682), .ZN(n690) );
  NOR2_X1 U758 ( .A1(G2090), .A2(G303), .ZN(n683) );
  XNOR2_X1 U759 ( .A(KEYINPUT100), .B(n683), .ZN(n684) );
  NAND2_X1 U760 ( .A1(n684), .A2(G8), .ZN(n685) );
  XNOR2_X1 U761 ( .A(KEYINPUT101), .B(n685), .ZN(n688) );
  INV_X1 U762 ( .A(n686), .ZN(n687) );
  NOR2_X1 U763 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U764 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U765 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U766 ( .A1(n694), .A2(n693), .ZN(n732) );
  NOR2_X1 U767 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U768 ( .A(n697), .B(KEYINPUT86), .ZN(n747) );
  XOR2_X1 U769 ( .A(KEYINPUT94), .B(KEYINPUT38), .Z(n699) );
  NAND2_X1 U770 ( .A1(G105), .A2(n989), .ZN(n698) );
  XNOR2_X1 U771 ( .A(n699), .B(n698), .ZN(n703) );
  NAND2_X1 U772 ( .A1(G141), .A2(n988), .ZN(n701) );
  NAND2_X1 U773 ( .A1(G117), .A2(n984), .ZN(n700) );
  NAND2_X1 U774 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U775 ( .A1(n703), .A2(n702), .ZN(n705) );
  NAND2_X1 U776 ( .A1(n985), .A2(G129), .ZN(n704) );
  NAND2_X1 U777 ( .A1(n705), .A2(n704), .ZN(n980) );
  NAND2_X1 U778 ( .A1(n980), .A2(G1996), .ZN(n706) );
  XNOR2_X1 U779 ( .A(n706), .B(KEYINPUT95), .ZN(n891) );
  NAND2_X1 U780 ( .A1(G119), .A2(n985), .ZN(n715) );
  NAND2_X1 U781 ( .A1(n988), .A2(G131), .ZN(n707) );
  XOR2_X1 U782 ( .A(KEYINPUT91), .B(n707), .Z(n709) );
  NAND2_X1 U783 ( .A1(n989), .A2(G95), .ZN(n708) );
  NAND2_X1 U784 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U785 ( .A(KEYINPUT92), .B(n710), .ZN(n713) );
  NAND2_X1 U786 ( .A1(n984), .A2(G107), .ZN(n711) );
  XOR2_X1 U787 ( .A(KEYINPUT90), .B(n711), .Z(n712) );
  NOR2_X1 U788 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U789 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U790 ( .A(n716), .B(KEYINPUT93), .Z(n999) );
  AND2_X1 U791 ( .A1(n999), .A2(G1991), .ZN(n887) );
  OR2_X1 U792 ( .A1(n891), .A2(n887), .ZN(n717) );
  NAND2_X1 U793 ( .A1(G140), .A2(n988), .ZN(n719) );
  NAND2_X1 U794 ( .A1(G104), .A2(n989), .ZN(n718) );
  NAND2_X1 U795 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U796 ( .A(KEYINPUT34), .B(n720), .ZN(n726) );
  NAND2_X1 U797 ( .A1(n984), .A2(G116), .ZN(n721) );
  XOR2_X1 U798 ( .A(KEYINPUT87), .B(n721), .Z(n723) );
  NAND2_X1 U799 ( .A1(n985), .A2(G128), .ZN(n722) );
  NAND2_X1 U800 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U801 ( .A(n724), .B(KEYINPUT35), .Z(n725) );
  NOR2_X1 U802 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U803 ( .A(KEYINPUT36), .B(n727), .Z(n728) );
  XNOR2_X1 U804 ( .A(KEYINPUT88), .B(n728), .ZN(n977) );
  XOR2_X1 U805 ( .A(G2067), .B(KEYINPUT37), .Z(n736) );
  NAND2_X1 U806 ( .A1(n977), .A2(n736), .ZN(n729) );
  XNOR2_X1 U807 ( .A(n729), .B(KEYINPUT89), .ZN(n916) );
  NAND2_X1 U808 ( .A1(n916), .A2(n747), .ZN(n744) );
  INV_X1 U809 ( .A(n744), .ZN(n730) );
  XNOR2_X1 U810 ( .A(KEYINPUT102), .B(n733), .ZN(n735) );
  XNOR2_X1 U811 ( .A(G1986), .B(G290), .ZN(n837) );
  NAND2_X1 U812 ( .A1(n837), .A2(n747), .ZN(n734) );
  NAND2_X1 U813 ( .A1(n735), .A2(n734), .ZN(n750) );
  NOR2_X1 U814 ( .A1(n977), .A2(n736), .ZN(n737) );
  XNOR2_X1 U815 ( .A(n737), .B(KEYINPUT105), .ZN(n897) );
  NOR2_X1 U816 ( .A1(G1996), .A2(n980), .ZN(n889) );
  NOR2_X1 U817 ( .A1(G1991), .A2(n999), .ZN(n886) );
  NOR2_X1 U818 ( .A1(G1986), .A2(G290), .ZN(n738) );
  XOR2_X1 U819 ( .A(n738), .B(KEYINPUT103), .Z(n739) );
  NOR2_X1 U820 ( .A1(n886), .A2(n739), .ZN(n740) );
  NOR2_X1 U821 ( .A1(n511), .A2(n740), .ZN(n741) );
  NOR2_X1 U822 ( .A1(n889), .A2(n741), .ZN(n742) );
  XNOR2_X1 U823 ( .A(KEYINPUT104), .B(n742), .ZN(n743) );
  XNOR2_X1 U824 ( .A(n743), .B(KEYINPUT39), .ZN(n745) );
  NAND2_X1 U825 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U826 ( .A1(n897), .A2(n746), .ZN(n748) );
  NAND2_X1 U827 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U828 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U829 ( .A(n751), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U830 ( .A(G2443), .B(G2446), .Z(n753) );
  XNOR2_X1 U831 ( .A(G2427), .B(G2451), .ZN(n752) );
  XNOR2_X1 U832 ( .A(n753), .B(n752), .ZN(n759) );
  XOR2_X1 U833 ( .A(G2430), .B(G2454), .Z(n755) );
  XOR2_X1 U834 ( .A(G1341), .B(n835), .Z(n754) );
  XNOR2_X1 U835 ( .A(n755), .B(n754), .ZN(n757) );
  XOR2_X1 U836 ( .A(G2435), .B(G2438), .Z(n756) );
  XNOR2_X1 U837 ( .A(n757), .B(n756), .ZN(n758) );
  XOR2_X1 U838 ( .A(n759), .B(n758), .Z(n760) );
  AND2_X1 U839 ( .A1(G14), .A2(n760), .ZN(G401) );
  AND2_X1 U840 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U841 ( .A(G57), .ZN(G237) );
  INV_X1 U842 ( .A(G82), .ZN(G220) );
  NAND2_X1 U843 ( .A1(G7), .A2(G661), .ZN(n761) );
  XOR2_X1 U844 ( .A(n761), .B(KEYINPUT10), .Z(n1017) );
  NAND2_X1 U845 ( .A1(n1017), .A2(G567), .ZN(n762) );
  XOR2_X1 U846 ( .A(KEYINPUT11), .B(n762), .Z(G234) );
  INV_X1 U847 ( .A(G860), .ZN(n769) );
  OR2_X1 U848 ( .A1(n1006), .A2(n769), .ZN(G153) );
  NOR2_X1 U849 ( .A1(n763), .A2(G868), .ZN(n765) );
  INV_X1 U850 ( .A(G868), .ZN(n766) );
  NOR2_X1 U851 ( .A1(n766), .A2(G301), .ZN(n764) );
  NOR2_X1 U852 ( .A1(n765), .A2(n764), .ZN(G284) );
  NOR2_X1 U853 ( .A1(G286), .A2(n766), .ZN(n768) );
  NOR2_X1 U854 ( .A1(G868), .A2(G299), .ZN(n767) );
  NOR2_X1 U855 ( .A1(n768), .A2(n767), .ZN(G297) );
  NAND2_X1 U856 ( .A1(n769), .A2(G559), .ZN(n770) );
  NAND2_X1 U857 ( .A1(n770), .A2(n1003), .ZN(n771) );
  XNOR2_X1 U858 ( .A(n771), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U859 ( .A1(G868), .A2(n1006), .ZN(n774) );
  NAND2_X1 U860 ( .A1(n1003), .A2(G868), .ZN(n772) );
  NOR2_X1 U861 ( .A1(G559), .A2(n772), .ZN(n773) );
  NOR2_X1 U862 ( .A1(n774), .A2(n773), .ZN(G282) );
  NAND2_X1 U863 ( .A1(G111), .A2(n984), .ZN(n781) );
  NAND2_X1 U864 ( .A1(G135), .A2(n988), .ZN(n776) );
  NAND2_X1 U865 ( .A1(G99), .A2(n989), .ZN(n775) );
  NAND2_X1 U866 ( .A1(n776), .A2(n775), .ZN(n779) );
  NAND2_X1 U867 ( .A1(n985), .A2(G123), .ZN(n777) );
  XOR2_X1 U868 ( .A(KEYINPUT18), .B(n777), .Z(n778) );
  NOR2_X1 U869 ( .A1(n779), .A2(n778), .ZN(n780) );
  NAND2_X1 U870 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U871 ( .A(n782), .B(KEYINPUT79), .ZN(n976) );
  XNOR2_X1 U872 ( .A(n976), .B(G2096), .ZN(n783) );
  INV_X1 U873 ( .A(G2100), .ZN(n948) );
  NAND2_X1 U874 ( .A1(n783), .A2(n948), .ZN(G156) );
  NAND2_X1 U875 ( .A1(n1003), .A2(G559), .ZN(n784) );
  XNOR2_X1 U876 ( .A(n784), .B(n1006), .ZN(n806) );
  NOR2_X1 U877 ( .A1(n806), .A2(G860), .ZN(n795) );
  NAND2_X1 U878 ( .A1(G67), .A2(n785), .ZN(n788) );
  NAND2_X1 U879 ( .A1(G55), .A2(n786), .ZN(n787) );
  NAND2_X1 U880 ( .A1(n788), .A2(n787), .ZN(n794) );
  NAND2_X1 U881 ( .A1(G93), .A2(n789), .ZN(n792) );
  NAND2_X1 U882 ( .A1(G80), .A2(n790), .ZN(n791) );
  NAND2_X1 U883 ( .A1(n792), .A2(n791), .ZN(n793) );
  NOR2_X1 U884 ( .A1(n794), .A2(n793), .ZN(n800) );
  XNOR2_X1 U885 ( .A(n795), .B(n800), .ZN(G145) );
  NOR2_X1 U886 ( .A1(G868), .A2(n800), .ZN(n796) );
  XNOR2_X1 U887 ( .A(n796), .B(KEYINPUT83), .ZN(n809) );
  XNOR2_X1 U888 ( .A(KEYINPUT81), .B(KEYINPUT19), .ZN(n798) );
  XNOR2_X1 U889 ( .A(G288), .B(KEYINPUT82), .ZN(n797) );
  XNOR2_X1 U890 ( .A(n798), .B(n797), .ZN(n799) );
  XNOR2_X1 U891 ( .A(n800), .B(n799), .ZN(n802) );
  XOR2_X1 U892 ( .A(G290), .B(G303), .Z(n801) );
  XNOR2_X1 U893 ( .A(n802), .B(n801), .ZN(n804) );
  XOR2_X1 U894 ( .A(n804), .B(n803), .Z(n805) );
  XNOR2_X1 U895 ( .A(n805), .B(G305), .ZN(n1002) );
  XNOR2_X1 U896 ( .A(n1002), .B(n806), .ZN(n807) );
  NAND2_X1 U897 ( .A1(G868), .A2(n807), .ZN(n808) );
  NAND2_X1 U898 ( .A1(n809), .A2(n808), .ZN(G295) );
  NAND2_X1 U899 ( .A1(G2084), .A2(G2078), .ZN(n810) );
  XOR2_X1 U900 ( .A(KEYINPUT20), .B(n810), .Z(n811) );
  NAND2_X1 U901 ( .A1(G2090), .A2(n811), .ZN(n812) );
  XNOR2_X1 U902 ( .A(KEYINPUT21), .B(n812), .ZN(n813) );
  NAND2_X1 U903 ( .A1(n813), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U904 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U905 ( .A(KEYINPUT73), .B(G132), .ZN(G219) );
  NOR2_X1 U906 ( .A1(G220), .A2(G219), .ZN(n814) );
  XOR2_X1 U907 ( .A(KEYINPUT22), .B(n814), .Z(n815) );
  XNOR2_X1 U908 ( .A(n815), .B(KEYINPUT84), .ZN(n816) );
  NOR2_X1 U909 ( .A1(G218), .A2(n816), .ZN(n817) );
  NAND2_X1 U910 ( .A1(G96), .A2(n817), .ZN(n826) );
  NAND2_X1 U911 ( .A1(n826), .A2(G2106), .ZN(n821) );
  NAND2_X1 U912 ( .A1(G120), .A2(G108), .ZN(n818) );
  NOR2_X1 U913 ( .A1(G237), .A2(n818), .ZN(n819) );
  NAND2_X1 U914 ( .A1(G69), .A2(n819), .ZN(n827) );
  NAND2_X1 U915 ( .A1(n827), .A2(G567), .ZN(n820) );
  NAND2_X1 U916 ( .A1(n821), .A2(n820), .ZN(n972) );
  NAND2_X1 U917 ( .A1(G661), .A2(G483), .ZN(n822) );
  NOR2_X1 U918 ( .A1(n972), .A2(n822), .ZN(n825) );
  NAND2_X1 U919 ( .A1(n825), .A2(G36), .ZN(G176) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n1017), .ZN(G217) );
  AND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n823) );
  NAND2_X1 U922 ( .A1(G661), .A2(n823), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n824) );
  NAND2_X1 U924 ( .A1(n825), .A2(n824), .ZN(G188) );
  NOR2_X1 U925 ( .A1(n827), .A2(n826), .ZN(G325) );
  XOR2_X1 U926 ( .A(KEYINPUT106), .B(G325), .Z(G261) );
  XOR2_X1 U927 ( .A(G108), .B(KEYINPUT116), .Z(G238) );
  NAND2_X1 U929 ( .A1(G124), .A2(n985), .ZN(n828) );
  XNOR2_X1 U930 ( .A(n828), .B(KEYINPUT44), .ZN(n830) );
  NAND2_X1 U931 ( .A1(n989), .A2(G100), .ZN(n829) );
  NAND2_X1 U932 ( .A1(n830), .A2(n829), .ZN(n834) );
  NAND2_X1 U933 ( .A1(G136), .A2(n988), .ZN(n832) );
  NAND2_X1 U934 ( .A1(G112), .A2(n984), .ZN(n831) );
  NAND2_X1 U935 ( .A1(n832), .A2(n831), .ZN(n833) );
  NOR2_X1 U936 ( .A1(n834), .A2(n833), .ZN(G162) );
  XNOR2_X1 U937 ( .A(KEYINPUT56), .B(G16), .ZN(n858) );
  XOR2_X1 U938 ( .A(n1003), .B(n835), .Z(n839) );
  XNOR2_X1 U939 ( .A(G1341), .B(n1006), .ZN(n836) );
  NOR2_X1 U940 ( .A1(n837), .A2(n836), .ZN(n838) );
  NAND2_X1 U941 ( .A1(n839), .A2(n838), .ZN(n846) );
  NAND2_X1 U942 ( .A1(n841), .A2(n840), .ZN(n843) );
  INV_X1 U943 ( .A(G1971), .ZN(n958) );
  NOR2_X1 U944 ( .A1(G166), .A2(n958), .ZN(n842) );
  NOR2_X1 U945 ( .A1(n843), .A2(n842), .ZN(n844) );
  XOR2_X1 U946 ( .A(KEYINPUT122), .B(n844), .Z(n845) );
  NOR2_X1 U947 ( .A1(n846), .A2(n845), .ZN(n856) );
  XOR2_X1 U948 ( .A(G299), .B(G1956), .Z(n848) );
  XOR2_X1 U949 ( .A(G301), .B(G1961), .Z(n847) );
  NAND2_X1 U950 ( .A1(n848), .A2(n847), .ZN(n854) );
  XNOR2_X1 U951 ( .A(G1966), .B(G168), .ZN(n850) );
  NAND2_X1 U952 ( .A1(n850), .A2(n849), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n851), .B(KEYINPUT121), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n852), .B(KEYINPUT57), .ZN(n853) );
  NOR2_X1 U955 ( .A1(n854), .A2(n853), .ZN(n855) );
  NAND2_X1 U956 ( .A1(n856), .A2(n855), .ZN(n857) );
  NAND2_X1 U957 ( .A1(n858), .A2(n857), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n859), .B(KEYINPUT123), .ZN(n885) );
  XNOR2_X1 U959 ( .A(KEYINPUT59), .B(G4), .ZN(n860) );
  XOR2_X1 U960 ( .A(n860), .B(G1348), .Z(n867) );
  XOR2_X1 U961 ( .A(G1341), .B(G19), .Z(n862) );
  XOR2_X1 U962 ( .A(G1956), .B(G20), .Z(n861) );
  NAND2_X1 U963 ( .A1(n862), .A2(n861), .ZN(n864) );
  XNOR2_X1 U964 ( .A(G6), .B(G1981), .ZN(n863) );
  NOR2_X1 U965 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U966 ( .A(KEYINPUT124), .B(n865), .Z(n866) );
  NOR2_X1 U967 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U968 ( .A(KEYINPUT60), .B(n868), .ZN(n870) );
  XOR2_X1 U969 ( .A(G1961), .B(G5), .Z(n869) );
  NAND2_X1 U970 ( .A1(n870), .A2(n869), .ZN(n873) );
  XOR2_X1 U971 ( .A(G21), .B(G1966), .Z(n871) );
  XNOR2_X1 U972 ( .A(KEYINPUT125), .B(n871), .ZN(n872) );
  NOR2_X1 U973 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U974 ( .A(KEYINPUT126), .B(n874), .ZN(n881) );
  XOR2_X1 U975 ( .A(G1976), .B(G23), .Z(n876) );
  XNOR2_X1 U976 ( .A(n958), .B(G22), .ZN(n875) );
  NAND2_X1 U977 ( .A1(n876), .A2(n875), .ZN(n878) );
  XNOR2_X1 U978 ( .A(G24), .B(G1986), .ZN(n877) );
  NOR2_X1 U979 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U980 ( .A(KEYINPUT58), .B(n879), .ZN(n880) );
  NAND2_X1 U981 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U982 ( .A(KEYINPUT61), .B(n882), .ZN(n883) );
  NOR2_X1 U983 ( .A1(n883), .A2(G16), .ZN(n884) );
  NOR2_X1 U984 ( .A1(n885), .A2(n884), .ZN(n921) );
  NOR2_X1 U985 ( .A1(n887), .A2(n886), .ZN(n914) );
  XOR2_X1 U986 ( .A(G2090), .B(G162), .Z(n888) );
  NOR2_X1 U987 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U988 ( .A(KEYINPUT51), .B(n890), .Z(n893) );
  NOR2_X1 U989 ( .A1(n891), .A2(n976), .ZN(n892) );
  NAND2_X1 U990 ( .A1(n893), .A2(n892), .ZN(n896) );
  XNOR2_X1 U991 ( .A(G2084), .B(G160), .ZN(n894) );
  XNOR2_X1 U992 ( .A(KEYINPUT117), .B(n894), .ZN(n895) );
  NOR2_X1 U993 ( .A1(n896), .A2(n895), .ZN(n898) );
  NAND2_X1 U994 ( .A1(n898), .A2(n897), .ZN(n912) );
  NAND2_X1 U995 ( .A1(n989), .A2(G103), .ZN(n899) );
  XNOR2_X1 U996 ( .A(n899), .B(KEYINPUT110), .ZN(n901) );
  NAND2_X1 U997 ( .A1(G139), .A2(n988), .ZN(n900) );
  NAND2_X1 U998 ( .A1(n901), .A2(n900), .ZN(n902) );
  XOR2_X1 U999 ( .A(KEYINPUT111), .B(n902), .Z(n907) );
  NAND2_X1 U1000 ( .A1(G115), .A2(n984), .ZN(n904) );
  NAND2_X1 U1001 ( .A1(G127), .A2(n985), .ZN(n903) );
  NAND2_X1 U1002 ( .A1(n904), .A2(n903), .ZN(n905) );
  XOR2_X1 U1003 ( .A(KEYINPUT47), .B(n905), .Z(n906) );
  NOR2_X1 U1004 ( .A1(n907), .A2(n906), .ZN(n996) );
  XOR2_X1 U1005 ( .A(G2072), .B(n996), .Z(n909) );
  XOR2_X1 U1006 ( .A(G164), .B(G2078), .Z(n908) );
  NOR2_X1 U1007 ( .A1(n909), .A2(n908), .ZN(n910) );
  XOR2_X1 U1008 ( .A(KEYINPUT50), .B(n910), .Z(n911) );
  NOR2_X1 U1009 ( .A1(n912), .A2(n911), .ZN(n913) );
  NAND2_X1 U1010 ( .A1(n914), .A2(n913), .ZN(n915) );
  NOR2_X1 U1011 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1012 ( .A(KEYINPUT52), .B(n917), .ZN(n918) );
  INV_X1 U1013 ( .A(KEYINPUT55), .ZN(n940) );
  NAND2_X1 U1014 ( .A1(n918), .A2(n940), .ZN(n919) );
  NAND2_X1 U1015 ( .A1(n919), .A2(G29), .ZN(n920) );
  NAND2_X1 U1016 ( .A1(n921), .A2(n920), .ZN(n946) );
  XOR2_X1 U1017 ( .A(G29), .B(KEYINPUT120), .Z(n943) );
  XOR2_X1 U1018 ( .A(G32), .B(G1996), .Z(n928) );
  XOR2_X1 U1019 ( .A(G25), .B(G1991), .Z(n922) );
  NAND2_X1 U1020 ( .A1(n922), .A2(G28), .ZN(n926) );
  XNOR2_X1 U1021 ( .A(G27), .B(n923), .ZN(n924) );
  XNOR2_X1 U1022 ( .A(KEYINPUT119), .B(n924), .ZN(n925) );
  NOR2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1024 ( .A1(n928), .A2(n927), .ZN(n933) );
  XNOR2_X1 U1025 ( .A(G2067), .B(G26), .ZN(n930) );
  XNOR2_X1 U1026 ( .A(G33), .B(G2072), .ZN(n929) );
  NOR2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1028 ( .A(KEYINPUT118), .B(n931), .Z(n932) );
  NOR2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1030 ( .A(KEYINPUT53), .B(n934), .Z(n937) );
  XOR2_X1 U1031 ( .A(G34), .B(KEYINPUT54), .Z(n935) );
  XNOR2_X1 U1032 ( .A(G2084), .B(n935), .ZN(n936) );
  NAND2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n939) );
  XNOR2_X1 U1034 ( .A(G35), .B(G2090), .ZN(n938) );
  NOR2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n941) );
  XOR2_X1 U1036 ( .A(n941), .B(n940), .Z(n942) );
  NAND2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1038 ( .A1(G11), .A2(n944), .ZN(n945) );
  NOR2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(n947), .B(KEYINPUT62), .ZN(G311) );
  XNOR2_X1 U1041 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1042 ( .A(G120), .ZN(G236) );
  XNOR2_X1 U1043 ( .A(G2678), .B(n948), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(G2067), .B(G2084), .ZN(n949) );
  XNOR2_X1 U1045 ( .A(n950), .B(n949), .ZN(n951) );
  XOR2_X1 U1046 ( .A(n951), .B(KEYINPUT107), .Z(n953) );
  XNOR2_X1 U1047 ( .A(G2090), .B(KEYINPUT42), .ZN(n952) );
  XNOR2_X1 U1048 ( .A(n953), .B(n952), .ZN(n957) );
  XOR2_X1 U1049 ( .A(G2096), .B(KEYINPUT43), .Z(n955) );
  XNOR2_X1 U1050 ( .A(G2078), .B(G2072), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(n955), .B(n954), .ZN(n956) );
  XOR2_X1 U1052 ( .A(n957), .B(n956), .Z(G227) );
  XOR2_X1 U1053 ( .A(n958), .B(G1976), .Z(n971) );
  XOR2_X1 U1054 ( .A(G2474), .B(KEYINPUT41), .Z(n961) );
  INV_X1 U1055 ( .A(G1996), .ZN(n959) );
  XOR2_X1 U1056 ( .A(n959), .B(G1986), .Z(n960) );
  XNOR2_X1 U1057 ( .A(n961), .B(n960), .ZN(n967) );
  XNOR2_X1 U1058 ( .A(G1981), .B(n962), .ZN(n965) );
  XOR2_X1 U1059 ( .A(G1966), .B(n963), .Z(n964) );
  XNOR2_X1 U1060 ( .A(n965), .B(n964), .ZN(n966) );
  XOR2_X1 U1061 ( .A(n967), .B(n966), .Z(n969) );
  XNOR2_X1 U1062 ( .A(G1991), .B(KEYINPUT108), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(n969), .B(n968), .ZN(n970) );
  XNOR2_X1 U1064 ( .A(n971), .B(n970), .ZN(G229) );
  INV_X1 U1065 ( .A(n972), .ZN(G319) );
  XOR2_X1 U1066 ( .A(KEYINPUT109), .B(KEYINPUT46), .Z(n974) );
  XNOR2_X1 U1067 ( .A(KEYINPUT112), .B(KEYINPUT48), .ZN(n973) );
  XNOR2_X1 U1068 ( .A(n974), .B(n973), .ZN(n975) );
  XNOR2_X1 U1069 ( .A(n976), .B(n975), .ZN(n979) );
  XNOR2_X1 U1070 ( .A(n977), .B(G162), .ZN(n978) );
  XNOR2_X1 U1071 ( .A(n979), .B(n978), .ZN(n983) );
  XNOR2_X1 U1072 ( .A(G164), .B(G160), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(n981), .B(n980), .ZN(n982) );
  XOR2_X1 U1074 ( .A(n983), .B(n982), .Z(n998) );
  NAND2_X1 U1075 ( .A1(G118), .A2(n984), .ZN(n987) );
  NAND2_X1 U1076 ( .A1(G130), .A2(n985), .ZN(n986) );
  NAND2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n994) );
  NAND2_X1 U1078 ( .A1(G142), .A2(n988), .ZN(n991) );
  NAND2_X1 U1079 ( .A1(G106), .A2(n989), .ZN(n990) );
  NAND2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  XOR2_X1 U1081 ( .A(KEYINPUT45), .B(n992), .Z(n993) );
  NOR2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1083 ( .A(n996), .B(n995), .ZN(n997) );
  XNOR2_X1 U1084 ( .A(n998), .B(n997), .ZN(n1000) );
  XNOR2_X1 U1085 ( .A(n1000), .B(n999), .ZN(n1001) );
  NOR2_X1 U1086 ( .A1(G37), .A2(n1001), .ZN(G395) );
  XOR2_X1 U1087 ( .A(KEYINPUT113), .B(n1002), .Z(n1005) );
  XOR2_X1 U1088 ( .A(n1003), .B(G286), .Z(n1004) );
  XNOR2_X1 U1089 ( .A(n1005), .B(n1004), .ZN(n1008) );
  XOR2_X1 U1090 ( .A(n1006), .B(G301), .Z(n1007) );
  XNOR2_X1 U1091 ( .A(n1008), .B(n1007), .ZN(n1009) );
  NOR2_X1 U1092 ( .A1(G37), .A2(n1009), .ZN(G397) );
  NOR2_X1 U1093 ( .A1(G227), .A2(G229), .ZN(n1010) );
  XOR2_X1 U1094 ( .A(KEYINPUT49), .B(n1010), .Z(n1011) );
  XNOR2_X1 U1095 ( .A(KEYINPUT114), .B(n1011), .ZN(n1016) );
  NOR2_X1 U1096 ( .A1(G395), .A2(G397), .ZN(n1012) );
  XOR2_X1 U1097 ( .A(KEYINPUT115), .B(n1012), .Z(n1013) );
  NAND2_X1 U1098 ( .A1(G319), .A2(n1013), .ZN(n1014) );
  NOR2_X1 U1099 ( .A1(G401), .A2(n1014), .ZN(n1015) );
  NAND2_X1 U1100 ( .A1(n1016), .A2(n1015), .ZN(G225) );
  INV_X1 U1101 ( .A(G225), .ZN(G308) );
  INV_X1 U1102 ( .A(G96), .ZN(G221) );
  INV_X1 U1103 ( .A(G69), .ZN(G235) );
  INV_X1 U1104 ( .A(n1017), .ZN(G223) );
endmodule

