//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 0 0 0 1 1 1 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 1 0 1 1 1 1 1 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1256, new_n1257, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(KEYINPUT64), .ZN(new_n205));
  INV_X1    g0005(.A(G77), .ZN(new_n206));
  NOR2_X1   g0006(.A1(G58), .A2(G68), .ZN(new_n207));
  INV_X1    g0007(.A(KEYINPUT64), .ZN(new_n208));
  NAND3_X1  g0008(.A1(new_n207), .A2(new_n208), .A3(new_n201), .ZN(new_n209));
  AND3_X1   g0009(.A1(new_n205), .A2(new_n206), .A3(new_n209), .ZN(G353));
  OAI21_X1  g0010(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0011(.A(G1), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT0), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n213), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(new_n207), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(G50), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  INV_X1    g0024(.A(G238), .ZN(new_n225));
  INV_X1    g0025(.A(G87), .ZN(new_n226));
  INV_X1    g0026(.A(G250), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n224), .B1(new_n203), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  INV_X1    g0030(.A(G97), .ZN(new_n231));
  INV_X1    g0031(.A(G257), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n229), .B1(new_n202), .B2(new_n230), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n215), .B1(new_n228), .B2(new_n233), .ZN(new_n234));
  OAI221_X1 g0034(.A(new_n218), .B1(new_n221), .B2(new_n223), .C1(KEYINPUT1), .C2(new_n234), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n235), .B1(KEYINPUT1), .B2(new_n234), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n201), .A2(G68), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n203), .A2(G50), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n247), .B(new_n252), .Z(G351));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G1), .A3(G13), .ZN(new_n255));
  INV_X1    g0055(.A(G41), .ZN(new_n256));
  OAI211_X1 g0056(.A(new_n212), .B(G45), .C1(new_n256), .C2(KEYINPUT5), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT5), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G41), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n255), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT79), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n261), .B1(new_n258), .B2(G41), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n256), .A2(KEYINPUT79), .A3(KEYINPUT5), .ZN(new_n263));
  INV_X1    g0063(.A(G45), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(G1), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n258), .A2(G41), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n262), .A2(new_n263), .A3(new_n265), .A4(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n255), .A2(G274), .ZN(new_n268));
  OAI22_X1  g0068(.A1(new_n260), .A2(new_n232), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  AND2_X1   g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NOR2_X1   g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  OAI211_X1 g0073(.A(G244), .B(new_n271), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT78), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT4), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G283), .ZN(new_n279));
  OAI211_X1 g0079(.A(G250), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n279), .B(new_n280), .C1(new_n274), .C2(new_n276), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n275), .B1(new_n274), .B2(new_n276), .ZN(new_n282));
  NOR3_X1   g0082(.A1(new_n278), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n270), .B1(new_n283), .B2(new_n255), .ZN(new_n284));
  INV_X1    g0084(.A(G169), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT3), .ZN(new_n287));
  INV_X1    g0087(.A(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n289), .A2(new_n213), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT7), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n289), .A2(KEYINPUT7), .A3(new_n213), .A4(new_n290), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n293), .A2(KEYINPUT75), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G107), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT67), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT67), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G107), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  OR2_X1    g0100(.A1(new_n294), .A2(KEYINPUT75), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n295), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n296), .A2(KEYINPUT6), .A3(G97), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n231), .A2(new_n296), .ZN(new_n304));
  NOR2_X1   g0104(.A1(G97), .A2(G107), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n303), .B1(new_n306), .B2(KEYINPUT6), .ZN(new_n307));
  NOR2_X1   g0107(.A1(G20), .A2(G33), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n307), .A2(G20), .B1(G77), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n302), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n219), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n212), .A2(G13), .A3(G20), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n231), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n314), .A2(new_n219), .A3(new_n311), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n317), .B1(new_n212), .B2(G33), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n316), .B1(new_n319), .B2(new_n231), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n313), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n269), .A2(KEYINPUT80), .ZN(new_n323));
  INV_X1    g0123(.A(G274), .ZN(new_n324));
  INV_X1    g0124(.A(new_n219), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n324), .B1(new_n325), .B2(new_n254), .ZN(new_n326));
  INV_X1    g0126(.A(new_n257), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n326), .A2(new_n327), .A3(new_n262), .A4(new_n263), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT80), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n328), .B(new_n329), .C1(new_n232), .C2(new_n260), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n323), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n274), .A2(new_n276), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT78), .ZN(new_n333));
  OR2_X1    g0133(.A1(new_n274), .A2(new_n276), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n280), .A2(new_n279), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n333), .A2(new_n334), .A3(new_n277), .A4(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n255), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G179), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n331), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  AND3_X1   g0140(.A1(new_n286), .A2(new_n322), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n320), .B1(new_n310), .B2(new_n312), .ZN(new_n342));
  OAI211_X1 g0142(.A(G190), .B(new_n270), .C1(new_n283), .C2(new_n255), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G200), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n345), .B1(new_n331), .B2(new_n338), .ZN(new_n346));
  OAI21_X1  g0146(.A(KEYINPUT81), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n283), .A2(new_n255), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n323), .A2(new_n330), .ZN(new_n349));
  OAI21_X1  g0149(.A(G200), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT81), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n350), .A2(new_n351), .A3(new_n342), .A4(new_n343), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n341), .B1(new_n347), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n315), .A2(new_n203), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n354), .B(KEYINPUT12), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n308), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n213), .A2(G33), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n356), .B1(new_n206), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n358), .A2(KEYINPUT11), .A3(new_n312), .ZN(new_n359));
  INV_X1    g0159(.A(new_n317), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n212), .A2(G20), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n360), .A2(G68), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n355), .A2(new_n359), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT11), .B1(new_n358), .B2(new_n312), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(G1), .B1(new_n256), .B2(new_n264), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n367), .A2(new_n255), .A3(G274), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n212), .B1(G41), .B2(G45), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n255), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n369), .B1(G238), .B2(new_n372), .ZN(new_n373));
  OAI211_X1 g0173(.A(G232), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT72), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n289), .A2(new_n290), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT72), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n376), .A2(new_n377), .A3(G232), .A4(G1698), .ZN(new_n378));
  NAND2_X1  g0178(.A1(G33), .A2(G97), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n376), .A2(G226), .A3(new_n271), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n375), .A2(new_n378), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n381), .A2(KEYINPUT73), .A3(new_n337), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT73), .B1(new_n381), .B2(new_n337), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n373), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT13), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT13), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n386), .B(new_n373), .C1(new_n382), .C2(new_n383), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT14), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n389), .A3(G169), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n385), .A2(G179), .A3(new_n387), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n389), .B1(new_n388), .B2(G169), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n366), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI211_X1 g0194(.A(G222), .B(new_n271), .C1(new_n272), .C2(new_n273), .ZN(new_n395));
  OAI211_X1 g0195(.A(G223), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n395), .B(new_n396), .C1(new_n206), .C2(new_n376), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n337), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n255), .A2(G226), .A3(new_n370), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n368), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT65), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n368), .A2(new_n399), .A3(KEYINPUT65), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n398), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(G200), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n398), .A2(G190), .A3(new_n402), .A4(new_n403), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT9), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n213), .B1(new_n205), .B2(new_n209), .ZN(new_n408));
  XNOR2_X1  g0208(.A(KEYINPUT8), .B(G58), .ZN(new_n409));
  INV_X1    g0209(.A(G150), .ZN(new_n410));
  INV_X1    g0210(.A(new_n308), .ZN(new_n411));
  OAI22_X1  g0211(.A1(new_n409), .A2(new_n357), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n312), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n201), .B1(new_n212), .B2(G20), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n360), .A2(new_n414), .B1(new_n201), .B2(new_n315), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n407), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  AND3_X1   g0216(.A1(new_n413), .A2(new_n407), .A3(new_n415), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n405), .B(new_n406), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT10), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT71), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT71), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n418), .A2(new_n421), .A3(KEYINPUT10), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n405), .A2(new_n406), .ZN(new_n423));
  INV_X1    g0223(.A(new_n416), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT70), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n413), .A2(new_n407), .A3(new_n415), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT10), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT70), .B1(new_n417), .B2(new_n416), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n423), .A2(new_n427), .A3(new_n428), .A4(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n420), .A2(new_n422), .A3(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n404), .A2(G179), .ZN(new_n432));
  XNOR2_X1  g0232(.A(new_n432), .B(KEYINPUT66), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n404), .A2(new_n285), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n413), .A2(new_n415), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT68), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n271), .B1(new_n289), .B2(new_n290), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n272), .A2(new_n273), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n438), .A2(G238), .B1(new_n300), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n376), .A2(G232), .A3(new_n271), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n337), .ZN(new_n443));
  INV_X1    g0243(.A(G244), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n368), .B1(new_n444), .B2(new_n371), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n437), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n255), .B1(new_n440), .B2(new_n441), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n448), .A2(KEYINPUT68), .A3(new_n445), .ZN(new_n449));
  OAI21_X1  g0249(.A(G190), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n409), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n451), .A2(new_n308), .B1(G20), .B2(G77), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT69), .ZN(new_n453));
  XNOR2_X1  g0253(.A(KEYINPUT15), .B(G87), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n453), .B1(new_n454), .B2(new_n357), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n452), .A2(KEYINPUT69), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n312), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n206), .B1(new_n212), .B2(G20), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n360), .A2(new_n458), .B1(new_n206), .B2(new_n315), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n443), .A2(new_n437), .A3(new_n446), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT68), .B1(new_n448), .B2(new_n445), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n460), .A2(G200), .A3(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n450), .A2(new_n457), .A3(new_n459), .A4(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n339), .B1(new_n447), .B2(new_n449), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n457), .A2(new_n459), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n460), .A2(new_n285), .A3(new_n461), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  AND3_X1   g0268(.A1(new_n431), .A2(new_n436), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n388), .A2(G200), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n385), .A2(G190), .A3(new_n387), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n470), .A2(new_n365), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT17), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n451), .A2(new_n361), .ZN(new_n474));
  OAI22_X1  g0274(.A1(new_n474), .A2(new_n317), .B1(new_n314), .B2(new_n451), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT76), .B1(new_n371), .B2(new_n230), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT76), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n255), .A2(new_n370), .A3(new_n478), .A4(G232), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  OR2_X1    g0280(.A1(G223), .A2(G1698), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(G226), .B2(new_n271), .ZN(new_n482));
  OAI22_X1  g0282(.A1(new_n482), .A2(new_n439), .B1(new_n288), .B2(new_n226), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n337), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n480), .A2(new_n484), .A3(new_n368), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n345), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(G190), .B2(new_n485), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT74), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n202), .A2(new_n203), .ZN(new_n489));
  OAI21_X1  g0289(.A(G20), .B1(new_n489), .B2(new_n207), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n308), .A2(G159), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n293), .A2(new_n294), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n492), .B1(new_n493), .B2(G68), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n488), .B1(new_n494), .B2(KEYINPUT16), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n203), .B1(new_n293), .B2(new_n294), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT16), .ZN(new_n497));
  NOR4_X1   g0297(.A1(new_n496), .A2(KEYINPUT74), .A3(new_n492), .A4(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n312), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n295), .A2(G68), .A3(new_n301), .ZN(new_n500));
  INV_X1    g0300(.A(new_n492), .ZN(new_n501));
  AOI21_X1  g0301(.A(KEYINPUT16), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n476), .B(new_n487), .C1(new_n499), .C2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n473), .B1(new_n503), .B2(KEYINPUT77), .ZN(new_n504));
  INV_X1    g0304(.A(new_n312), .ZN(new_n505));
  AOI21_X1  g0305(.A(KEYINPUT7), .B1(new_n439), .B2(new_n213), .ZN(new_n506));
  INV_X1    g0306(.A(new_n294), .ZN(new_n507));
  OAI21_X1  g0307(.A(G68), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n508), .A2(KEYINPUT16), .A3(new_n501), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT74), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n494), .A2(new_n488), .A3(KEYINPUT16), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n505), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n502), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n475), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT77), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT17), .A4(new_n487), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n485), .A2(new_n339), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n369), .B1(new_n483), .B2(new_n337), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n285), .B1(new_n518), .B2(new_n480), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(KEYINPUT18), .B1(new_n514), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n476), .B1(new_n499), .B2(new_n502), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT18), .ZN(new_n523));
  INV_X1    g0323(.A(new_n520), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AND4_X1   g0325(.A1(new_n504), .A2(new_n516), .A3(new_n521), .A4(new_n525), .ZN(new_n526));
  AND4_X1   g0326(.A1(new_n394), .A2(new_n469), .A3(new_n472), .A4(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(G116), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n311), .A2(new_n219), .B1(G20), .B2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n279), .B(new_n213), .C1(G33), .C2(new_n231), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT20), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n529), .A2(KEYINPUT20), .A3(new_n530), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n318), .A2(G116), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n315), .A2(new_n528), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  OAI211_X1 g0339(.A(G270), .B(new_n255), .C1(new_n257), .C2(new_n259), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n268), .B2(new_n267), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(G264), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n543));
  OAI211_X1 g0343(.A(G257), .B(new_n271), .C1(new_n272), .C2(new_n273), .ZN(new_n544));
  INV_X1    g0344(.A(G303), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n543), .B(new_n544), .C1(new_n545), .C2(new_n376), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n337), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n542), .A2(new_n547), .A3(G190), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n541), .B1(new_n337), .B2(new_n546), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n539), .B(new_n548), .C1(new_n345), .C2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n542), .A2(new_n547), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n538), .A2(new_n551), .A3(G169), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT21), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n538), .A2(new_n549), .A3(G179), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n538), .A2(new_n551), .A3(KEYINPUT21), .A4(G169), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n550), .A2(new_n554), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT86), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n556), .A2(new_n555), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n560), .A2(KEYINPUT86), .A3(new_n554), .A4(new_n550), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n227), .A2(new_n271), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n232), .A2(G1698), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n563), .B(new_n564), .C1(new_n272), .C2(new_n273), .ZN(new_n565));
  NAND2_X1  g0365(.A1(G33), .A2(G294), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(KEYINPUT89), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(KEYINPUT89), .B1(new_n565), .B2(new_n566), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n337), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(G264), .B(new_n255), .C1(new_n257), .C2(new_n259), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n328), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G179), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n565), .A2(new_n566), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT89), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n255), .B1(new_n579), .B2(new_n567), .ZN(new_n580));
  OAI21_X1  g0380(.A(KEYINPUT90), .B1(new_n580), .B2(new_n572), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT90), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n570), .A2(new_n573), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n581), .A2(new_n583), .A3(G169), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n576), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n213), .B(G87), .C1(new_n272), .C2(new_n273), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT22), .ZN(new_n587));
  XNOR2_X1  g0387(.A(new_n586), .B(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT23), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n589), .A2(new_n296), .A3(G20), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT87), .ZN(new_n591));
  XNOR2_X1  g0391(.A(new_n590), .B(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n213), .A2(G33), .A3(G116), .ZN(new_n593));
  OAI21_X1  g0393(.A(KEYINPUT23), .B1(new_n300), .B2(new_n213), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(KEYINPUT24), .B1(new_n588), .B2(new_n595), .ZN(new_n596));
  XNOR2_X1  g0396(.A(new_n586), .B(KEYINPUT22), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n594), .A2(new_n593), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT24), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .A4(new_n592), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n312), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT25), .ZN(new_n603));
  AOI211_X1 g0403(.A(G107), .B(new_n314), .C1(KEYINPUT88), .C2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n603), .A2(KEYINPUT88), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n604), .A2(new_n605), .ZN(new_n607));
  OAI22_X1  g0407(.A1(new_n606), .A2(new_n607), .B1(new_n296), .B2(new_n319), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n602), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n585), .A2(new_n610), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n213), .B(G68), .C1(new_n272), .C2(new_n273), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT19), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT83), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT83), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(KEYINPUT19), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n357), .A2(new_n231), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n612), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n379), .B1(new_n614), .B2(new_n616), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n226), .A2(new_n231), .ZN(new_n621));
  OAI22_X1  g0421(.A1(new_n620), .A2(G20), .B1(new_n300), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT84), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n619), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI221_X1 g0424(.A(KEYINPUT84), .B1(new_n300), .B2(new_n621), .C1(new_n620), .C2(G20), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n505), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n225), .A2(new_n271), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n444), .A2(G1698), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n627), .B(new_n628), .C1(new_n272), .C2(new_n273), .ZN(new_n629));
  NAND2_X1  g0429(.A1(G33), .A2(G116), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n255), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(KEYINPUT82), .A2(G250), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n264), .B2(G1), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n255), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n212), .A2(new_n324), .A3(G45), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n227), .A2(KEYINPUT82), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n631), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n639), .A2(new_n345), .ZN(new_n640));
  INV_X1    g0440(.A(new_n454), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n641), .A2(new_n314), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n319), .A2(new_n226), .ZN(new_n643));
  NOR4_X1   g0443(.A1(new_n626), .A2(new_n640), .A3(new_n642), .A4(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n639), .A2(G190), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT85), .ZN(new_n646));
  XNOR2_X1  g0446(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n622), .A2(new_n623), .ZN(new_n648));
  INV_X1    g0448(.A(new_n619), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(new_n625), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n642), .B1(new_n650), .B2(new_n312), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n318), .A2(new_n641), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n639), .A2(G169), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n654), .B1(new_n339), .B2(new_n639), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n644), .A2(new_n647), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n608), .B1(new_n601), .B2(new_n312), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n575), .A2(G200), .ZN(new_n658));
  AOI21_X1  g0458(.A(G190), .B1(new_n581), .B2(new_n583), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n611), .A2(new_n656), .A3(new_n660), .ZN(new_n661));
  AND4_X1   g0461(.A1(new_n353), .A2(new_n527), .A3(new_n562), .A4(new_n661), .ZN(G372));
  INV_X1    g0462(.A(new_n436), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT94), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n514), .A2(KEYINPUT18), .A3(new_n520), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n523), .B1(new_n522), .B2(new_n524), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n521), .A2(KEYINPUT94), .A3(new_n525), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n388), .A2(G169), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(KEYINPUT14), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n671), .A2(new_n391), .A3(new_n390), .ZN(new_n672));
  INV_X1    g0472(.A(new_n467), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n672), .A2(new_n366), .B1(new_n472), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n504), .A2(new_n516), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n669), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n663), .B1(new_n676), .B2(new_n431), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n347), .A2(new_n352), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n286), .A2(new_n322), .A3(new_n340), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(new_n680), .A3(new_n660), .ZN(new_n681));
  INV_X1    g0481(.A(new_n640), .ZN(new_n682));
  INV_X1    g0482(.A(new_n643), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n651), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT91), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n651), .A2(KEYINPUT91), .A3(new_n682), .A4(new_n683), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(new_n647), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n653), .A2(new_n655), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(KEYINPUT92), .B1(new_n681), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n645), .B(KEYINPUT85), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n692), .B1(new_n644), .B2(KEYINPUT91), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n693), .A2(new_n686), .B1(new_n653), .B2(new_n655), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT92), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n353), .A2(new_n694), .A3(new_n695), .A4(new_n660), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n560), .A2(new_n554), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT93), .ZN(new_n698));
  AND3_X1   g0498(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT93), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n611), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n691), .A2(new_n696), .A3(new_n703), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n690), .A2(KEYINPUT26), .A3(new_n680), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n689), .B1(new_n692), .B2(new_n684), .ZN(new_n706));
  OAI21_X1  g0506(.A(KEYINPUT26), .B1(new_n706), .B2(new_n680), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n689), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n704), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n678), .B1(new_n527), .B2(new_n710), .ZN(new_n711));
  XOR2_X1   g0511(.A(new_n711), .B(KEYINPUT95), .Z(G369));
  INV_X1    g0512(.A(G13), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n713), .A2(G1), .A3(G20), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT96), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT27), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G213), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n715), .A2(new_n716), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(G343), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n562), .B1(new_n539), .B2(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n698), .A2(new_n701), .A3(new_n538), .A4(new_n723), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G330), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n611), .A2(new_n660), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(new_n657), .B2(new_n724), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n657), .B1(new_n584), .B2(new_n576), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(new_n723), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  OR3_X1    g0534(.A1(new_n728), .A2(new_n734), .A3(KEYINPUT97), .ZN(new_n735));
  OAI21_X1  g0535(.A(KEYINPUT97), .B1(new_n728), .B2(new_n734), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n699), .A2(new_n723), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n729), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n739), .B1(new_n611), .B2(new_n723), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n737), .A2(new_n740), .ZN(G399));
  INV_X1    g0541(.A(new_n216), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G41), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n300), .A2(G116), .A3(new_n621), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n744), .A2(G1), .A3(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(new_n223), .B2(new_n744), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT28), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT29), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n688), .A2(KEYINPUT26), .A3(new_n341), .A4(new_n689), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT26), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(new_n706), .B2(new_n680), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n688), .B1(new_n731), .B2(new_n697), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n753), .B(new_n689), .C1(new_n681), .C2(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n749), .B1(new_n755), .B2(new_n724), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n723), .B1(new_n704), .B2(new_n709), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n756), .B1(new_n757), .B2(new_n749), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n661), .A2(new_n562), .A3(new_n353), .A4(new_n724), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT30), .ZN(new_n761));
  INV_X1    g0561(.A(new_n571), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n631), .A2(new_n762), .A3(new_n638), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n549), .A2(new_n570), .A3(new_n763), .A4(G179), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n761), .B1(new_n764), .B2(new_n284), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n551), .A2(new_n339), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n634), .A2(new_n637), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n629), .A2(new_n630), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n767), .B(new_n571), .C1(new_n768), .C2(new_n255), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n580), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n269), .B1(new_n336), .B2(new_n337), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n766), .A2(new_n770), .A3(new_n771), .A4(KEYINPUT30), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n339), .B1(new_n631), .B2(new_n638), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n773), .B1(new_n542), .B2(new_n547), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n574), .B(new_n774), .C1(new_n348), .C2(new_n349), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n765), .A2(new_n772), .A3(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT98), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n765), .A2(new_n775), .A3(new_n772), .A4(KEYINPUT98), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n778), .A2(new_n723), .A3(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT31), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n776), .A2(KEYINPUT31), .A3(new_n723), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n760), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G330), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n759), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n748), .B1(new_n787), .B2(G1), .ZN(G364));
  NOR2_X1   g0588(.A1(new_n713), .A2(G20), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n212), .B1(new_n789), .B2(G45), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n743), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n742), .A2(new_n439), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n794), .A2(G355), .B1(new_n528), .B2(new_n742), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n742), .A2(new_n376), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(G45), .B2(new_n223), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n252), .A2(new_n264), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n795), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G13), .A2(G33), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(G20), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n219), .B1(G20), .B2(new_n285), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n793), .B1(new_n799), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n803), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n213), .A2(G190), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT99), .ZN(new_n808));
  NOR3_X1   g0608(.A1(new_n808), .A2(G179), .A3(G200), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G159), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT32), .Z(new_n811));
  NAND3_X1  g0611(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(G190), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n813), .A2(KEYINPUT101), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n813), .A2(KEYINPUT101), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(G68), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n339), .A2(G200), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n807), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n376), .B1(new_n820), .B2(new_n206), .ZN(new_n821));
  INV_X1    g0621(.A(G190), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n812), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(G179), .A2(G200), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n213), .B1(new_n825), .B2(G190), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n824), .A2(new_n201), .B1(new_n826), .B2(new_n231), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n213), .A2(new_n822), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n819), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n821), .B(new_n827), .C1(G58), .C2(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n828), .A2(new_n339), .A3(G200), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n832), .A2(KEYINPUT100), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(KEYINPUT100), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NOR3_X1   g0636(.A1(new_n808), .A2(G179), .A3(new_n345), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n836), .A2(G87), .B1(new_n837), .B2(G107), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n811), .A2(new_n818), .A3(new_n831), .A4(new_n838), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n836), .A2(G303), .B1(new_n837), .B2(G283), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n809), .A2(G329), .ZN(new_n841));
  XNOR2_X1  g0641(.A(KEYINPUT33), .B(G317), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n817), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(G322), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n439), .B1(new_n829), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(G326), .ZN(new_n846));
  INV_X1    g0646(.A(G294), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n824), .A2(new_n846), .B1(new_n826), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n820), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n845), .B(new_n848), .C1(G311), .C2(new_n849), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n840), .A2(new_n841), .A3(new_n843), .A4(new_n850), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n839), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n802), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n805), .B1(new_n806), .B2(new_n852), .C1(new_n727), .C2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n728), .A2(new_n793), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n727), .A2(G330), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(G396));
  NAND2_X1  g0657(.A1(new_n468), .A2(new_n724), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(new_n704), .B2(new_n709), .ZN(new_n859));
  INV_X1    g0659(.A(new_n757), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n723), .A2(new_n465), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n463), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n467), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n673), .A2(new_n724), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n859), .B1(new_n860), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n786), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT103), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n868), .B(new_n793), .C1(new_n786), .C2(new_n866), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n803), .A2(new_n800), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n793), .B1(new_n206), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n809), .ZN(new_n872));
  INV_X1    g0672(.A(G132), .ZN(new_n873));
  OAI22_X1  g0673(.A1(new_n872), .A2(new_n873), .B1(new_n201), .B2(new_n835), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n837), .A2(G68), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n875), .B(new_n376), .C1(new_n202), .C2(new_n826), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT34), .ZN(new_n877));
  AOI22_X1  g0677(.A1(G143), .A2(new_n830), .B1(new_n849), .B2(G159), .ZN(new_n878));
  INV_X1    g0678(.A(G137), .ZN(new_n879));
  OAI221_X1 g0679(.A(new_n878), .B1(new_n879), .B2(new_n824), .C1(new_n410), .C2(new_n816), .ZN(new_n880));
  AOI211_X1 g0680(.A(new_n874), .B(new_n876), .C1(new_n877), .C2(new_n880), .ZN(new_n881));
  OR2_X1    g0681(.A1(new_n880), .A2(new_n877), .ZN(new_n882));
  AOI22_X1  g0682(.A1(G294), .A2(new_n830), .B1(new_n849), .B2(G116), .ZN(new_n883));
  OAI221_X1 g0683(.A(new_n883), .B1(new_n231), .B2(new_n826), .C1(new_n545), .C2(new_n824), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n837), .A2(G87), .ZN(new_n885));
  INV_X1    g0685(.A(G311), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n885), .B1(new_n872), .B2(new_n886), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n884), .B(new_n887), .C1(G283), .C2(new_n817), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n439), .B1(new_n835), .B2(new_n296), .ZN(new_n889));
  XOR2_X1   g0689(.A(new_n889), .B(KEYINPUT102), .Z(new_n890));
  AOI22_X1  g0690(.A1(new_n881), .A2(new_n882), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n865), .ZN(new_n892));
  OAI221_X1 g0692(.A(new_n871), .B1(new_n806), .B2(new_n891), .C1(new_n892), .C2(new_n801), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n869), .A2(new_n893), .ZN(G384));
  AND4_X1   g0694(.A1(KEYINPUT31), .A2(new_n778), .A3(new_n723), .A4(new_n779), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n724), .B1(new_n776), .B2(new_n777), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT31), .B1(new_n896), .B2(new_n779), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n865), .B1(new_n898), .B2(new_n760), .ZN(new_n899));
  INV_X1    g0699(.A(new_n472), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n366), .B(new_n723), .C1(new_n672), .C2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n723), .A2(new_n366), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n394), .A2(new_n472), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT104), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n497), .B1(new_n496), .B2(new_n492), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n312), .B(new_n906), .C1(new_n495), .C2(new_n498), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n476), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n520), .A2(new_n721), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n514), .A2(new_n487), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT37), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n905), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n522), .A2(new_n524), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n522), .A2(new_n720), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n913), .A2(new_n914), .A3(new_n911), .A4(new_n503), .ZN(new_n915));
  INV_X1    g0715(.A(new_n503), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n907), .A2(new_n476), .B1(new_n520), .B2(new_n721), .ZN(new_n917));
  OAI211_X1 g0717(.A(KEYINPUT104), .B(KEYINPUT37), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n912), .A2(new_n915), .A3(new_n918), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n504), .A2(new_n521), .A3(new_n516), .A4(new_n525), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n721), .B1(new_n907), .B2(new_n476), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AND3_X1   g0722(.A1(new_n919), .A2(KEYINPUT38), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT38), .B1(new_n919), .B2(new_n922), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n899), .B(new_n904), .C1(new_n923), .C2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT40), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n925), .A2(KEYINPUT105), .A3(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT105), .B1(new_n925), .B2(new_n926), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT38), .ZN(new_n931));
  INV_X1    g0731(.A(new_n675), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n914), .B1(new_n669), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n913), .A2(new_n914), .A3(new_n503), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(new_n911), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n931), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n919), .A2(KEYINPUT38), .A3(new_n922), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n899), .A2(new_n904), .A3(KEYINPUT40), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n928), .A2(new_n930), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n896), .A2(KEYINPUT31), .A3(new_n779), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n760), .A2(new_n782), .A3(new_n941), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n527), .A2(new_n942), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n940), .A2(new_n943), .ZN(new_n945));
  INV_X1    g0745(.A(G330), .ZN(new_n946));
  NOR3_X1   g0746(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT39), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n938), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n672), .A2(new_n366), .A3(new_n724), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NOR3_X1   g0751(.A1(new_n923), .A2(new_n924), .A3(new_n948), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n949), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n864), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n904), .B1(new_n859), .B2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n923), .A2(new_n924), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n667), .A2(new_n668), .A3(new_n721), .ZN(new_n959));
  AND3_X1   g0759(.A1(new_n954), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n527), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n677), .B1(new_n758), .B2(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n960), .B(new_n962), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n947), .A2(new_n963), .B1(new_n212), .B2(new_n789), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(new_n963), .B2(new_n947), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n528), .B(new_n221), .C1(new_n307), .C2(KEYINPUT35), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(KEYINPUT35), .B2(new_n307), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT36), .Z(new_n968));
  OR3_X1    g0768(.A1(new_n223), .A2(new_n206), .A3(new_n489), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n212), .B(G13), .C1(new_n969), .C2(new_n248), .ZN(new_n970));
  OR3_X1    g0770(.A1(new_n965), .A2(new_n968), .A3(new_n970), .ZN(G367));
  INV_X1    g0771(.A(new_n796), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n804), .B1(new_n216), .B2(new_n454), .C1(new_n972), .C2(new_n243), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n973), .A2(new_n792), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n651), .A2(new_n683), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n723), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n694), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n689), .B2(new_n976), .ZN(new_n978));
  AOI21_X1  g0778(.A(KEYINPUT46), .B1(new_n836), .B2(G116), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(G294), .B2(new_n817), .ZN(new_n980));
  INV_X1    g0780(.A(new_n837), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n981), .A2(new_n231), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(G317), .B2(new_n809), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n439), .B1(new_n829), .B2(new_n545), .ZN(new_n984));
  INV_X1    g0784(.A(new_n300), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n985), .A2(new_n826), .B1(new_n824), .B2(new_n886), .ZN(new_n986));
  AOI211_X1 g0786(.A(new_n984), .B(new_n986), .C1(G283), .C2(new_n849), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n836), .A2(KEYINPUT46), .A3(G116), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n980), .A2(new_n983), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n981), .A2(new_n206), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n990), .A2(new_n439), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT109), .Z(new_n992));
  AOI22_X1  g0792(.A1(new_n836), .A2(G58), .B1(new_n809), .B2(G137), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n826), .A2(new_n203), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n829), .A2(new_n410), .B1(new_n820), .B2(new_n201), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n994), .B(new_n995), .C1(G143), .C2(new_n823), .ZN(new_n996));
  INV_X1    g0796(.A(G159), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n993), .B(new_n996), .C1(new_n997), .C2(new_n816), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n989), .B1(new_n992), .B2(new_n998), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT47), .Z(new_n1000));
  OAI221_X1 g0800(.A(new_n974), .B1(new_n853), .B2(new_n978), .C1(new_n1000), .C2(new_n806), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n679), .B(new_n680), .C1(new_n342), .C2(new_n724), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n341), .A2(new_n723), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1004), .A2(new_n739), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT42), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n611), .B1(new_n347), .B2(new_n352), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n724), .B1(new_n1007), .B2(new_n341), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n978), .B(KEYINPUT43), .Z(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT106), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1006), .A2(new_n1008), .A3(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1009), .A2(KEYINPUT106), .A3(new_n1010), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1004), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n737), .A2(KEYINPUT107), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n737), .A2(new_n1018), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT107), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1017), .A2(new_n1022), .A3(new_n1021), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n743), .B(KEYINPUT41), .Z(new_n1027));
  NAND2_X1  g0827(.A1(new_n1004), .A2(new_n740), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT44), .Z(new_n1029));
  NOR2_X1   g0829(.A1(new_n1004), .A2(new_n740), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT45), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1032), .A2(KEYINPUT108), .A3(new_n737), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n739), .B1(new_n733), .B2(new_n738), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(new_n728), .Z(new_n1035));
  NAND3_X1  g0835(.A1(new_n735), .A2(KEYINPUT108), .A3(new_n736), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1036), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1033), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1027), .B1(new_n1038), .B2(new_n787), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1039), .A2(new_n791), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1001), .B1(new_n1026), .B2(new_n1040), .ZN(G387));
  AOI22_X1  g0841(.A1(G317), .A2(new_n830), .B1(new_n849), .B2(G303), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n844), .B2(new_n824), .C1(new_n816), .C2(new_n886), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT48), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1046));
  INV_X1    g0846(.A(G283), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n835), .A2(new_n847), .B1(new_n1047), .B2(new_n826), .ZN(new_n1048));
  OR3_X1    g0848(.A1(new_n1045), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT49), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n439), .B1(new_n872), .B2(new_n846), .C1(new_n528), .C2(new_n981), .ZN(new_n1053));
  OR3_X1    g0853(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n835), .A2(new_n206), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(KEYINPUT110), .B(G150), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1055), .B(new_n982), .C1(new_n809), .C2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n826), .A2(new_n454), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n376), .B1(new_n820), .B2(new_n203), .C1(new_n201), .C2(new_n829), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1058), .B(new_n1059), .C1(G159), .C2(new_n823), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1057), .B(new_n1060), .C1(new_n409), .C2(new_n816), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n806), .B1(new_n1054), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n796), .B1(new_n240), .B2(new_n264), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n794), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1063), .B1(new_n745), .B2(new_n1064), .ZN(new_n1065));
  OR3_X1    g0865(.A1(new_n409), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1066));
  AOI21_X1  g0866(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1067));
  OAI21_X1  g0867(.A(KEYINPUT50), .B1(new_n409), .B2(G50), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1066), .A2(new_n745), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1065), .A2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(G107), .B2(new_n216), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n793), .B(new_n1062), .C1(new_n804), .C2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n734), .A2(new_n802), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1035), .A2(new_n791), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n787), .A2(new_n1035), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n743), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n787), .A2(new_n1035), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1074), .B1(new_n1076), .B2(new_n1077), .ZN(G393));
  AOI21_X1  g0878(.A(new_n744), .B1(new_n1033), .B2(new_n1037), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1079), .A2(new_n787), .A3(new_n1035), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n796), .A2(new_n247), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1081), .B(new_n804), .C1(new_n231), .C2(new_n216), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n792), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1083), .B(KEYINPUT111), .Z(new_n1084));
  OAI221_X1 g0884(.A(new_n439), .B1(new_n826), .B2(new_n528), .C1(new_n847), .C2(new_n820), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n872), .A2(new_n844), .B1(new_n1047), .B2(new_n835), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1085), .B(new_n1086), .C1(G107), .C2(new_n837), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT52), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n823), .A2(G317), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n886), .B2(new_n829), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n817), .A2(G303), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1087), .B(new_n1091), .C1(new_n1088), .C2(new_n1090), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n824), .A2(new_n410), .B1(new_n829), .B2(new_n997), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT51), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n817), .A2(G50), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n826), .A2(new_n206), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n439), .B(new_n1096), .C1(new_n451), .C2(new_n849), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1094), .A2(new_n1095), .A3(new_n885), .A4(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n836), .A2(G68), .B1(new_n809), .B2(G143), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT112), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1092), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1084), .B1(new_n1101), .B2(new_n803), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n1018), .B2(new_n853), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n791), .B1(new_n1075), .B2(new_n743), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1032), .B(new_n737), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1080), .B(new_n1103), .C1(new_n1104), .C2(new_n1105), .ZN(G390));
  AND2_X1   g0906(.A1(new_n901), .A2(new_n903), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n858), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n710), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1107), .B1(new_n1109), .B2(new_n864), .ZN(new_n1110));
  AOI21_X1  g0910(.A(KEYINPUT39), .B1(new_n936), .B2(new_n937), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n1110), .A2(new_n951), .B1(new_n1111), .B2(new_n952), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n786), .A2(new_n892), .A3(new_n904), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n951), .B1(new_n936), .B2(new_n937), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT113), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n689), .B1(new_n681), .B2(new_n754), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n750), .A2(new_n752), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n724), .B(new_n863), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n864), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n904), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1114), .A2(new_n1115), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1115), .B1(new_n1114), .B2(new_n1120), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1112), .B(new_n1113), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1120), .A2(new_n938), .A3(new_n950), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(KEYINPUT113), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1114), .A2(new_n1115), .A3(new_n1120), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n949), .A2(new_n953), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n956), .A2(new_n950), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n1125), .A2(new_n1126), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT114), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n942), .A2(G330), .A3(new_n892), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1130), .B1(new_n1107), .B2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n899), .A2(new_n904), .A3(KEYINPUT114), .A4(G330), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1123), .B1(new_n1129), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1107), .B1(new_n785), .B2(new_n865), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1132), .A2(new_n1136), .A3(new_n1133), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1109), .A2(new_n864), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1107), .A2(new_n1131), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1113), .A2(new_n864), .A3(new_n1118), .A4(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n900), .B1(new_n672), .B2(new_n366), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n431), .A2(new_n468), .A3(new_n436), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1144), .A2(new_n920), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n942), .A2(G330), .A3(new_n1143), .A4(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(KEYINPUT115), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT115), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n527), .A2(new_n1148), .A3(G330), .A4(new_n942), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1150), .B(new_n677), .C1(new_n758), .C2(new_n961), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1142), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n744), .B1(new_n1135), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1151), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1123), .B(new_n1155), .C1(new_n1129), .C2(new_n1134), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n870), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n875), .B1(new_n226), .B2(new_n835), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n439), .B1(new_n820), .B2(new_n231), .C1(new_n528), .C2(new_n829), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1096), .B(new_n1160), .C1(G283), .C2(new_n823), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n985), .B2(new_n816), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1159), .B(new_n1162), .C1(G294), .C2(new_n809), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n809), .A2(G125), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1164), .B(new_n376), .C1(new_n981), .C2(new_n201), .ZN(new_n1165));
  XOR2_X1   g0965(.A(new_n1165), .B(KEYINPUT116), .Z(new_n1166));
  NAND2_X1  g0966(.A1(new_n836), .A2(new_n1056), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT53), .ZN(new_n1168));
  INV_X1    g0968(.A(G128), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n824), .A2(new_n1169), .B1(new_n829), .B2(new_n873), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT117), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n816), .A2(new_n879), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT54), .B(G143), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n820), .A2(new_n1173), .B1(new_n826), .B2(new_n997), .ZN(new_n1174));
  NOR4_X1   g0974(.A1(new_n1168), .A2(new_n1171), .A3(new_n1172), .A4(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1163), .B1(new_n1166), .B2(new_n1175), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n792), .B1(new_n451), .B2(new_n1158), .C1(new_n1176), .C2(new_n806), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n1127), .B2(new_n800), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT118), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1123), .B(new_n791), .C1(new_n1129), .C2(new_n1134), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1157), .A2(new_n1182), .ZN(G378));
  AOI21_X1  g0983(.A(new_n946), .B1(new_n939), .B2(new_n938), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n927), .B2(new_n929), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n431), .A2(new_n436), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n720), .A2(new_n435), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1186), .B(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1188), .B(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1185), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1190), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1184), .B(new_n1192), .C1(new_n927), .C2(new_n929), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n960), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1191), .A2(new_n960), .A3(new_n1193), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1190), .A2(new_n800), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n792), .B1(G50), .B2(new_n1158), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n376), .A2(G41), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1201), .B1(new_n296), .B2(new_n829), .C1(new_n454), .C2(new_n820), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n994), .B(new_n1202), .C1(G116), .C2(new_n823), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n231), .B2(new_n816), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n872), .A2(new_n1047), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n981), .A2(new_n202), .ZN(new_n1206));
  NOR4_X1   g1006(.A1(new_n1204), .A2(new_n1055), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  OR2_X1    g1007(.A1(new_n1207), .A2(KEYINPUT58), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n826), .A2(new_n410), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n829), .A2(new_n1169), .B1(new_n820), .B2(new_n879), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1209), .B(new_n1210), .C1(G125), .C2(new_n823), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1211), .B1(new_n835), .B2(new_n1173), .C1(new_n873), .C2(new_n816), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1212), .A2(KEYINPUT59), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(KEYINPUT59), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(KEYINPUT119), .B(G124), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n288), .B(new_n256), .C1(new_n872), .C2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G159), .B2(new_n837), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1213), .A2(new_n1214), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1207), .A2(KEYINPUT58), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1201), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1220), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1208), .A2(new_n1218), .A3(new_n1219), .A4(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1200), .B1(new_n1222), .B2(new_n803), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1198), .A2(new_n791), .B1(new_n1199), .B2(new_n1223), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n1191), .A2(new_n960), .A3(new_n1193), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n960), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1226));
  OAI21_X1  g1026(.A(KEYINPUT57), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  AND2_X1   g1027(.A1(new_n1156), .A2(new_n1152), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n743), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1156), .A2(new_n1152), .ZN(new_n1230));
  AOI21_X1  g1030(.A(KEYINPUT57), .B1(new_n1198), .B2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1224), .B1(new_n1229), .B2(new_n1231), .ZN(G375));
  XNOR2_X1  g1032(.A(new_n790), .B(KEYINPUT120), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1107), .A2(new_n800), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n792), .B1(G68), .B2(new_n1158), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n376), .B1(new_n820), .B2(new_n410), .C1(new_n879), .C2(new_n829), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n824), .A2(new_n873), .B1(new_n826), .B2(new_n201), .ZN(new_n1237));
  NOR3_X1   g1037(.A1(new_n1206), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n816), .B2(new_n1173), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n872), .A2(new_n1169), .B1(new_n997), .B2(new_n835), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT121), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n990), .B1(G97), .B2(new_n836), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1242), .B1(new_n545), .B2(new_n872), .ZN(new_n1243));
  OAI221_X1 g1043(.A(new_n439), .B1(new_n829), .B2(new_n1047), .C1(new_n985), .C2(new_n820), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n1058), .B(new_n1244), .C1(G294), .C2(new_n823), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1245), .B1(new_n528), .B2(new_n816), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n1239), .A2(new_n1241), .B1(new_n1243), .B2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1235), .B1(new_n1247), .B2(new_n803), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n1142), .A2(new_n1233), .B1(new_n1234), .B2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT122), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1249), .B(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1027), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1139), .A2(new_n1151), .A3(new_n1141), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1153), .A2(new_n1252), .A3(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1251), .A2(new_n1254), .ZN(G381));
  OR2_X1    g1055(.A1(G393), .A2(G396), .ZN(new_n1256));
  OR4_X1    g1056(.A1(G384), .A2(G387), .A3(new_n1256), .A4(G390), .ZN(new_n1257));
  OR4_X1    g1057(.A1(G378), .A2(new_n1257), .A3(G375), .A4(G381), .ZN(G407));
  AOI21_X1  g1058(.A(new_n1181), .B1(new_n1156), .B2(new_n1154), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n722), .A2(G213), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1262));
  OAI211_X1 g1062(.A(G407), .B(G213), .C1(G375), .C2(new_n1262), .ZN(G409));
  INV_X1    g1063(.A(KEYINPUT124), .ZN(new_n1264));
  XOR2_X1   g1064(.A(G393), .B(G396), .Z(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1024), .B(new_n1025), .C1(new_n1039), .C2(new_n791), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1267), .A2(new_n1001), .A3(G390), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(G390), .B1(new_n1267), .B2(new_n1001), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1266), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(G390), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(G387), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1273), .A2(new_n1265), .A3(new_n1268), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1271), .A2(KEYINPUT123), .A3(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT123), .B1(new_n1271), .B2(new_n1274), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT61), .ZN(new_n1278));
  OAI211_X1 g1078(.A(G378), .B(new_n1224), .C1(new_n1229), .C2(new_n1231), .ZN(new_n1279));
  AND3_X1   g1079(.A1(new_n1198), .A2(new_n1252), .A3(new_n1230), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1233), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1199), .A2(new_n1223), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1259), .B1(new_n1280), .B2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1261), .B1(new_n1279), .B2(new_n1284), .ZN(new_n1285));
  AND2_X1   g1085(.A1(new_n869), .A2(new_n893), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(new_n1249), .B(KEYINPUT122), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1139), .A2(new_n1151), .A3(KEYINPUT60), .A4(new_n1141), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n743), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1153), .A2(KEYINPUT60), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1289), .B1(new_n1290), .B2(new_n1253), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1286), .B1(new_n1287), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1291), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1293), .A2(new_n1251), .A3(G384), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1292), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(G2897), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1260), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1292), .B(new_n1294), .C1(new_n1296), .C2(new_n1260), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1278), .B1(new_n1285), .B2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT62), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1295), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1302), .B1(new_n1285), .B2(new_n1303), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1301), .A2(new_n1304), .ZN(new_n1305));
  AOI211_X1 g1105(.A(new_n1261), .B(new_n1295), .C1(new_n1279), .C2(new_n1284), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1302), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1277), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1285), .A2(KEYINPUT63), .A3(new_n1303), .ZN(new_n1309));
  OAI211_X1 g1109(.A(new_n1309), .B(new_n1278), .C1(new_n1285), .C2(new_n1300), .ZN(new_n1310));
  AND2_X1   g1110(.A1(new_n1271), .A2(new_n1274), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1311), .B1(new_n1306), .B2(KEYINPUT63), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1310), .A2(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1264), .B1(new_n1308), .B2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1301), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1285), .A2(new_n1303), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT63), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1315), .A2(new_n1318), .A3(new_n1311), .A4(new_n1309), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1316), .A2(KEYINPUT62), .ZN(new_n1320));
  NOR3_X1   g1120(.A1(new_n1320), .A2(new_n1301), .A3(new_n1304), .ZN(new_n1321));
  OAI211_X1 g1121(.A(KEYINPUT124), .B(new_n1319), .C1(new_n1321), .C2(new_n1277), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1314), .A2(new_n1322), .ZN(G405));
  NAND2_X1  g1123(.A1(G375), .A2(new_n1259), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1324), .A2(new_n1295), .A3(new_n1279), .ZN(new_n1325));
  AND2_X1   g1125(.A1(new_n1325), .A2(KEYINPUT126), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1325), .A2(KEYINPUT126), .ZN(new_n1327));
  OR2_X1    g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1324), .A2(new_n1279), .ZN(new_n1329));
  AND3_X1   g1129(.A1(new_n1329), .A2(KEYINPUT125), .A3(new_n1303), .ZN(new_n1330));
  AOI21_X1  g1130(.A(KEYINPUT125), .B1(new_n1329), .B2(new_n1303), .ZN(new_n1331));
  OR2_X1    g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  OAI21_X1  g1132(.A(KEYINPUT127), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT127), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1277), .A2(new_n1334), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1328), .A2(new_n1332), .A3(new_n1333), .A4(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1333), .ZN(new_n1337));
  OAI22_X1  g1137(.A1(new_n1327), .A2(new_n1326), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1336), .A2(new_n1339), .ZN(G402));
endmodule


