//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n993, new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041;
  XNOR2_X1  g000(.A(G110), .B(G140), .ZN(new_n187));
  INV_X1    g001(.A(G227), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G953), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT77), .ZN(new_n191));
  INV_X1    g005(.A(G104), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT3), .B1(new_n192), .B2(G107), .ZN(new_n193));
  AOI21_X1  g007(.A(G101), .B1(new_n192), .B2(G107), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n196), .A3(G104), .ZN(new_n197));
  AND3_X1   g011(.A1(new_n193), .A2(new_n194), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G101), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n196), .A2(G104), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n192), .A2(G107), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n199), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n191), .B1(new_n198), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT64), .B1(new_n204), .B2(G146), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(G143), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n204), .A2(G146), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n205), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n204), .A2(G146), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT1), .ZN(new_n212));
  OAI21_X1  g026(.A(G128), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(G143), .B(G146), .ZN(new_n214));
  INV_X1    g028(.A(G128), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(KEYINPUT1), .ZN(new_n216));
  AOI22_X1  g030(.A1(new_n210), .A2(new_n213), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n202), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n193), .A2(new_n194), .A3(new_n197), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT77), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n203), .A2(new_n217), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n214), .A2(new_n216), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n207), .A2(G143), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n215), .B1(new_n223), .B2(KEYINPUT1), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n222), .B1(new_n214), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(new_n219), .A3(new_n218), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n221), .A2(KEYINPUT78), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(KEYINPUT78), .B1(new_n221), .B2(new_n226), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT11), .ZN(new_n229));
  INV_X1    g043(.A(G134), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n229), .B1(new_n230), .B2(G137), .ZN(new_n231));
  INV_X1    g045(.A(G137), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(KEYINPUT11), .A3(G134), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n230), .A2(G137), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n231), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G131), .ZN(new_n236));
  AND2_X1   g050(.A1(KEYINPUT65), .A2(G131), .ZN(new_n237));
  NOR2_X1   g051(.A1(KEYINPUT65), .A2(G131), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n239), .A2(new_n231), .A3(new_n233), .A4(new_n234), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n236), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NOR3_X1   g056(.A1(new_n227), .A2(new_n228), .A3(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT79), .B1(new_n243), .B2(KEYINPUT12), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n221), .A2(new_n226), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT78), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n221), .A2(KEYINPUT78), .A3(new_n226), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(new_n241), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT79), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT12), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n242), .A2(new_n251), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n244), .A2(new_n252), .B1(new_n245), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n203), .A2(new_n220), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT10), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n217), .A2(new_n256), .ZN(new_n257));
  AOI22_X1  g071(.A1(new_n255), .A2(new_n257), .B1(new_n226), .B2(new_n256), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n193), .A2(new_n197), .A3(new_n201), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G101), .ZN(new_n260));
  OAI21_X1  g074(.A(KEYINPUT76), .B1(new_n260), .B2(KEYINPUT4), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT76), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n259), .A2(new_n262), .A3(new_n263), .A4(G101), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  AND2_X1   g079(.A1(KEYINPUT0), .A2(G128), .ZN(new_n266));
  NOR2_X1   g080(.A1(KEYINPUT0), .A2(G128), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI22_X1  g082(.A1(new_n210), .A2(new_n268), .B1(new_n266), .B2(new_n214), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n260), .A2(KEYINPUT4), .A3(new_n219), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n265), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n258), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n272), .A2(new_n241), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n190), .B1(new_n254), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n190), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n272), .A2(new_n241), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n274), .A2(G469), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G469), .ZN(new_n279));
  INV_X1    g093(.A(G902), .ZN(new_n280));
  INV_X1    g094(.A(new_n275), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n244), .A2(new_n252), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n245), .A2(new_n253), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n190), .ZN(new_n285));
  INV_X1    g099(.A(new_n273), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n285), .B1(new_n286), .B2(new_n276), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n279), .B(new_n280), .C1(new_n284), .C2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(G469), .A2(G902), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n278), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G221), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT75), .ZN(new_n292));
  INV_X1    g106(.A(G234), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n293), .A2(KEYINPUT9), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n293), .A2(KEYINPUT9), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n292), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(KEYINPUT9), .B(G234), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT75), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n291), .B1(new_n299), .B2(new_n280), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n290), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G237), .ZN(new_n304));
  INV_X1    g118(.A(G953), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n305), .A3(G214), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n204), .ZN(new_n307));
  NOR2_X1   g121(.A1(G237), .A2(G953), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(G143), .A3(G214), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n239), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT17), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n307), .A2(new_n239), .A3(new_n309), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G140), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G125), .ZN(new_n317));
  INV_X1    g131(.A(G125), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G140), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n317), .A2(new_n319), .A3(KEYINPUT16), .ZN(new_n320));
  OR3_X1    g134(.A1(new_n318), .A2(KEYINPUT16), .A3(G140), .ZN(new_n321));
  AND3_X1   g135(.A1(new_n320), .A2(G146), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(G146), .B1(new_n320), .B2(new_n321), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n315), .B(new_n324), .C1(new_n313), .C2(new_n312), .ZN(new_n325));
  XOR2_X1   g139(.A(G113), .B(G122), .Z(new_n326));
  XOR2_X1   g140(.A(KEYINPUT88), .B(G104), .Z(new_n327));
  XOR2_X1   g141(.A(new_n326), .B(new_n327), .Z(new_n328));
  AND2_X1   g142(.A1(new_n317), .A2(new_n319), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n329), .B(new_n207), .ZN(new_n330));
  NAND2_X1  g144(.A1(KEYINPUT18), .A2(G131), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n307), .A2(new_n309), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n331), .ZN(new_n333));
  AOI21_X1  g147(.A(KEYINPUT85), .B1(new_n310), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT85), .ZN(new_n335));
  AOI211_X1 g149(.A(new_n335), .B(new_n331), .C1(new_n307), .C2(new_n309), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n330), .B(new_n332), .C1(new_n334), .C2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n325), .A2(new_n328), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT89), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n325), .A2(new_n337), .A3(KEYINPUT89), .A4(new_n328), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n312), .A2(new_n314), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n320), .A2(new_n321), .A3(G146), .ZN(new_n344));
  NAND2_X1  g158(.A1(KEYINPUT86), .A2(KEYINPUT19), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n329), .A2(new_n345), .ZN(new_n346));
  XOR2_X1   g160(.A(KEYINPUT86), .B(KEYINPUT19), .Z(new_n347));
  OAI21_X1  g161(.A(new_n346), .B1(new_n329), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n344), .B1(new_n348), .B2(G146), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n337), .B1(new_n343), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT87), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n328), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n337), .B(KEYINPUT87), .C1(new_n343), .C2(new_n349), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n342), .A2(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(G475), .A2(G902), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT90), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n359), .B1(new_n342), .B2(new_n355), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n358), .B1(KEYINPUT20), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n356), .A2(KEYINPUT90), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT20), .ZN(new_n363));
  INV_X1    g177(.A(new_n357), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n364), .B1(new_n342), .B2(new_n355), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n362), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n325), .A2(new_n337), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n342), .B1(new_n328), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n280), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n361), .A2(new_n366), .B1(G475), .B2(new_n369), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n305), .A2(G217), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n296), .A2(new_n298), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT93), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n296), .A2(new_n298), .A3(KEYINPUT93), .A4(new_n371), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n204), .A2(G128), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n215), .A2(G143), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n376), .A2(new_n377), .A3(new_n230), .ZN(new_n378));
  INV_X1    g192(.A(G116), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G122), .ZN(new_n380));
  INV_X1    g194(.A(G122), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G116), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n380), .A2(new_n382), .A3(new_n196), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n381), .A2(G116), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n379), .A2(G122), .ZN(new_n385));
  OAI21_X1  g199(.A(G107), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n378), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT13), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n376), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n204), .A2(KEYINPUT13), .A3(G128), .ZN(new_n390));
  AND3_X1   g204(.A1(new_n389), .A2(new_n377), .A3(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n387), .B1(new_n230), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n230), .B1(new_n376), .B2(new_n377), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n383), .B1(new_n378), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(KEYINPUT14), .B1(new_n381), .B2(G116), .ZN(new_n395));
  OAI21_X1  g209(.A(KEYINPUT91), .B1(new_n395), .B2(new_n384), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT91), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n397), .B(new_n380), .C1(new_n385), .C2(KEYINPUT14), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n396), .B(new_n398), .C1(KEYINPUT14), .C2(new_n380), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n394), .B1(new_n399), .B2(G107), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT92), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n392), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n380), .A2(KEYINPUT14), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n380), .B1(new_n385), .B2(KEYINPUT14), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n403), .B1(new_n404), .B2(KEYINPUT91), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n196), .B1(new_n405), .B2(new_n398), .ZN(new_n406));
  NOR3_X1   g220(.A1(new_n406), .A2(KEYINPUT92), .A3(new_n394), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n374), .B(new_n375), .C1(new_n402), .C2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT94), .ZN(new_n409));
  OAI21_X1  g223(.A(KEYINPUT92), .B1(new_n406), .B2(new_n394), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n400), .A2(new_n401), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n374), .A2(new_n375), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n410), .A2(new_n411), .A3(new_n412), .A4(new_n392), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n408), .A2(new_n409), .A3(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n402), .A2(new_n407), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(KEYINPUT94), .A3(new_n412), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(new_n280), .A3(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G478), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n418), .A2(KEYINPUT15), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n417), .B(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n305), .A2(G952), .ZN(new_n422));
  NAND2_X1  g236(.A1(G234), .A2(G237), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(KEYINPUT21), .B(G898), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n425), .B(KEYINPUT95), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n423), .A2(G902), .A3(G953), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n424), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  XOR2_X1   g242(.A(new_n428), .B(KEYINPUT96), .Z(new_n429));
  NAND3_X1  g243(.A1(new_n370), .A2(new_n421), .A3(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(G214), .B1(G237), .B2(G902), .ZN(new_n431));
  XOR2_X1   g245(.A(new_n431), .B(KEYINPUT80), .Z(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(G110), .B(G122), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  OR2_X1    g249(.A1(KEYINPUT66), .A2(G119), .ZN(new_n436));
  NAND2_X1  g250(.A1(KEYINPUT66), .A2(G119), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(G116), .A3(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n438), .A2(KEYINPUT67), .ZN(new_n439));
  INV_X1    g253(.A(G119), .ZN(new_n440));
  OAI21_X1  g254(.A(KEYINPUT67), .B1(new_n440), .B2(G116), .ZN(new_n441));
  AND2_X1   g255(.A1(KEYINPUT66), .A2(G119), .ZN(new_n442));
  NOR2_X1   g256(.A1(KEYINPUT66), .A2(G119), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n441), .B1(new_n444), .B2(G116), .ZN(new_n445));
  OAI21_X1  g259(.A(KEYINPUT5), .B1(new_n439), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G113), .B1(new_n438), .B2(KEYINPUT5), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(KEYINPUT2), .B(G113), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n451), .B1(new_n439), .B2(new_n445), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n449), .A2(KEYINPUT81), .A3(new_n452), .A4(new_n255), .ZN(new_n453));
  INV_X1    g267(.A(new_n441), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n438), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT67), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n444), .A2(new_n456), .A3(G116), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n455), .A2(new_n457), .A3(new_n450), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n452), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(new_n265), .A3(new_n270), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n453), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n450), .B1(new_n455), .B2(new_n457), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n462), .B1(new_n446), .B2(new_n448), .ZN(new_n463));
  AOI21_X1  g277(.A(KEYINPUT81), .B1(new_n463), .B2(new_n255), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n435), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT81), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT5), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n467), .B1(new_n455), .B2(new_n457), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n452), .B1(new_n468), .B2(new_n447), .ZN(new_n469));
  INV_X1    g283(.A(new_n255), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n471), .A2(new_n434), .A3(new_n460), .A4(new_n453), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n465), .A2(KEYINPUT6), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT6), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n474), .B(new_n435), .C1(new_n461), .C2(new_n464), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n210), .A2(new_n213), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n222), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n477), .A2(G125), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n269), .A2(new_n318), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  XOR2_X1   g294(.A(KEYINPUT82), .B(G224), .Z(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n305), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT83), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n481), .A2(KEYINPUT83), .A3(new_n305), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n480), .B(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n473), .A2(new_n475), .A3(new_n487), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n484), .A2(KEYINPUT7), .A3(new_n485), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n490), .B1(new_n479), .B2(new_n478), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n480), .A2(new_n489), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n469), .B1(new_n198), .B2(new_n202), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n494), .B1(new_n470), .B2(new_n469), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n434), .B(KEYINPUT8), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(G902), .B1(new_n497), .B2(new_n472), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n488), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(G210), .B1(G237), .B2(G902), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n500), .A2(KEYINPUT84), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n501), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n503), .B1(new_n488), .B2(new_n498), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n433), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n430), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G131), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n232), .A2(G134), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n507), .B1(new_n508), .B2(new_n234), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n231), .A2(new_n233), .A3(new_n234), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n509), .B1(new_n510), .B2(new_n239), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n477), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT30), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n241), .A2(new_n269), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n513), .B1(new_n512), .B2(new_n514), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n459), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n512), .A2(new_n514), .A3(new_n458), .A4(new_n452), .ZN(new_n518));
  XOR2_X1   g332(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n519));
  NAND2_X1  g333(.A1(new_n308), .A2(G210), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT26), .B(G101), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n521), .B(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n517), .A2(new_n518), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT31), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n512), .A2(new_n514), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n459), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT28), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n528), .B1(new_n529), .B2(new_n518), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n518), .A2(new_n529), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n523), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT31), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n517), .A2(new_n533), .A3(new_n518), .A4(new_n524), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n526), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G472), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(new_n536), .A3(new_n280), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT69), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT32), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n535), .A2(KEYINPUT69), .A3(new_n536), .A4(new_n280), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n530), .A2(new_n531), .A3(new_n523), .ZN(new_n543));
  OR2_X1    g357(.A1(new_n543), .A2(KEYINPUT29), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n517), .A2(new_n518), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n546), .A2(new_n524), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n280), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT70), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n518), .A2(new_n549), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n452), .A2(new_n458), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n551), .A2(KEYINPUT70), .A3(new_n514), .A4(new_n512), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n550), .A2(new_n552), .A3(new_n528), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n531), .B1(new_n553), .B2(KEYINPUT28), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n554), .A2(KEYINPUT29), .A3(new_n524), .ZN(new_n555));
  OAI21_X1  g369(.A(G472), .B1(new_n548), .B2(new_n555), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n535), .A2(KEYINPUT32), .A3(new_n536), .A4(new_n280), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT71), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n557), .A2(new_n558), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n542), .B(new_n556), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT22), .B(G137), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n291), .A2(new_n293), .A3(G953), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n562), .B(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(G128), .B1(new_n442), .B2(new_n443), .ZN(new_n565));
  NOR2_X1   g379(.A1(G119), .A2(G128), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(KEYINPUT23), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(G110), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n215), .B1(new_n442), .B2(new_n443), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT23), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n568), .A2(new_n569), .A3(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT24), .B(G110), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n565), .A2(new_n567), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n329), .A2(new_n207), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n344), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n574), .B1(new_n565), .B2(new_n567), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n320), .A2(new_n321), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n207), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n581), .B1(new_n583), .B2(new_n344), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n568), .A2(new_n572), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(G110), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n564), .B1(new_n580), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT73), .ZN(new_n589));
  INV_X1    g403(.A(new_n574), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n215), .B1(new_n436), .B2(new_n437), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n590), .B1(new_n591), .B2(new_n566), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n592), .B1(new_n322), .B2(new_n323), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n569), .B1(new_n568), .B2(new_n572), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n578), .B1(new_n573), .B2(new_n575), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n589), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n580), .A2(new_n587), .A3(KEYINPUT73), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n588), .B1(new_n599), .B2(new_n564), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(G902), .B1(new_n293), .B2(G217), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT74), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n604), .B(KEYINPUT25), .C1(new_n600), .C2(G902), .ZN(new_n605));
  OAI21_X1  g419(.A(G217), .B1(new_n293), .B2(G902), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(KEYINPUT72), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n564), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n609), .B1(new_n597), .B2(new_n598), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n280), .B1(new_n610), .B2(new_n588), .ZN(new_n611));
  AOI21_X1  g425(.A(KEYINPUT25), .B1(new_n611), .B2(new_n604), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n603), .B1(new_n608), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n303), .A2(new_n506), .A3(new_n561), .A4(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G101), .ZN(G3));
  NAND2_X1  g430(.A1(new_n499), .A2(new_n500), .ZN(new_n617));
  INV_X1    g431(.A(new_n500), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n488), .A2(new_n498), .A3(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n617), .A2(new_n433), .A3(new_n429), .A4(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT97), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n412), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n374), .A2(KEYINPUT97), .A3(new_n375), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(KEYINPUT98), .B1(new_n415), .B2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n626), .B1(new_n415), .B2(new_n412), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n410), .A2(new_n411), .A3(new_n392), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT98), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n628), .A2(new_n629), .A3(new_n622), .A4(new_n623), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n625), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(KEYINPUT99), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT99), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n625), .A2(new_n627), .A3(new_n633), .A4(new_n630), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n414), .A2(new_n416), .ZN(new_n635));
  AOI22_X1  g449(.A1(new_n632), .A2(new_n634), .B1(new_n635), .B2(new_n626), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n418), .A2(G902), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n417), .A2(new_n418), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n417), .A2(KEYINPUT100), .A3(new_n418), .ZN(new_n641));
  AOI22_X1  g455(.A1(new_n636), .A2(new_n637), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n620), .A2(new_n642), .A3(new_n370), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n535), .A2(new_n280), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(G472), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n539), .A2(new_n541), .A3(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n646), .A2(new_n613), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n303), .A2(new_n643), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT34), .B(G104), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G6));
  NAND2_X1  g464(.A1(new_n369), .A2(G475), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n358), .A2(KEYINPUT20), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n365), .A2(new_n363), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n620), .A2(new_n421), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n303), .A2(new_n655), .A3(new_n647), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT35), .B(G107), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G9));
  INV_X1    g472(.A(new_n599), .ZN(new_n659));
  OR2_X1    g473(.A1(new_n564), .A2(KEYINPUT36), .ZN(new_n660));
  OR2_X1    g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n661), .A2(new_n602), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n663), .B1(new_n608), .B2(new_n612), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n646), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n303), .A2(new_n506), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT37), .B(G110), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G12));
  INV_X1    g483(.A(G900), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n423), .A2(new_n670), .A3(G902), .A4(G953), .ZN(new_n671));
  OR2_X1    g485(.A1(new_n671), .A2(KEYINPUT101), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(KEYINPUT101), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n672), .A2(new_n424), .A3(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n651), .B(new_n675), .C1(new_n652), .C2(new_n653), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(new_n421), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n290), .A2(new_n677), .A3(new_n301), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n432), .B1(new_n499), .B2(new_n500), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n619), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n678), .A2(new_n561), .A3(new_n681), .A4(new_n664), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  NOR2_X1   g497(.A1(new_n502), .A2(new_n504), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n365), .B1(new_n362), .B2(new_n363), .ZN(new_n687));
  AND4_X1   g501(.A1(new_n359), .A2(new_n356), .A3(new_n363), .A4(new_n357), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n651), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n420), .ZN(new_n690));
  NOR4_X1   g504(.A1(new_n686), .A2(new_n432), .A3(new_n664), .A4(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n674), .B(KEYINPUT39), .Z(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  OR3_X1    g507(.A1(new_n302), .A2(KEYINPUT40), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(KEYINPUT40), .B1(new_n302), .B2(new_n693), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n553), .A2(new_n523), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n525), .ZN(new_n697));
  AOI21_X1  g511(.A(G902), .B1(new_n697), .B2(KEYINPUT103), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n698), .B1(KEYINPUT103), .B2(new_n697), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(G472), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n542), .B(new_n700), .C1(new_n559), .C2(new_n560), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n691), .A2(new_n694), .A3(new_n695), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G143), .ZN(G45));
  NAND2_X1  g517(.A1(new_n632), .A2(new_n634), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n635), .A2(new_n626), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n704), .A2(new_n705), .A3(new_n637), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n640), .A2(new_n641), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(new_n689), .A3(new_n675), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n302), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n710), .A2(new_n561), .A3(new_n681), .A4(new_n664), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G146), .ZN(G48));
  AND3_X1   g526(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n250), .B1(new_n249), .B2(new_n251), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n283), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n287), .B1(new_n715), .B2(new_n275), .ZN(new_n716));
  OAI21_X1  g530(.A(G469), .B1(new_n716), .B2(G902), .ZN(new_n717));
  AND3_X1   g531(.A1(new_n717), .A2(new_n301), .A3(new_n288), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n643), .A2(new_n561), .A3(new_n614), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT41), .B(G113), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G15));
  NAND4_X1  g535(.A1(new_n655), .A2(new_n561), .A3(new_n614), .A4(new_n718), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G116), .ZN(G18));
  INV_X1    g537(.A(KEYINPUT104), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n718), .A2(new_n724), .A3(new_n681), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n717), .A2(new_n301), .A3(new_n288), .ZN(new_n726));
  OAI21_X1  g540(.A(KEYINPUT104), .B1(new_n726), .B2(new_n680), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n430), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n561), .A2(new_n729), .A3(new_n664), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G119), .ZN(G21));
  NAND4_X1  g546(.A1(new_n717), .A2(new_n301), .A3(new_n288), .A4(new_n429), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n689), .A2(new_n679), .A3(new_n420), .A4(new_n619), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT107), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n526), .B(new_n534), .C1(new_n554), .C2(new_n524), .ZN(new_n737));
  NOR2_X1   g551(.A1(G472), .A2(G902), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(KEYINPUT105), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT105), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n737), .A2(new_n741), .A3(new_n738), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(KEYINPUT106), .B(G472), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n744), .B1(new_n535), .B2(new_n280), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  AND4_X1   g560(.A1(new_n736), .A2(new_n743), .A3(new_n614), .A4(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n745), .B1(new_n740), .B2(new_n742), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n736), .B1(new_n748), .B2(new_n614), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n735), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G122), .ZN(G24));
  AND3_X1   g565(.A1(new_n737), .A2(new_n741), .A3(new_n738), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n741), .B1(new_n737), .B2(new_n738), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n664), .B(new_n746), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT108), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n743), .A2(KEYINPUT108), .A3(new_n664), .A4(new_n746), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n709), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n728), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G125), .ZN(G27));
  NOR3_X1   g574(.A1(new_n502), .A2(new_n432), .A3(new_n504), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n561), .A2(new_n614), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n302), .A2(KEYINPUT109), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT109), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n290), .A2(new_n764), .A3(new_n301), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n762), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n709), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT42), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n761), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n769), .B1(new_n763), .B2(new_n765), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n556), .A2(new_n557), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n537), .A2(new_n540), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n614), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT42), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n773), .A2(new_n774), .A3(new_n709), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n770), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g591(.A(KEYINPUT110), .B1(new_n768), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n763), .A2(new_n765), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n561), .A2(new_n614), .A3(new_n761), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n779), .A2(new_n780), .A3(new_n767), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n774), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT110), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n783), .A3(new_n776), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n778), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(new_n507), .ZN(G33));
  NAND3_X1  g600(.A1(new_n779), .A2(new_n780), .A3(new_n677), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G134), .ZN(G36));
  INV_X1    g602(.A(new_n288), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n274), .A2(new_n277), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT45), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n274), .A2(KEYINPUT45), .A3(new_n277), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(G469), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n289), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT46), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n789), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n794), .A2(KEYINPUT46), .A3(new_n289), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n300), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n799), .A2(new_n692), .ZN(new_n800));
  OAI21_X1  g614(.A(KEYINPUT43), .B1(new_n642), .B2(new_n689), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT43), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n708), .A2(new_n802), .A3(new_n370), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n646), .A2(new_n664), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT44), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(KEYINPUT44), .B1(new_n804), .B2(new_n805), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n808), .A2(new_n769), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n800), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G137), .ZN(G39));
  NOR2_X1   g626(.A1(KEYINPUT111), .A2(KEYINPUT47), .ZN(new_n813));
  OR2_X1    g627(.A1(new_n799), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n799), .A2(new_n815), .ZN(new_n816));
  NOR4_X1   g630(.A1(new_n561), .A2(new_n769), .A3(new_n709), .A4(new_n614), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n814), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G140), .ZN(G42));
  NOR2_X1   g633(.A1(G952), .A2(G953), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n764), .B1(new_n290), .B2(new_n301), .ZN(new_n822));
  INV_X1    g636(.A(new_n765), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n758), .B(new_n761), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n769), .A2(new_n420), .A3(new_n676), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n825), .A2(new_n561), .A3(new_n303), .A4(new_n664), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n787), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT114), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n787), .A2(new_n824), .A3(KEYINPUT114), .A4(new_n826), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XOR2_X1   g645(.A(new_n674), .B(KEYINPUT115), .Z(new_n832));
  NAND2_X1  g646(.A1(new_n665), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n734), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n303), .A2(new_n701), .A3(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n759), .A2(new_n711), .A3(new_n682), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT52), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n561), .A2(new_n681), .A3(new_n664), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n838), .B1(new_n678), .B2(new_n710), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT52), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n839), .A2(new_n759), .A3(new_n840), .A4(new_n835), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n831), .A2(new_n837), .A3(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n731), .A2(new_n719), .A3(new_n722), .A4(new_n750), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT112), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n844), .B1(new_n642), .B2(new_n370), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n708), .A2(KEYINPUT112), .A3(new_n689), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n370), .A2(new_n420), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n433), .B(new_n429), .C1(new_n502), .C2(new_n504), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n848), .A2(new_n303), .A3(new_n647), .A4(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n851), .A2(new_n667), .A3(new_n615), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(KEYINPUT113), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n302), .A2(new_n505), .A3(new_n430), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n561), .A2(new_n614), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n854), .B1(new_n855), .B2(new_n666), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT113), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n856), .A2(new_n857), .A3(new_n851), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n843), .B1(new_n853), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(new_n778), .A3(new_n784), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n821), .B1(new_n842), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n837), .A2(new_n841), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n862), .B1(new_n829), .B2(new_n830), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n561), .A2(new_n729), .A3(new_n664), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n864), .B1(new_n725), .B2(new_n727), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n750), .A2(new_n719), .ZN(new_n866));
  INV_X1    g680(.A(new_n722), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  AND4_X1   g682(.A1(new_n857), .A2(new_n851), .A3(new_n667), .A4(new_n615), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n857), .B1(new_n856), .B2(new_n851), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT53), .B1(new_n768), .B2(new_n777), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n863), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n861), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n783), .B1(new_n782), .B2(new_n776), .ZN(new_n877));
  AOI221_X4 g691(.A(KEYINPUT110), .B1(new_n770), .B2(new_n775), .C1(new_n781), .C2(new_n774), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n871), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n863), .A2(new_n879), .A3(KEYINPUT53), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n875), .B1(new_n880), .B2(new_n861), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n876), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n747), .A2(new_n749), .ZN(new_n883));
  INV_X1    g697(.A(new_n424), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n801), .A2(new_n884), .A3(new_n803), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n885), .A2(KEYINPUT116), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(KEYINPUT116), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n883), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n728), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n718), .A2(new_n761), .ZN(new_n890));
  NOR4_X1   g704(.A1(new_n890), .A2(new_n701), .A3(new_n613), .A4(new_n424), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n891), .A2(new_n689), .A3(new_n708), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n889), .A2(new_n422), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n890), .B1(new_n886), .B2(new_n887), .ZN(new_n894));
  INV_X1    g708(.A(new_n773), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n896), .A2(KEYINPUT48), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(KEYINPUT48), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n893), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n717), .A2(new_n288), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n900), .A2(new_n301), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n901), .B1(new_n814), .B2(new_n816), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n888), .A2(new_n761), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n756), .A2(new_n757), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n708), .A2(new_n689), .ZN(new_n906));
  AOI22_X1  g720(.A1(new_n894), .A2(new_n905), .B1(new_n891), .B2(new_n906), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n686), .A2(new_n432), .A3(new_n718), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n888), .A2(KEYINPUT50), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT50), .B1(new_n888), .B2(new_n908), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n907), .B(KEYINPUT51), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n899), .B1(new_n904), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT118), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT117), .B1(new_n902), .B2(new_n903), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT117), .ZN(new_n917));
  INV_X1    g731(.A(new_n903), .ZN(new_n918));
  INV_X1    g732(.A(new_n816), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n799), .A2(new_n813), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n917), .B(new_n918), .C1(new_n921), .C2(new_n901), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n907), .B(KEYINPUT118), .C1(new_n909), .C2(new_n910), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n915), .A2(new_n916), .A3(new_n922), .A4(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT51), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n912), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n820), .B1(new_n882), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n642), .A2(new_n689), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n300), .A2(new_n432), .ZN(new_n929));
  AND4_X1   g743(.A1(new_n614), .A2(new_n686), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n701), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n900), .B(KEYINPUT49), .Z(new_n932));
  NAND3_X1  g746(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(KEYINPUT119), .B1(new_n927), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n880), .A2(new_n861), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(KEYINPUT54), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n861), .A2(new_n874), .A3(new_n875), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n926), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n820), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT119), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n941), .A2(new_n942), .A3(new_n933), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n935), .A2(new_n943), .ZN(G75));
  NOR2_X1   g758(.A1(new_n305), .A2(G952), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n861), .A2(new_n874), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n947), .A2(new_n280), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT56), .B1(new_n948), .B2(G210), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n473), .A2(new_n475), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(new_n487), .ZN(new_n951));
  XNOR2_X1  g765(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n951), .B(new_n952), .Z(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n946), .B1(new_n949), .B2(new_n954), .ZN(new_n955));
  AOI211_X1 g769(.A(KEYINPUT56), .B(new_n953), .C1(new_n948), .C2(G210), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n955), .A2(new_n956), .ZN(G51));
  NAND2_X1  g771(.A1(new_n861), .A2(new_n874), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(KEYINPUT54), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n938), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n289), .B(KEYINPUT57), .Z(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(new_n287), .B2(new_n284), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n794), .B(KEYINPUT121), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n948), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n945), .B1(new_n963), .B2(new_n965), .ZN(G54));
  NAND2_X1  g780(.A1(KEYINPUT58), .A2(G475), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n948), .A2(KEYINPUT122), .A3(new_n356), .A4(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT122), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n958), .A2(G902), .A3(new_n968), .ZN(new_n971));
  INV_X1    g785(.A(new_n356), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n945), .B1(new_n971), .B2(new_n972), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n969), .A2(new_n973), .A3(new_n974), .ZN(G60));
  INV_X1    g789(.A(new_n636), .ZN(new_n976));
  NAND2_X1  g790(.A1(G478), .A2(G902), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT59), .Z(new_n978));
  OAI21_X1  g792(.A(new_n976), .B1(new_n882), .B2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n978), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n960), .A2(new_n636), .A3(new_n980), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n979), .A2(new_n946), .A3(new_n981), .ZN(G63));
  NAND2_X1  g796(.A1(new_n661), .A2(new_n662), .ZN(new_n983));
  NAND2_X1  g797(.A1(G217), .A2(G902), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT60), .ZN(new_n985));
  OR3_X1    g799(.A1(new_n947), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n600), .B1(new_n947), .B2(new_n985), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n986), .A2(new_n946), .A3(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT61), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n986), .A2(KEYINPUT61), .A3(new_n946), .A4(new_n987), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n991), .ZN(G66));
  NAND2_X1  g806(.A1(new_n426), .A2(new_n481), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(G953), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n994), .B1(new_n859), .B2(G953), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n950), .B1(G898), .B2(new_n305), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n995), .B(new_n996), .ZN(G69));
  OAI21_X1  g811(.A(G953), .B1(new_n188), .B2(new_n670), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(new_n734), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n800), .A2(new_n1000), .A3(new_n895), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n839), .A2(new_n759), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n1002), .A2(new_n787), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n818), .A2(new_n1001), .A3(new_n1003), .A4(new_n811), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n305), .B1(new_n1004), .B2(new_n785), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n515), .A2(new_n516), .ZN(new_n1006));
  XOR2_X1   g820(.A(new_n348), .B(KEYINPUT123), .Z(new_n1007));
  XNOR2_X1  g821(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  OAI211_X1 g822(.A(new_n1005), .B(new_n1008), .C1(G900), .C2(new_n305), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT124), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n780), .A2(new_n303), .A3(new_n692), .A4(new_n848), .ZN(new_n1011));
  AND2_X1   g825(.A1(new_n811), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1002), .A2(new_n702), .ZN(new_n1013));
  OR2_X1    g827(.A1(new_n1013), .A2(KEYINPUT62), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1013), .A2(KEYINPUT62), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n1012), .A2(new_n818), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1008), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n1016), .A2(new_n305), .A3(new_n1017), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1009), .A2(new_n1010), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1010), .B1(new_n1009), .B2(new_n1018), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n999), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g836(.A(new_n1021), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1023), .A2(new_n998), .A3(new_n1019), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1022), .A2(new_n1024), .ZN(G72));
  NOR2_X1   g839(.A1(new_n545), .A2(new_n524), .ZN(new_n1026));
  NOR3_X1   g840(.A1(new_n1004), .A2(new_n785), .A3(new_n871), .ZN(new_n1027));
  NAND2_X1  g841(.A1(G472), .A2(G902), .ZN(new_n1028));
  XOR2_X1   g842(.A(new_n1028), .B(KEYINPUT63), .Z(new_n1029));
  INV_X1    g843(.A(new_n1029), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1026), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n1029), .B1(new_n1016), .B2(new_n871), .ZN(new_n1032));
  INV_X1    g846(.A(KEYINPUT125), .ZN(new_n1033));
  NOR2_X1   g847(.A1(new_n546), .A2(new_n523), .ZN(new_n1034));
  AND3_X1   g848(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1033), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1036));
  OAI211_X1 g850(.A(new_n946), .B(new_n1031), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  NOR3_X1   g851(.A1(new_n1034), .A2(new_n1030), .A3(new_n1026), .ZN(new_n1038));
  AND2_X1   g852(.A1(new_n936), .A2(new_n1038), .ZN(new_n1039));
  OR2_X1    g853(.A1(new_n1039), .A2(KEYINPUT126), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1039), .A2(KEYINPUT126), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n1037), .B1(new_n1040), .B2(new_n1041), .ZN(G57));
endmodule


