//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 1 0 0 0 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 0 0 1 0 1 1 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n544,
    new_n545, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT66), .Z(G259));
  XOR2_X1   g020(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(G125), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI211_X1 g040(.A(G137), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n460), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n465), .A2(new_n469), .ZN(G160));
  OR2_X1    g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(G2105), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G136), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n460), .B1(new_n471), .B2(new_n472), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  OR2_X1    g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n477), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n474), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G162));
  OAI21_X1  g055(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G114), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(new_n482), .B2(G2105), .ZN(new_n483));
  AND2_X1   g058(.A1(G126), .A2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n484), .B1(new_n461), .B2(new_n462), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT68), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(new_n484), .C1(new_n461), .C2(new_n462), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n483), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  OAI211_X1 g064(.A(G138), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  XNOR2_X1  g066(.A(KEYINPUT3), .B(G2104), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n492), .A2(new_n493), .A3(G138), .A4(new_n460), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n489), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  INV_X1    g072(.A(G651), .ZN(new_n498));
  XNOR2_X1  g073(.A(KEYINPUT5), .B(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G62), .ZN(new_n500));
  NAND2_X1  g075(.A1(G75), .A2(G543), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OR2_X1    g077(.A1(new_n502), .A2(KEYINPUT69), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(KEYINPUT69), .ZN(new_n504));
  XOR2_X1   g079(.A(KEYINPUT5), .B(G543), .Z(new_n505));
  AND2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n509), .A2(G88), .B1(new_n511), .B2(G50), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n503), .A2(new_n504), .A3(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(G166));
  NAND3_X1  g089(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n515), .B(KEYINPUT7), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G51), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n516), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n517), .A2(G89), .ZN(new_n521));
  NAND2_X1  g096(.A1(G63), .A2(G651), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n505), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OR3_X1    g098(.A1(new_n520), .A2(new_n523), .A3(KEYINPUT70), .ZN(new_n524));
  OAI21_X1  g099(.A(KEYINPUT70), .B1(new_n520), .B2(new_n523), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(G168));
  NAND2_X1  g101(.A1(new_n499), .A2(new_n517), .ZN(new_n527));
  INV_X1    g102(.A(G90), .ZN(new_n528));
  INV_X1    g103(.A(G52), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n527), .A2(new_n528), .B1(new_n518), .B2(new_n529), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n499), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n531), .A2(new_n498), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n530), .A2(new_n532), .ZN(G301));
  INV_X1    g108(.A(G301), .ZN(G171));
  INV_X1    g109(.A(G81), .ZN(new_n535));
  INV_X1    g110(.A(G43), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n527), .A2(new_n535), .B1(new_n518), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n499), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n498), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  NAND4_X1  g117(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g118(.A1(G1), .A2(G3), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT8), .ZN(new_n545));
  NAND4_X1  g120(.A1(G319), .A2(G483), .A3(G661), .A4(new_n545), .ZN(G188));
  AOI22_X1  g121(.A1(new_n499), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G91), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n547), .A2(new_n498), .B1(new_n527), .B2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  AND2_X1   g125(.A1(KEYINPUT71), .A2(G53), .ZN(new_n551));
  OAI211_X1 g126(.A(G543), .B(new_n551), .C1(new_n506), .C2(new_n507), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(KEYINPUT9), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT9), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n517), .A2(new_n554), .A3(G543), .A4(new_n551), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n556), .A2(KEYINPUT72), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT72), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n558), .B1(new_n553), .B2(new_n555), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n550), .B1(new_n557), .B2(new_n559), .ZN(G299));
  INV_X1    g135(.A(G168), .ZN(G286));
  INV_X1    g136(.A(KEYINPUT73), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n512), .B1(KEYINPUT69), .B2(new_n502), .ZN(new_n563));
  INV_X1    g138(.A(new_n504), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n503), .A2(KEYINPUT73), .A3(new_n512), .A4(new_n504), .ZN(new_n566));
  AND2_X1   g141(.A1(new_n565), .A2(new_n566), .ZN(G303));
  NAND3_X1  g142(.A1(new_n517), .A2(G49), .A3(G543), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT74), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n568), .B(new_n569), .ZN(new_n570));
  OR2_X1    g145(.A1(new_n499), .A2(G74), .ZN(new_n571));
  AOI22_X1  g146(.A1(G651), .A2(new_n571), .B1(new_n509), .B2(G87), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(G288));
  INV_X1    g148(.A(G86), .ZN(new_n574));
  INV_X1    g149(.A(G48), .ZN(new_n575));
  OAI22_X1  g150(.A1(new_n527), .A2(new_n574), .B1(new_n518), .B2(new_n575), .ZN(new_n576));
  AND2_X1   g151(.A1(G73), .A2(G543), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n577), .B1(new_n499), .B2(G61), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n578), .A2(new_n498), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G305));
  AND2_X1   g156(.A1(new_n499), .A2(G60), .ZN(new_n582));
  AND2_X1   g157(.A1(G72), .A2(G543), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT75), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n585), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n509), .A2(G85), .B1(new_n511), .B2(G47), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n509), .A2(KEYINPUT10), .A3(G92), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n592));
  INV_X1    g167(.A(G92), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n527), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G66), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n505), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n598), .A2(G651), .B1(new_n511), .B2(G54), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n590), .B1(new_n601), .B2(G868), .ZN(G284));
  OAI21_X1  g177(.A(new_n590), .B1(new_n601), .B2(G868), .ZN(G321));
  NOR2_X1   g178(.A1(G299), .A2(G868), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n604), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g180(.A(new_n604), .B1(G868), .B2(G168), .ZN(G280));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n601), .B1(new_n607), .B2(G860), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT76), .ZN(G148));
  NAND2_X1  g184(.A1(new_n601), .A2(new_n607), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  OR3_X1    g187(.A1(new_n611), .A2(KEYINPUT77), .A3(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(KEYINPUT77), .B1(new_n611), .B2(new_n612), .ZN(new_n614));
  OAI211_X1 g189(.A(new_n613), .B(new_n614), .C1(G868), .C2(new_n541), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g191(.A1(new_n475), .A2(G123), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT80), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n473), .A2(G135), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT79), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n460), .A2(G111), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n618), .B(new_n620), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT81), .Z(new_n624));
  OR2_X1    g199(.A1(new_n624), .A2(G2096), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(G2096), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n492), .A2(new_n467), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT12), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2100), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT78), .B(KEYINPUT13), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n625), .A2(new_n626), .A3(new_n631), .ZN(G156));
  INV_X1    g207(.A(KEYINPUT14), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2427), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(new_n636), .B2(new_n635), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n638), .B(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(G14), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n647), .B1(new_n646), .B2(new_n644), .ZN(G401));
  XOR2_X1   g223(.A(G2067), .B(G2678), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT82), .ZN(new_n650));
  NOR2_X1   g225(.A1(G2072), .A2(G2078), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n442), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  NOR3_X1   g229(.A1(new_n650), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT18), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n652), .A2(KEYINPUT83), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n652), .A2(KEYINPUT83), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n650), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n652), .B(KEYINPUT17), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n659), .B(new_n654), .C1(new_n650), .C2(new_n660), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n650), .A2(new_n653), .A3(new_n660), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n656), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2096), .B(G2100), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(G227));
  XNOR2_X1  g240(.A(G1961), .B(G1966), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT85), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1956), .B(G2474), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n670), .A2(new_n671), .A3(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT86), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n675), .B1(new_n670), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n678), .B1(new_n677), .B2(new_n670), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n679), .A2(KEYINPUT20), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n679), .A2(KEYINPUT20), .ZN(new_n681));
  OAI221_X1 g256(.A(new_n676), .B1(new_n675), .B2(new_n671), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1991), .B(G1996), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1981), .B(G1986), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT87), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n684), .B(new_n688), .ZN(G229));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G23), .ZN(new_n691));
  INV_X1    g266(.A(G288), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(new_n690), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT90), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT33), .B(G1976), .Z(new_n695));
  XOR2_X1   g270(.A(new_n694), .B(new_n695), .Z(new_n696));
  NAND2_X1  g271(.A1(G166), .A2(G16), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G16), .B2(G22), .ZN(new_n698));
  INV_X1    g273(.A(G1971), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(G6), .A2(G16), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(new_n580), .B2(G16), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT32), .B(G1981), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n698), .A2(new_n699), .ZN(new_n705));
  NAND4_X1  g280(.A1(new_n696), .A2(new_n700), .A3(new_n704), .A4(new_n705), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n706), .A2(KEYINPUT34), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(KEYINPUT34), .ZN(new_n708));
  OR2_X1    g283(.A1(G16), .A2(G24), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G290), .B2(new_n690), .ZN(new_n710));
  INV_X1    g285(.A(G1986), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G25), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT88), .Z(new_n716));
  NAND2_X1  g291(.A1(new_n473), .A2(G131), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n475), .A2(G119), .ZN(new_n718));
  OR2_X1    g293(.A1(G95), .A2(G2105), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n719), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n716), .B1(new_n721), .B2(G29), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT35), .B(G1991), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT89), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(KEYINPUT91), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n725), .B2(new_n722), .ZN(new_n727));
  AND3_X1   g302(.A1(new_n712), .A2(new_n713), .A3(new_n727), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n707), .A2(new_n708), .A3(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT36), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n714), .A2(G35), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G162), .B2(new_n714), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT29), .ZN(new_n734));
  OAI22_X1  g309(.A1(new_n624), .A2(new_n714), .B1(G2090), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n690), .A2(G21), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G168), .B2(new_n690), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n735), .B1(G1966), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n734), .A2(G2090), .ZN(new_n739));
  NOR2_X1   g314(.A1(G4), .A2(G16), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT92), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n600), .B2(new_n690), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G1348), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n714), .A2(G32), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n475), .A2(G129), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT96), .Z(new_n746));
  NAND3_X1  g321(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT98), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT26), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n467), .A2(G105), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n750), .A2(KEYINPUT97), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(KEYINPUT97), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n751), .A2(new_n752), .B1(G141), .B2(new_n473), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n746), .A2(new_n749), .A3(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n744), .B1(new_n755), .B2(new_n714), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT27), .B(G1996), .Z(new_n757));
  XOR2_X1   g332(.A(new_n756), .B(new_n757), .Z(new_n758));
  AND4_X1   g333(.A1(new_n738), .A2(new_n739), .A3(new_n743), .A4(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(G16), .A2(G19), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n541), .B2(G16), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT93), .B(G1341), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT25), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n492), .A2(G127), .ZN(new_n766));
  NAND2_X1  g341(.A1(G115), .A2(G2104), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n460), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AOI211_X1 g343(.A(new_n765), .B(new_n768), .C1(G139), .C2(new_n473), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n769), .A2(new_n714), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n714), .A2(G33), .ZN(new_n771));
  OR3_X1    g346(.A1(new_n770), .A2(G2072), .A3(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(G2072), .B1(new_n770), .B2(new_n771), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT24), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n714), .B1(new_n774), .B2(G34), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n774), .B2(G34), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G160), .B2(G29), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n772), .B(new_n773), .C1(G2084), .C2(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(G5), .A2(G16), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT100), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G301), .B2(new_n690), .ZN(new_n781));
  INV_X1    g356(.A(G1961), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n777), .A2(G2084), .ZN(new_n784));
  NOR2_X1   g359(.A1(KEYINPUT31), .A2(G11), .ZN(new_n785));
  AND2_X1   g360(.A1(KEYINPUT31), .A2(G11), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT30), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n787), .A2(G28), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n714), .B1(new_n787), .B2(G28), .ZN(new_n789));
  OAI221_X1 g364(.A(new_n784), .B1(new_n785), .B2(new_n786), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  NOR3_X1   g365(.A1(new_n778), .A2(new_n783), .A3(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(G27), .A2(G29), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G164), .B2(G29), .ZN(new_n793));
  INV_X1    g368(.A(G2078), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n737), .A2(G1966), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT99), .Z(new_n797));
  AND4_X1   g372(.A1(new_n763), .A2(new_n791), .A3(new_n795), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n690), .A2(G20), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT23), .ZN(new_n800));
  INV_X1    g375(.A(G299), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(new_n690), .ZN(new_n802));
  INV_X1    g377(.A(G1956), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n473), .A2(G140), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT94), .ZN(new_n806));
  OAI21_X1  g381(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n807));
  INV_X1    g382(.A(G116), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(G2105), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n475), .B2(G128), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(G29), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT95), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n714), .A2(G26), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT28), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(G2067), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n759), .A2(new_n798), .A3(new_n804), .A4(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT101), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n729), .A2(new_n730), .ZN(new_n822));
  AND3_X1   g397(.A1(new_n731), .A2(new_n821), .A3(new_n822), .ZN(G311));
  NAND3_X1  g398(.A1(new_n731), .A2(new_n821), .A3(new_n822), .ZN(G150));
  AOI22_X1  g399(.A1(new_n509), .A2(G93), .B1(new_n511), .B2(G55), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n499), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n498), .B2(new_n826), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT103), .B(G860), .Z(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT37), .Z(new_n831));
  NAND2_X1  g406(.A1(new_n601), .A2(G559), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT38), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n540), .B(new_n827), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT39), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT102), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n828), .B1(new_n835), .B2(new_n836), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n831), .B1(new_n838), .B2(new_n839), .ZN(G145));
  XOR2_X1   g415(.A(new_n624), .B(G160), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(G162), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n473), .A2(G142), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n460), .A2(G118), .ZN(new_n845));
  OAI21_X1  g420(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n846));
  AND3_X1   g421(.A1(new_n475), .A2(KEYINPUT105), .A3(G130), .ZN(new_n847));
  AOI21_X1  g422(.A(KEYINPUT105), .B1(new_n475), .B2(G130), .ZN(new_n848));
  OAI221_X1 g423(.A(new_n844), .B1(new_n845), .B2(new_n846), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT106), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n628), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n851), .A2(new_n721), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n721), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n811), .B(G164), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n754), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n769), .A2(KEYINPUT104), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n769), .A2(KEYINPUT104), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n856), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n854), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n854), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n858), .A2(new_n860), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n862), .B1(KEYINPUT107), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT107), .ZN(new_n867));
  NOR3_X1   g442(.A1(new_n863), .A2(new_n864), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n843), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n842), .A2(new_n861), .A3(new_n865), .ZN(new_n870));
  INV_X1    g445(.A(G37), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  AND3_X1   g448(.A1(new_n869), .A2(new_n873), .A3(KEYINPUT40), .ZN(new_n874));
  AOI21_X1  g449(.A(KEYINPUT40), .B1(new_n869), .B2(new_n873), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(new_n875), .ZN(G395));
  NAND2_X1  g451(.A1(new_n827), .A2(new_n612), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n601), .B(G299), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT41), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n834), .B(new_n611), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n881), .B1(new_n878), .B2(new_n880), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT42), .ZN(new_n883));
  XNOR2_X1  g458(.A(G166), .B(G290), .ZN(new_n884));
  XNOR2_X1  g459(.A(G288), .B(new_n580), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n883), .B(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n877), .B1(new_n888), .B2(new_n612), .ZN(G295));
  OAI21_X1  g464(.A(new_n877), .B1(new_n888), .B2(new_n612), .ZN(G331));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n891));
  OR2_X1    g466(.A1(G168), .A2(KEYINPUT109), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n834), .ZN(new_n893));
  AOI21_X1  g468(.A(G301), .B1(G168), .B2(KEYINPUT109), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n894), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n879), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n895), .A2(new_n878), .A3(new_n896), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n886), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n901), .A2(G37), .ZN(new_n902));
  XOR2_X1   g477(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n903));
  NAND3_X1  g478(.A1(new_n899), .A2(new_n886), .A3(new_n900), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n903), .B1(new_n902), .B2(new_n904), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n891), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n908));
  INV_X1    g483(.A(new_n904), .ZN(new_n909));
  NOR3_X1   g484(.A1(new_n909), .A2(G37), .A3(new_n901), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n908), .B(KEYINPUT44), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n907), .A2(new_n912), .ZN(G397));
  AOI21_X1  g488(.A(G1384), .B1(new_n489), .B2(new_n495), .ZN(new_n914));
  XOR2_X1   g489(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(G40), .ZN(new_n918));
  NOR3_X1   g493(.A1(new_n465), .A2(new_n469), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G1996), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(KEYINPUT46), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n811), .B(new_n817), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n925), .A2(new_n755), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n924), .B1(new_n920), .B2(new_n926), .ZN(new_n927));
  XOR2_X1   g502(.A(new_n927), .B(KEYINPUT126), .Z(new_n928));
  OR2_X1    g503(.A1(new_n928), .A2(KEYINPUT47), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(KEYINPUT47), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n754), .B(new_n922), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n931), .A2(new_n925), .ZN(new_n932));
  INV_X1    g507(.A(new_n721), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n932), .A2(new_n725), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n806), .A2(new_n817), .A3(new_n810), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n920), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n725), .B(new_n721), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n932), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(new_n921), .ZN(new_n939));
  NOR3_X1   g514(.A1(new_n920), .A2(G1986), .A3(G290), .ZN(new_n940));
  XOR2_X1   g515(.A(new_n940), .B(KEYINPUT48), .Z(new_n941));
  AOI21_X1  g516(.A(new_n936), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n929), .A2(new_n930), .A3(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(G1981), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n580), .A2(new_n944), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n578), .A2(new_n498), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n509), .A2(G86), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n511), .A2(G48), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n946), .A2(new_n944), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT113), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n580), .A2(KEYINPUT113), .A3(new_n944), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n945), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n953), .A2(KEYINPUT49), .ZN(new_n954));
  INV_X1    g529(.A(G8), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n955), .B1(new_n914), .B2(new_n919), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n956), .B1(new_n953), .B2(KEYINPUT49), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(G288), .A2(G1976), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n959), .A2(new_n960), .B1(new_n951), .B2(new_n952), .ZN(new_n961));
  INV_X1    g536(.A(new_n956), .ZN(new_n962));
  INV_X1    g537(.A(G1384), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n496), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT112), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(new_n965), .A3(new_n915), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT112), .B1(new_n914), .B2(new_n916), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n463), .A2(new_n464), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(G2105), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n969), .A2(G40), .A3(new_n468), .A4(new_n466), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n970), .B1(new_n914), .B2(KEYINPUT45), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n966), .A2(new_n967), .A3(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n496), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT50), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n974), .B(new_n919), .C1(new_n975), .C2(new_n914), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G2090), .ZN(new_n978));
  AOI22_X1  g553(.A1(new_n972), .A2(new_n699), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n979), .A2(new_n955), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n565), .A2(G8), .A3(new_n566), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT55), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n981), .B(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n692), .A2(G1976), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n956), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT52), .ZN(new_n987));
  INV_X1    g562(.A(G1976), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT52), .B1(G288), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n985), .A2(new_n989), .A3(new_n956), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n987), .B(new_n990), .C1(new_n954), .C2(new_n957), .ZN(new_n991));
  OAI22_X1  g566(.A1(new_n961), .A2(new_n962), .B1(new_n984), .B2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n991), .B1(new_n983), .B2(new_n980), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT114), .B1(new_n980), .B2(new_n983), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n981), .B(KEYINPUT55), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n995), .B(new_n996), .C1(new_n955), .C2(new_n979), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n974), .A2(new_n919), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n975), .B1(new_n496), .B2(new_n963), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n998), .A2(G2084), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT45), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n964), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n915), .A2(G1384), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n970), .B1(new_n496), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(G1966), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(G8), .B1(new_n1000), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1006), .A2(G286), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n993), .A2(new_n994), .A3(new_n997), .A4(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT63), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n979), .A2(new_n955), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n995), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n993), .A2(KEYINPUT63), .A3(new_n1012), .A4(new_n1007), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n992), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G1966), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n496), .A2(new_n1003), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n919), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n914), .A2(KEYINPUT45), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1015), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT120), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n964), .A2(KEYINPUT50), .ZN(new_n1021));
  INV_X1    g596(.A(G2084), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n970), .B1(new_n496), .B2(new_n973), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1019), .A2(new_n1020), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1020), .B1(new_n1019), .B2(new_n1024), .ZN(new_n1026));
  NAND2_X1  g601(.A1(G286), .A2(G8), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1006), .A2(new_n1029), .A3(new_n1027), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT121), .B1(new_n1032), .B2(G8), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT120), .B1(new_n1000), .B2(new_n1005), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1019), .A2(new_n1020), .A3(new_n1024), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1034), .A2(KEYINPUT121), .A3(G8), .A4(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n1027), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT51), .B1(new_n1033), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT122), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1031), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI211_X1 g615(.A(KEYINPUT122), .B(KEYINPUT51), .C1(new_n1033), .C2(new_n1037), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1028), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT56), .B(G2072), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n966), .A2(new_n967), .A3(new_n971), .A4(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n803), .B1(new_n998), .B2(new_n999), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n553), .A2(new_n555), .ZN(new_n1047));
  NOR3_X1   g622(.A1(new_n549), .A2(new_n1047), .A3(KEYINPUT57), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1048), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1046), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n914), .A2(new_n817), .A3(new_n919), .ZN(new_n1053));
  INV_X1    g628(.A(G1348), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1053), .B1(new_n976), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1052), .B1(new_n1055), .B2(new_n600), .ZN(new_n1056));
  AOI21_X1  g631(.A(G1348), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1057));
  OAI211_X1 g632(.A(KEYINPUT116), .B(new_n601), .C1(new_n1057), .C2(new_n1053), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1051), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1044), .A2(new_n1049), .A3(new_n1045), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1044), .A2(new_n1045), .A3(KEYINPUT115), .A4(new_n1049), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1059), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT117), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1059), .A2(new_n1064), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT118), .B1(new_n1046), .B2(new_n1050), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n1070));
  AOI211_X1 g645(.A(new_n1070), .B(new_n1049), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT61), .B1(new_n1072), .B2(new_n1064), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n600), .A2(KEYINPUT119), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT119), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1075), .B1(new_n595), .B2(new_n599), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1055), .A2(KEYINPUT60), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT60), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1079), .B1(new_n1057), .B2(new_n1053), .ZN(new_n1080));
  NOR3_X1   g655(.A1(new_n1057), .A2(new_n1079), .A3(new_n1053), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1076), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1078), .B(new_n1080), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1051), .A2(KEYINPUT61), .A3(new_n1060), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n966), .A2(new_n967), .A3(new_n971), .A4(new_n922), .ZN(new_n1086));
  XOR2_X1   g661(.A(KEYINPUT58), .B(G1341), .Z(new_n1087));
  OAI21_X1  g662(.A(new_n1087), .B1(new_n964), .B2(new_n970), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1085), .B1(new_n1089), .B2(new_n541), .ZN(new_n1090));
  AOI211_X1 g665(.A(KEYINPUT59), .B(new_n540), .C1(new_n1086), .C2(new_n1088), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1083), .B(new_n1084), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1066), .B(new_n1068), .C1(new_n1073), .C2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT125), .ZN(new_n1094));
  INV_X1    g669(.A(new_n991), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n997), .A2(new_n984), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n996), .B1(new_n1011), .B2(new_n995), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1094), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n966), .A2(new_n967), .A3(new_n971), .A4(new_n794), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n782), .B1(new_n998), .B2(new_n999), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1100), .A2(G2078), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1002), .A2(new_n1004), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NOR3_X1   g680(.A1(new_n1101), .A2(G171), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1103), .B1(new_n919), .B2(KEYINPUT124), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1108), .B1(KEYINPUT124), .B2(new_n919), .ZN(new_n1109));
  AOI211_X1 g684(.A(new_n1001), .B(G1384), .C1(new_n489), .C2(new_n495), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n917), .A2(new_n1110), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n1109), .A2(new_n1111), .B1(new_n976), .B2(new_n782), .ZN(new_n1112));
  AOI21_X1  g687(.A(G301), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n1106), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1105), .B1(new_n1100), .B2(new_n1099), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1116), .B1(new_n1117), .B2(G301), .ZN(new_n1118));
  OAI211_X1 g693(.A(KEYINPUT123), .B(G171), .C1(new_n1101), .C2(new_n1105), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1107), .A2(new_n1112), .A3(G301), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1115), .B1(new_n1121), .B2(new_n1114), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n993), .A2(new_n994), .A3(KEYINPUT125), .A4(new_n997), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1093), .A2(new_n1098), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1014), .B1(new_n1042), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1098), .A2(new_n1123), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1028), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1036), .A2(new_n1027), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1034), .A2(G8), .A3(new_n1035), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1029), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1030), .B1(new_n1133), .B2(KEYINPUT122), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1041), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1128), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1127), .B1(new_n1136), .B2(KEYINPUT62), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1042), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1125), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(G290), .B(new_n711), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n939), .B1(new_n920), .B2(new_n1141), .ZN(new_n1142));
  XOR2_X1   g717(.A(new_n1142), .B(KEYINPUT111), .Z(new_n1143));
  OAI21_X1  g718(.A(new_n943), .B1(new_n1140), .B2(new_n1143), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g719(.A1(new_n905), .A2(new_n906), .ZN(new_n1146));
  INV_X1    g720(.A(G319), .ZN(new_n1147));
  NOR3_X1   g721(.A1(G401), .A2(new_n1147), .A3(G227), .ZN(new_n1148));
  XNOR2_X1  g722(.A(new_n1148), .B(KEYINPUT127), .ZN(new_n1149));
  NOR2_X1   g723(.A1(G229), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g724(.A1(new_n865), .A2(KEYINPUT107), .ZN(new_n1151));
  NAND2_X1  g725(.A1(new_n1151), .A2(new_n861), .ZN(new_n1152));
  INV_X1    g726(.A(new_n868), .ZN(new_n1153));
  AOI21_X1  g727(.A(new_n842), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g728(.A(new_n1150), .B1(new_n1154), .B2(new_n872), .ZN(new_n1155));
  NOR2_X1   g729(.A1(new_n1146), .A2(new_n1155), .ZN(G308));
  OAI221_X1 g730(.A(new_n1150), .B1(new_n1154), .B2(new_n872), .C1(new_n905), .C2(new_n906), .ZN(G225));
endmodule


