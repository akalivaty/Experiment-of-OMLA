

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591;

  XNOR2_X1 U326 ( .A(n412), .B(n411), .ZN(n573) );
  XNOR2_X1 U327 ( .A(n410), .B(KEYINPUT119), .ZN(n411) );
  XNOR2_X1 U328 ( .A(n309), .B(n308), .ZN(n533) );
  XNOR2_X1 U329 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U330 ( .A(n359), .B(n358), .ZN(n360) );
  NOR2_X1 U331 ( .A1(n533), .A2(n453), .ZN(n567) );
  XNOR2_X1 U332 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U333 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  XOR2_X1 U334 ( .A(G183GAT), .B(G176GAT), .Z(n295) );
  XNOR2_X1 U335 ( .A(G190GAT), .B(G99GAT), .ZN(n294) );
  XNOR2_X1 U336 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U337 ( .A(KEYINPUT20), .B(KEYINPUT81), .Z(n297) );
  XNOR2_X1 U338 ( .A(G169GAT), .B(KEYINPUT80), .ZN(n296) );
  XNOR2_X1 U339 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U340 ( .A(n299), .B(n298), .ZN(n309) );
  XNOR2_X1 U341 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n300) );
  XNOR2_X1 U342 ( .A(n300), .B(KEYINPUT17), .ZN(n326) );
  XOR2_X1 U343 ( .A(n326), .B(KEYINPUT82), .Z(n302) );
  NAND2_X1 U344 ( .A1(G227GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U345 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U346 ( .A(G113GAT), .B(KEYINPUT0), .Z(n432) );
  XNOR2_X1 U347 ( .A(n303), .B(n432), .ZN(n307) );
  XOR2_X1 U348 ( .A(G120GAT), .B(G71GAT), .Z(n356) );
  XOR2_X1 U349 ( .A(G134GAT), .B(n356), .Z(n305) );
  XOR2_X1 U350 ( .A(G15GAT), .B(G127GAT), .Z(n370) );
  XNOR2_X1 U351 ( .A(G43GAT), .B(n370), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U353 ( .A(n307), .B(n306), .ZN(n308) );
  INV_X1 U354 ( .A(G92GAT), .ZN(n310) );
  NAND2_X1 U355 ( .A1(G64GAT), .A2(n310), .ZN(n313) );
  INV_X1 U356 ( .A(G64GAT), .ZN(n311) );
  NAND2_X1 U357 ( .A1(n311), .A2(G92GAT), .ZN(n312) );
  NAND2_X1 U358 ( .A1(n313), .A2(n312), .ZN(n315) );
  XNOR2_X1 U359 ( .A(G176GAT), .B(G204GAT), .ZN(n314) );
  XNOR2_X1 U360 ( .A(n315), .B(n314), .ZN(n352) );
  XOR2_X1 U361 ( .A(G169GAT), .B(G8GAT), .Z(n338) );
  XOR2_X1 U362 ( .A(n352), .B(n338), .Z(n317) );
  NAND2_X1 U363 ( .A1(G226GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U364 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U365 ( .A(n318), .B(KEYINPUT90), .Z(n320) );
  XOR2_X1 U366 ( .A(G183GAT), .B(KEYINPUT76), .Z(n362) );
  XNOR2_X1 U367 ( .A(n362), .B(KEYINPUT89), .ZN(n319) );
  XNOR2_X1 U368 ( .A(n320), .B(n319), .ZN(n322) );
  XNOR2_X1 U369 ( .A(G36GAT), .B(G190GAT), .ZN(n321) );
  XNOR2_X1 U370 ( .A(n321), .B(KEYINPUT75), .ZN(n398) );
  XOR2_X1 U371 ( .A(n322), .B(n398), .Z(n328) );
  XOR2_X1 U372 ( .A(KEYINPUT83), .B(G218GAT), .Z(n324) );
  XNOR2_X1 U373 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n323) );
  XNOR2_X1 U374 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U375 ( .A(G197GAT), .B(n325), .Z(n427) );
  XNOR2_X1 U376 ( .A(n326), .B(n427), .ZN(n327) );
  XNOR2_X1 U377 ( .A(n328), .B(n327), .ZN(n519) );
  XOR2_X1 U378 ( .A(G1GAT), .B(G15GAT), .Z(n330) );
  XNOR2_X1 U379 ( .A(G197GAT), .B(G113GAT), .ZN(n329) );
  XNOR2_X1 U380 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U381 ( .A(KEYINPUT68), .B(KEYINPUT29), .Z(n332) );
  XNOR2_X1 U382 ( .A(KEYINPUT66), .B(KEYINPUT67), .ZN(n331) );
  XNOR2_X1 U383 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U384 ( .A(n334), .B(n333), .ZN(n347) );
  XOR2_X1 U385 ( .A(G22GAT), .B(G141GAT), .Z(n336) );
  XNOR2_X1 U386 ( .A(G50GAT), .B(G36GAT), .ZN(n335) );
  XNOR2_X1 U387 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U388 ( .A(n338), .B(n337), .Z(n340) );
  NAND2_X1 U389 ( .A1(G229GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U390 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U391 ( .A(n341), .B(KEYINPUT30), .Z(n345) );
  XOR2_X1 U392 ( .A(G29GAT), .B(G43GAT), .Z(n343) );
  XNOR2_X1 U393 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n342) );
  XNOR2_X1 U394 ( .A(n343), .B(n342), .ZN(n386) );
  XNOR2_X1 U395 ( .A(n386), .B(KEYINPUT69), .ZN(n344) );
  XNOR2_X1 U396 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U397 ( .A(n347), .B(n346), .ZN(n575) );
  XNOR2_X1 U398 ( .A(KEYINPUT70), .B(KEYINPUT33), .ZN(n349) );
  AND2_X1 U399 ( .A1(G230GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U400 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U401 ( .A(n350), .B(KEYINPUT32), .Z(n354) );
  XNOR2_X1 U402 ( .A(G106GAT), .B(G78GAT), .ZN(n351) );
  XNOR2_X1 U403 ( .A(n351), .B(G148GAT), .ZN(n421) );
  XNOR2_X1 U404 ( .A(n352), .B(n421), .ZN(n353) );
  XNOR2_X1 U405 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U406 ( .A(n355), .B(KEYINPUT31), .ZN(n359) );
  XOR2_X1 U407 ( .A(KEYINPUT13), .B(G57GAT), .Z(n363) );
  XOR2_X1 U408 ( .A(n363), .B(KEYINPUT71), .Z(n357) );
  XOR2_X1 U409 ( .A(G99GAT), .B(G85GAT), .Z(n383) );
  XNOR2_X1 U410 ( .A(n360), .B(n383), .ZN(n580) );
  XOR2_X1 U411 ( .A(KEYINPUT41), .B(n580), .Z(n553) );
  NAND2_X1 U412 ( .A1(n575), .A2(n553), .ZN(n361) );
  XNOR2_X1 U413 ( .A(n361), .B(KEYINPUT46), .ZN(n381) );
  XOR2_X1 U414 ( .A(n363), .B(n362), .Z(n365) );
  XNOR2_X1 U415 ( .A(G211GAT), .B(G78GAT), .ZN(n364) );
  XNOR2_X1 U416 ( .A(n365), .B(n364), .ZN(n369) );
  XOR2_X1 U417 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n367) );
  NAND2_X1 U418 ( .A1(G231GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U419 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U420 ( .A(n369), .B(n368), .Z(n372) );
  XOR2_X1 U421 ( .A(G22GAT), .B(G155GAT), .Z(n415) );
  XNOR2_X1 U422 ( .A(n370), .B(n415), .ZN(n371) );
  XNOR2_X1 U423 ( .A(n372), .B(n371), .ZN(n380) );
  XOR2_X1 U424 ( .A(KEYINPUT12), .B(G64GAT), .Z(n374) );
  XNOR2_X1 U425 ( .A(G8GAT), .B(G71GAT), .ZN(n373) );
  XNOR2_X1 U426 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U427 ( .A(KEYINPUT15), .B(KEYINPUT77), .Z(n376) );
  XNOR2_X1 U428 ( .A(G1GAT), .B(KEYINPUT14), .ZN(n375) );
  XNOR2_X1 U429 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U430 ( .A(n378), .B(n377), .Z(n379) );
  XNOR2_X1 U431 ( .A(n380), .B(n379), .ZN(n477) );
  NAND2_X1 U432 ( .A1(n381), .A2(n477), .ZN(n382) );
  XNOR2_X1 U433 ( .A(n382), .B(KEYINPUT107), .ZN(n401) );
  XOR2_X1 U434 ( .A(KEYINPUT65), .B(KEYINPUT64), .Z(n385) );
  XOR2_X1 U435 ( .A(G134GAT), .B(KEYINPUT74), .Z(n431) );
  XNOR2_X1 U436 ( .A(n383), .B(n431), .ZN(n384) );
  XNOR2_X1 U437 ( .A(n385), .B(n384), .ZN(n390) );
  XOR2_X1 U438 ( .A(n386), .B(KEYINPUT11), .Z(n388) );
  NAND2_X1 U439 ( .A1(G232GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U440 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U441 ( .A(n390), .B(n389), .Z(n392) );
  XNOR2_X1 U442 ( .A(G218GAT), .B(G92GAT), .ZN(n391) );
  XNOR2_X1 U443 ( .A(n392), .B(n391), .ZN(n396) );
  XOR2_X1 U444 ( .A(KEYINPUT73), .B(KEYINPUT10), .Z(n394) );
  XNOR2_X1 U445 ( .A(G106GAT), .B(KEYINPUT9), .ZN(n393) );
  XNOR2_X1 U446 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U447 ( .A(n396), .B(n395), .Z(n400) );
  XNOR2_X1 U448 ( .A(G50GAT), .B(KEYINPUT72), .ZN(n397) );
  XNOR2_X1 U449 ( .A(n397), .B(G162GAT), .ZN(n422) );
  XNOR2_X1 U450 ( .A(n422), .B(n398), .ZN(n399) );
  XNOR2_X1 U451 ( .A(n400), .B(n399), .ZN(n454) );
  NAND2_X1 U452 ( .A1(n401), .A2(n454), .ZN(n402) );
  XNOR2_X1 U453 ( .A(n402), .B(KEYINPUT47), .ZN(n408) );
  XOR2_X1 U454 ( .A(KEYINPUT45), .B(KEYINPUT108), .Z(n404) );
  INV_X1 U455 ( .A(n477), .ZN(n585) );
  XOR2_X1 U456 ( .A(KEYINPUT36), .B(n454), .Z(n587) );
  NAND2_X1 U457 ( .A1(n585), .A2(n587), .ZN(n403) );
  XNOR2_X1 U458 ( .A(n404), .B(n403), .ZN(n405) );
  INV_X1 U459 ( .A(n575), .ZN(n550) );
  NAND2_X1 U460 ( .A1(n405), .A2(n550), .ZN(n406) );
  NOR2_X1 U461 ( .A1(n580), .A2(n406), .ZN(n407) );
  NOR2_X1 U462 ( .A1(n408), .A2(n407), .ZN(n409) );
  XNOR2_X1 U463 ( .A(n409), .B(KEYINPUT48), .ZN(n529) );
  NOR2_X1 U464 ( .A1(n519), .A2(n529), .ZN(n412) );
  INV_X1 U465 ( .A(KEYINPUT54), .ZN(n410) );
  XOR2_X1 U466 ( .A(KEYINPUT24), .B(KEYINPUT85), .Z(n417) );
  XOR2_X1 U467 ( .A(KEYINPUT2), .B(KEYINPUT84), .Z(n414) );
  XNOR2_X1 U468 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n413) );
  XNOR2_X1 U469 ( .A(n414), .B(n413), .ZN(n440) );
  XNOR2_X1 U470 ( .A(n440), .B(n415), .ZN(n416) );
  XNOR2_X1 U471 ( .A(n417), .B(n416), .ZN(n426) );
  XOR2_X1 U472 ( .A(KEYINPUT23), .B(G204GAT), .Z(n419) );
  NAND2_X1 U473 ( .A1(G228GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U474 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U475 ( .A(n420), .B(KEYINPUT22), .Z(n424) );
  XNOR2_X1 U476 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U477 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U478 ( .A(n426), .B(n425), .ZN(n428) );
  XOR2_X1 U479 ( .A(n428), .B(n427), .Z(n472) );
  XOR2_X1 U480 ( .A(KEYINPUT1), .B(KEYINPUT87), .Z(n430) );
  XNOR2_X1 U481 ( .A(KEYINPUT88), .B(KEYINPUT4), .ZN(n429) );
  XNOR2_X1 U482 ( .A(n430), .B(n429), .ZN(n436) );
  XOR2_X1 U483 ( .A(n431), .B(G162GAT), .Z(n434) );
  XNOR2_X1 U484 ( .A(G29GAT), .B(n432), .ZN(n433) );
  XNOR2_X1 U485 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U486 ( .A(n436), .B(n435), .Z(n438) );
  NAND2_X1 U487 ( .A1(G225GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U488 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U489 ( .A(n439), .B(KEYINPUT86), .Z(n442) );
  XNOR2_X1 U490 ( .A(n440), .B(KEYINPUT6), .ZN(n441) );
  XNOR2_X1 U491 ( .A(n442), .B(n441), .ZN(n450) );
  XOR2_X1 U492 ( .A(KEYINPUT5), .B(G57GAT), .Z(n444) );
  XNOR2_X1 U493 ( .A(G1GAT), .B(G120GAT), .ZN(n443) );
  XNOR2_X1 U494 ( .A(n444), .B(n443), .ZN(n448) );
  XOR2_X1 U495 ( .A(G85GAT), .B(G155GAT), .Z(n446) );
  XNOR2_X1 U496 ( .A(G127GAT), .B(G148GAT), .ZN(n445) );
  XNOR2_X1 U497 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U498 ( .A(n448), .B(n447), .Z(n449) );
  XNOR2_X1 U499 ( .A(n450), .B(n449), .ZN(n517) );
  INV_X1 U500 ( .A(n517), .ZN(n570) );
  NOR2_X1 U501 ( .A1(n472), .A2(n570), .ZN(n451) );
  AND2_X1 U502 ( .A1(n573), .A2(n451), .ZN(n452) );
  XNOR2_X1 U503 ( .A(n452), .B(KEYINPUT55), .ZN(n453) );
  INV_X1 U504 ( .A(n454), .ZN(n563) );
  NAND2_X1 U505 ( .A1(n567), .A2(n563), .ZN(n458) );
  XOR2_X1 U506 ( .A(KEYINPUT58), .B(KEYINPUT122), .Z(n456) );
  INV_X1 U507 ( .A(G190GAT), .ZN(n455) );
  XNOR2_X1 U508 ( .A(n553), .B(KEYINPUT100), .ZN(n535) );
  NAND2_X1 U509 ( .A1(n567), .A2(n535), .ZN(n461) );
  XOR2_X1 U510 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n459) );
  XNOR2_X1 U511 ( .A(n459), .B(G176GAT), .ZN(n460) );
  XNOR2_X1 U512 ( .A(n461), .B(n460), .ZN(G1349GAT) );
  NOR2_X1 U513 ( .A1(n580), .A2(n550), .ZN(n493) );
  NOR2_X1 U514 ( .A1(n533), .A2(n519), .ZN(n462) );
  NOR2_X1 U515 ( .A1(n472), .A2(n462), .ZN(n463) );
  XNOR2_X1 U516 ( .A(n463), .B(KEYINPUT93), .ZN(n464) );
  XNOR2_X1 U517 ( .A(n464), .B(KEYINPUT25), .ZN(n469) );
  XOR2_X1 U518 ( .A(n519), .B(KEYINPUT27), .Z(n473) );
  XOR2_X1 U519 ( .A(KEYINPUT26), .B(KEYINPUT91), .Z(n466) );
  NAND2_X1 U520 ( .A1(n533), .A2(n472), .ZN(n465) );
  XNOR2_X1 U521 ( .A(n466), .B(n465), .ZN(n571) );
  INV_X1 U522 ( .A(n571), .ZN(n548) );
  NAND2_X1 U523 ( .A1(n473), .A2(n548), .ZN(n467) );
  XOR2_X1 U524 ( .A(KEYINPUT92), .B(n467), .Z(n468) );
  NOR2_X1 U525 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U526 ( .A(n470), .B(KEYINPUT94), .ZN(n471) );
  NOR2_X1 U527 ( .A1(n570), .A2(n471), .ZN(n476) );
  XOR2_X1 U528 ( .A(KEYINPUT28), .B(n472), .Z(n531) );
  NAND2_X1 U529 ( .A1(n533), .A2(n531), .ZN(n474) );
  NAND2_X1 U530 ( .A1(n570), .A2(n473), .ZN(n528) );
  NOR2_X1 U531 ( .A1(n474), .A2(n528), .ZN(n475) );
  NOR2_X1 U532 ( .A1(n476), .A2(n475), .ZN(n490) );
  NOR2_X1 U533 ( .A1(n563), .A2(n477), .ZN(n478) );
  XOR2_X1 U534 ( .A(KEYINPUT16), .B(n478), .Z(n479) );
  NOR2_X1 U535 ( .A1(n490), .A2(n479), .ZN(n480) );
  XOR2_X1 U536 ( .A(KEYINPUT95), .B(n480), .Z(n505) );
  NAND2_X1 U537 ( .A1(n493), .A2(n505), .ZN(n488) );
  NOR2_X1 U538 ( .A1(n517), .A2(n488), .ZN(n481) );
  XOR2_X1 U539 ( .A(G1GAT), .B(n481), .Z(n482) );
  XNOR2_X1 U540 ( .A(KEYINPUT34), .B(n482), .ZN(G1324GAT) );
  NOR2_X1 U541 ( .A1(n519), .A2(n488), .ZN(n483) );
  XOR2_X1 U542 ( .A(G8GAT), .B(n483), .Z(G1325GAT) );
  NOR2_X1 U543 ( .A1(n488), .A2(n533), .ZN(n487) );
  XOR2_X1 U544 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n485) );
  XNOR2_X1 U545 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n484) );
  XNOR2_X1 U546 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U547 ( .A(n487), .B(n486), .ZN(G1326GAT) );
  NOR2_X1 U548 ( .A1(n531), .A2(n488), .ZN(n489) );
  XOR2_X1 U549 ( .A(G22GAT), .B(n489), .Z(G1327GAT) );
  NOR2_X1 U550 ( .A1(n585), .A2(n490), .ZN(n491) );
  NAND2_X1 U551 ( .A1(n587), .A2(n491), .ZN(n492) );
  XNOR2_X1 U552 ( .A(KEYINPUT37), .B(n492), .ZN(n516) );
  NAND2_X1 U553 ( .A1(n516), .A2(n493), .ZN(n494) );
  XNOR2_X1 U554 ( .A(KEYINPUT38), .B(n494), .ZN(n502) );
  NOR2_X1 U555 ( .A1(n502), .A2(n517), .ZN(n497) );
  XNOR2_X1 U556 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n495), .B(KEYINPUT98), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n497), .B(n496), .ZN(G1328GAT) );
  NOR2_X1 U559 ( .A1(n519), .A2(n502), .ZN(n498) );
  XOR2_X1 U560 ( .A(G36GAT), .B(n498), .Z(G1329GAT) );
  XNOR2_X1 U561 ( .A(KEYINPUT99), .B(KEYINPUT40), .ZN(n500) );
  NOR2_X1 U562 ( .A1(n533), .A2(n502), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U564 ( .A(G43GAT), .B(n501), .ZN(G1330GAT) );
  NOR2_X1 U565 ( .A1(n502), .A2(n531), .ZN(n503) );
  XOR2_X1 U566 ( .A(G50GAT), .B(n503), .Z(G1331GAT) );
  NAND2_X1 U567 ( .A1(n535), .A2(n550), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n504), .B(KEYINPUT101), .ZN(n515) );
  NAND2_X1 U569 ( .A1(n505), .A2(n515), .ZN(n511) );
  NOR2_X1 U570 ( .A1(n517), .A2(n511), .ZN(n508) );
  XOR2_X1 U571 ( .A(KEYINPUT102), .B(KEYINPUT42), .Z(n506) );
  XNOR2_X1 U572 ( .A(G57GAT), .B(n506), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n508), .B(n507), .ZN(G1332GAT) );
  NOR2_X1 U574 ( .A1(n519), .A2(n511), .ZN(n509) );
  XOR2_X1 U575 ( .A(G64GAT), .B(n509), .Z(G1333GAT) );
  NOR2_X1 U576 ( .A1(n533), .A2(n511), .ZN(n510) );
  XOR2_X1 U577 ( .A(G71GAT), .B(n510), .Z(G1334GAT) );
  NOR2_X1 U578 ( .A1(n531), .A2(n511), .ZN(n513) );
  XNOR2_X1 U579 ( .A(KEYINPUT103), .B(KEYINPUT43), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U581 ( .A(G78GAT), .B(n514), .Z(G1335GAT) );
  NAND2_X1 U582 ( .A1(n516), .A2(n515), .ZN(n525) );
  NOR2_X1 U583 ( .A1(n517), .A2(n525), .ZN(n518) );
  XOR2_X1 U584 ( .A(G85GAT), .B(n518), .Z(G1336GAT) );
  NOR2_X1 U585 ( .A1(n519), .A2(n525), .ZN(n520) );
  XOR2_X1 U586 ( .A(KEYINPUT104), .B(n520), .Z(n521) );
  XNOR2_X1 U587 ( .A(G92GAT), .B(n521), .ZN(G1337GAT) );
  NOR2_X1 U588 ( .A1(n533), .A2(n525), .ZN(n523) );
  XNOR2_X1 U589 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n522) );
  XNOR2_X1 U590 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U591 ( .A(G99GAT), .B(n524), .ZN(G1338GAT) );
  NOR2_X1 U592 ( .A1(n531), .A2(n525), .ZN(n526) );
  XOR2_X1 U593 ( .A(KEYINPUT44), .B(n526), .Z(n527) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n527), .ZN(G1339GAT) );
  NOR2_X1 U595 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U596 ( .A(KEYINPUT109), .B(n530), .Z(n549) );
  NAND2_X1 U597 ( .A1(n549), .A2(n531), .ZN(n532) );
  NOR2_X1 U598 ( .A1(n533), .A2(n532), .ZN(n543) );
  NAND2_X1 U599 ( .A1(n575), .A2(n543), .ZN(n534) );
  XNOR2_X1 U600 ( .A(G113GAT), .B(n534), .ZN(G1340GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT110), .B(KEYINPUT49), .Z(n537) );
  NAND2_X1 U602 ( .A1(n543), .A2(n535), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U604 ( .A(G120GAT), .B(n538), .ZN(G1341GAT) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(KEYINPUT111), .ZN(n542) );
  XOR2_X1 U606 ( .A(KEYINPUT112), .B(KEYINPUT50), .Z(n540) );
  NAND2_X1 U607 ( .A1(n543), .A2(n585), .ZN(n539) );
  XNOR2_X1 U608 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(G1342GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT113), .B(KEYINPUT51), .Z(n545) );
  NAND2_X1 U611 ( .A1(n543), .A2(n563), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(n547) );
  XOR2_X1 U613 ( .A(G134GAT), .B(KEYINPUT114), .Z(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NAND2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n552) );
  NOR2_X1 U616 ( .A1(n550), .A2(n552), .ZN(n551) );
  XOR2_X1 U617 ( .A(G141GAT), .B(n551), .Z(G1344GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT116), .Z(n555) );
  INV_X1 U619 ( .A(n552), .ZN(n562) );
  NAND2_X1 U620 ( .A1(n562), .A2(n553), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U622 ( .A(n556), .B(KEYINPUT52), .Z(n558) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(KEYINPUT115), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1345GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n560) );
  NAND2_X1 U626 ( .A1(n562), .A2(n585), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(G155GAT), .B(n561), .ZN(G1346GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U631 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n566) );
  NAND2_X1 U632 ( .A1(n575), .A2(n567), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(G1348GAT) );
  XOR2_X1 U634 ( .A(G183GAT), .B(KEYINPUT121), .Z(n569) );
  NAND2_X1 U635 ( .A1(n567), .A2(n585), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(G1350GAT) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  AND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U639 ( .A(KEYINPUT123), .B(n574), .Z(n588) );
  NAND2_X1 U640 ( .A1(n588), .A2(n575), .ZN(n579) );
  XOR2_X1 U641 ( .A(KEYINPUT124), .B(KEYINPUT59), .Z(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n582) );
  NAND2_X1 U646 ( .A1(n588), .A2(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n584) );
  XOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT125), .Z(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NAND2_X1 U650 ( .A1(n588), .A2(n585), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U652 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n590) );
  NAND2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

