

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U548 ( .A1(G2104), .A2(n518), .ZN(n866) );
  NOR2_X1 U549 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X2 U550 ( .A1(n524), .A2(n523), .ZN(G160) );
  AND2_X1 U551 ( .A1(n815), .A2(n814), .ZN(n514) );
  INV_X1 U552 ( .A(KEYINPUT27), .ZN(n713) );
  XNOR2_X1 U553 ( .A(n714), .B(n713), .ZN(n716) );
  NOR2_X1 U554 ( .A1(G299), .A2(n725), .ZN(n717) );
  OR2_X1 U555 ( .A1(n724), .A2(n723), .ZN(n728) );
  AND2_X1 U556 ( .A1(n728), .A2(n727), .ZN(n729) );
  NOR2_X1 U557 ( .A1(G1384), .A2(G164), .ZN(n697) );
  NAND2_X1 U558 ( .A1(G160), .A2(G40), .ZN(n698) );
  NAND2_X1 U559 ( .A1(n816), .A2(n514), .ZN(n825) );
  NOR2_X1 U560 ( .A1(G651), .A2(n640), .ZN(n646) );
  NOR2_X1 U561 ( .A1(G651), .A2(G543), .ZN(n654) );
  NAND2_X1 U562 ( .A1(n522), .A2(n521), .ZN(n523) );
  NAND2_X1 U563 ( .A1(n518), .A2(G2104), .ZN(n515) );
  XNOR2_X2 U564 ( .A(n515), .B(KEYINPUT67), .ZN(n872) );
  NAND2_X1 U565 ( .A1(G101), .A2(n872), .ZN(n516) );
  XNOR2_X1 U566 ( .A(n516), .B(KEYINPUT23), .ZN(n524) );
  NOR2_X1 U567 ( .A1(G2105), .A2(G2104), .ZN(n517) );
  XOR2_X2 U568 ( .A(KEYINPUT17), .B(n517), .Z(n870) );
  NAND2_X1 U569 ( .A1(n870), .A2(G137), .ZN(n522) );
  INV_X1 U570 ( .A(G2105), .ZN(n518) );
  NAND2_X1 U571 ( .A1(G125), .A2(n866), .ZN(n520) );
  AND2_X1 U572 ( .A1(G2105), .A2(G2104), .ZN(n867) );
  NAND2_X1 U573 ( .A1(G113), .A2(n867), .ZN(n519) );
  AND2_X1 U574 ( .A1(n520), .A2(n519), .ZN(n521) );
  INV_X1 U575 ( .A(G651), .ZN(n529) );
  NOR2_X1 U576 ( .A1(G543), .A2(n529), .ZN(n525) );
  XOR2_X1 U577 ( .A(KEYINPUT1), .B(n525), .Z(n645) );
  NAND2_X1 U578 ( .A1(G65), .A2(n645), .ZN(n527) );
  XOR2_X1 U579 ( .A(KEYINPUT0), .B(G543), .Z(n640) );
  NAND2_X1 U580 ( .A1(G53), .A2(n646), .ZN(n526) );
  NAND2_X1 U581 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U582 ( .A(KEYINPUT70), .B(n528), .Z(n533) );
  NOR2_X1 U583 ( .A1(n640), .A2(n529), .ZN(n649) );
  NAND2_X1 U584 ( .A1(n649), .A2(G78), .ZN(n531) );
  NAND2_X1 U585 ( .A1(G91), .A2(n654), .ZN(n530) );
  AND2_X1 U586 ( .A1(n531), .A2(n530), .ZN(n532) );
  NAND2_X1 U587 ( .A1(n533), .A2(n532), .ZN(G299) );
  NAND2_X1 U588 ( .A1(n867), .A2(G114), .ZN(n534) );
  XNOR2_X1 U589 ( .A(n534), .B(KEYINPUT88), .ZN(n536) );
  NAND2_X1 U590 ( .A1(G138), .A2(n870), .ZN(n535) );
  NAND2_X1 U591 ( .A1(n536), .A2(n535), .ZN(n540) );
  NAND2_X1 U592 ( .A1(G126), .A2(n866), .ZN(n538) );
  NAND2_X1 U593 ( .A1(G102), .A2(n872), .ZN(n537) );
  NAND2_X1 U594 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U595 ( .A1(n540), .A2(n539), .ZN(G164) );
  NAND2_X1 U596 ( .A1(G77), .A2(n649), .ZN(n542) );
  NAND2_X1 U597 ( .A1(G90), .A2(n654), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U599 ( .A(n543), .B(KEYINPUT9), .ZN(n545) );
  NAND2_X1 U600 ( .A1(G52), .A2(n646), .ZN(n544) );
  NAND2_X1 U601 ( .A1(n545), .A2(n544), .ZN(n548) );
  NAND2_X1 U602 ( .A1(n645), .A2(G64), .ZN(n546) );
  XOR2_X1 U603 ( .A(KEYINPUT68), .B(n546), .Z(n547) );
  NOR2_X1 U604 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U605 ( .A(KEYINPUT69), .B(n549), .Z(G171) );
  INV_X1 U606 ( .A(G171), .ZN(G301) );
  NAND2_X1 U607 ( .A1(G60), .A2(n645), .ZN(n551) );
  NAND2_X1 U608 ( .A1(G85), .A2(n654), .ZN(n550) );
  NAND2_X1 U609 ( .A1(n551), .A2(n550), .ZN(n555) );
  NAND2_X1 U610 ( .A1(G72), .A2(n649), .ZN(n553) );
  NAND2_X1 U611 ( .A1(G47), .A2(n646), .ZN(n552) );
  NAND2_X1 U612 ( .A1(n553), .A2(n552), .ZN(n554) );
  OR2_X1 U613 ( .A1(n555), .A2(n554), .ZN(G290) );
  XOR2_X1 U614 ( .A(G2443), .B(G2446), .Z(n557) );
  XNOR2_X1 U615 ( .A(G2427), .B(G2451), .ZN(n556) );
  XNOR2_X1 U616 ( .A(n557), .B(n556), .ZN(n563) );
  XOR2_X1 U617 ( .A(G2430), .B(G2454), .Z(n559) );
  XNOR2_X1 U618 ( .A(G1348), .B(G1341), .ZN(n558) );
  XNOR2_X1 U619 ( .A(n559), .B(n558), .ZN(n561) );
  XOR2_X1 U620 ( .A(G2435), .B(G2438), .Z(n560) );
  XNOR2_X1 U621 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U622 ( .A(n563), .B(n562), .Z(n564) );
  AND2_X1 U623 ( .A1(G14), .A2(n564), .ZN(G401) );
  AND2_X1 U624 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U625 ( .A(G69), .ZN(G235) );
  INV_X1 U626 ( .A(G132), .ZN(G219) );
  INV_X1 U627 ( .A(G82), .ZN(G220) );
  NAND2_X1 U628 ( .A1(G88), .A2(n654), .ZN(n565) );
  XNOR2_X1 U629 ( .A(n565), .B(KEYINPUT82), .ZN(n567) );
  NAND2_X1 U630 ( .A1(n645), .A2(G62), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n571) );
  NAND2_X1 U632 ( .A1(G75), .A2(n649), .ZN(n569) );
  NAND2_X1 U633 ( .A1(G50), .A2(n646), .ZN(n568) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U635 ( .A1(n571), .A2(n570), .ZN(G166) );
  NAND2_X1 U636 ( .A1(n654), .A2(G89), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n572), .B(KEYINPUT4), .ZN(n574) );
  NAND2_X1 U638 ( .A1(G76), .A2(n649), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(KEYINPUT5), .ZN(n580) );
  NAND2_X1 U641 ( .A1(G63), .A2(n645), .ZN(n577) );
  NAND2_X1 U642 ( .A1(G51), .A2(n646), .ZN(n576) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U644 ( .A(KEYINPUT6), .B(n578), .Z(n579) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U647 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U648 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n583) );
  NAND2_X1 U649 ( .A1(G7), .A2(G661), .ZN(n582) );
  XNOR2_X1 U650 ( .A(n583), .B(n582), .ZN(G223) );
  INV_X1 U651 ( .A(G223), .ZN(n833) );
  AND2_X1 U652 ( .A1(G567), .A2(n833), .ZN(n584) );
  XNOR2_X1 U653 ( .A(n584), .B(KEYINPUT11), .ZN(G234) );
  XOR2_X1 U654 ( .A(KEYINPUT72), .B(KEYINPUT14), .Z(n586) );
  NAND2_X1 U655 ( .A1(G56), .A2(n645), .ZN(n585) );
  XNOR2_X1 U656 ( .A(n586), .B(n585), .ZN(n594) );
  NAND2_X1 U657 ( .A1(n654), .A2(G81), .ZN(n587) );
  XNOR2_X1 U658 ( .A(n587), .B(KEYINPUT12), .ZN(n589) );
  NAND2_X1 U659 ( .A1(G68), .A2(n649), .ZN(n588) );
  NAND2_X1 U660 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U661 ( .A(n590), .B(KEYINPUT13), .ZN(n592) );
  NAND2_X1 U662 ( .A1(G43), .A2(n646), .ZN(n591) );
  NAND2_X1 U663 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U664 ( .A1(n594), .A2(n593), .ZN(n912) );
  INV_X1 U665 ( .A(n912), .ZN(n615) );
  XNOR2_X1 U666 ( .A(G860), .B(KEYINPUT73), .ZN(n611) );
  OR2_X1 U667 ( .A1(n615), .A2(n611), .ZN(G153) );
  NAND2_X1 U668 ( .A1(G301), .A2(G868), .ZN(n595) );
  XNOR2_X1 U669 ( .A(n595), .B(KEYINPUT74), .ZN(n605) );
  INV_X1 U670 ( .A(G868), .ZN(n608) );
  NAND2_X1 U671 ( .A1(n646), .A2(G54), .ZN(n602) );
  NAND2_X1 U672 ( .A1(G79), .A2(n649), .ZN(n597) );
  NAND2_X1 U673 ( .A1(G66), .A2(n645), .ZN(n596) );
  NAND2_X1 U674 ( .A1(n597), .A2(n596), .ZN(n600) );
  NAND2_X1 U675 ( .A1(G92), .A2(n654), .ZN(n598) );
  XNOR2_X1 U676 ( .A(KEYINPUT75), .B(n598), .ZN(n599) );
  NOR2_X1 U677 ( .A1(n600), .A2(n599), .ZN(n601) );
  NAND2_X1 U678 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U679 ( .A(KEYINPUT15), .B(n603), .Z(n923) );
  NAND2_X1 U680 ( .A1(n608), .A2(n923), .ZN(n604) );
  NAND2_X1 U681 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U682 ( .A(KEYINPUT76), .B(n606), .ZN(G284) );
  NOR2_X1 U683 ( .A1(G868), .A2(G299), .ZN(n607) );
  XOR2_X1 U684 ( .A(KEYINPUT77), .B(n607), .Z(n610) );
  NOR2_X1 U685 ( .A1(G286), .A2(n608), .ZN(n609) );
  NOR2_X1 U686 ( .A1(n610), .A2(n609), .ZN(G297) );
  NAND2_X1 U687 ( .A1(n611), .A2(G559), .ZN(n612) );
  INV_X1 U688 ( .A(n923), .ZN(n634) );
  NAND2_X1 U689 ( .A1(n612), .A2(n634), .ZN(n613) );
  XNOR2_X1 U690 ( .A(n613), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U691 ( .A1(n634), .A2(G868), .ZN(n614) );
  NOR2_X1 U692 ( .A1(G559), .A2(n614), .ZN(n617) );
  NOR2_X1 U693 ( .A1(G868), .A2(n615), .ZN(n616) );
  NOR2_X1 U694 ( .A1(n617), .A2(n616), .ZN(G282) );
  NAND2_X1 U695 ( .A1(G111), .A2(n867), .ZN(n619) );
  NAND2_X1 U696 ( .A1(G135), .A2(n870), .ZN(n618) );
  NAND2_X1 U697 ( .A1(n619), .A2(n618), .ZN(n625) );
  NAND2_X1 U698 ( .A1(G99), .A2(n872), .ZN(n620) );
  XNOR2_X1 U699 ( .A(n620), .B(KEYINPUT78), .ZN(n623) );
  NAND2_X1 U700 ( .A1(G123), .A2(n866), .ZN(n621) );
  XNOR2_X1 U701 ( .A(n621), .B(KEYINPUT18), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U703 ( .A1(n625), .A2(n624), .ZN(n965) );
  XNOR2_X1 U704 ( .A(G2096), .B(n965), .ZN(n627) );
  INV_X1 U705 ( .A(G2100), .ZN(n626) );
  NAND2_X1 U706 ( .A1(n627), .A2(n626), .ZN(G156) );
  NAND2_X1 U707 ( .A1(G67), .A2(n645), .ZN(n629) );
  NAND2_X1 U708 ( .A1(G55), .A2(n646), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U710 ( .A1(G80), .A2(n649), .ZN(n631) );
  NAND2_X1 U711 ( .A1(G93), .A2(n654), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U713 ( .A1(n633), .A2(n632), .ZN(n667) );
  NAND2_X1 U714 ( .A1(n634), .A2(G559), .ZN(n664) );
  XOR2_X1 U715 ( .A(n912), .B(n664), .Z(n635) );
  NOR2_X1 U716 ( .A1(G860), .A2(n635), .ZN(n636) );
  XNOR2_X1 U717 ( .A(n667), .B(n636), .ZN(G145) );
  NAND2_X1 U718 ( .A1(G49), .A2(n646), .ZN(n638) );
  NAND2_X1 U719 ( .A1(G74), .A2(G651), .ZN(n637) );
  NAND2_X1 U720 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U721 ( .A1(n645), .A2(n639), .ZN(n643) );
  NAND2_X1 U722 ( .A1(G87), .A2(n640), .ZN(n641) );
  XOR2_X1 U723 ( .A(KEYINPUT79), .B(n641), .Z(n642) );
  NAND2_X1 U724 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U725 ( .A(KEYINPUT80), .B(n644), .ZN(G288) );
  NAND2_X1 U726 ( .A1(G61), .A2(n645), .ZN(n648) );
  NAND2_X1 U727 ( .A1(G48), .A2(n646), .ZN(n647) );
  NAND2_X1 U728 ( .A1(n648), .A2(n647), .ZN(n653) );
  XOR2_X1 U729 ( .A(KEYINPUT2), .B(KEYINPUT81), .Z(n651) );
  NAND2_X1 U730 ( .A1(n649), .A2(G73), .ZN(n650) );
  XOR2_X1 U731 ( .A(n651), .B(n650), .Z(n652) );
  NOR2_X1 U732 ( .A1(n653), .A2(n652), .ZN(n656) );
  NAND2_X1 U733 ( .A1(n654), .A2(G86), .ZN(n655) );
  NAND2_X1 U734 ( .A1(n656), .A2(n655), .ZN(G305) );
  XNOR2_X1 U735 ( .A(G288), .B(G305), .ZN(n657) );
  XNOR2_X1 U736 ( .A(n657), .B(G299), .ZN(n660) );
  XOR2_X1 U737 ( .A(KEYINPUT83), .B(KEYINPUT19), .Z(n658) );
  XNOR2_X1 U738 ( .A(G290), .B(n658), .ZN(n659) );
  XOR2_X1 U739 ( .A(n660), .B(n659), .Z(n662) );
  XNOR2_X1 U740 ( .A(G166), .B(n667), .ZN(n661) );
  XNOR2_X1 U741 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U742 ( .A(n912), .B(n663), .ZN(n881) );
  XOR2_X1 U743 ( .A(n881), .B(n664), .Z(n665) );
  NAND2_X1 U744 ( .A1(G868), .A2(n665), .ZN(n666) );
  XNOR2_X1 U745 ( .A(n666), .B(KEYINPUT84), .ZN(n669) );
  OR2_X1 U746 ( .A1(n667), .A2(G868), .ZN(n668) );
  NAND2_X1 U747 ( .A1(n669), .A2(n668), .ZN(G295) );
  NAND2_X1 U748 ( .A1(G2078), .A2(G2084), .ZN(n670) );
  XOR2_X1 U749 ( .A(KEYINPUT20), .B(n670), .Z(n671) );
  NAND2_X1 U750 ( .A1(G2090), .A2(n671), .ZN(n672) );
  XNOR2_X1 U751 ( .A(KEYINPUT21), .B(n672), .ZN(n673) );
  NAND2_X1 U752 ( .A1(n673), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U753 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U754 ( .A1(G220), .A2(G219), .ZN(n674) );
  XOR2_X1 U755 ( .A(KEYINPUT22), .B(n674), .Z(n675) );
  NOR2_X1 U756 ( .A1(G218), .A2(n675), .ZN(n676) );
  NAND2_X1 U757 ( .A1(G96), .A2(n676), .ZN(n838) );
  NAND2_X1 U758 ( .A1(G2106), .A2(n838), .ZN(n677) );
  XNOR2_X1 U759 ( .A(n677), .B(KEYINPUT85), .ZN(n682) );
  NAND2_X1 U760 ( .A1(G120), .A2(G108), .ZN(n678) );
  NOR2_X1 U761 ( .A1(G235), .A2(n678), .ZN(n679) );
  NAND2_X1 U762 ( .A1(n679), .A2(G57), .ZN(n680) );
  XNOR2_X1 U763 ( .A(KEYINPUT86), .B(n680), .ZN(n837) );
  AND2_X1 U764 ( .A1(n837), .A2(G567), .ZN(n681) );
  NOR2_X1 U765 ( .A1(n682), .A2(n681), .ZN(G319) );
  INV_X1 U766 ( .A(G319), .ZN(n684) );
  NAND2_X1 U767 ( .A1(G661), .A2(G483), .ZN(n683) );
  NOR2_X1 U768 ( .A1(n684), .A2(n683), .ZN(n836) );
  NAND2_X1 U769 ( .A1(n836), .A2(G36), .ZN(n685) );
  XOR2_X1 U770 ( .A(KEYINPUT87), .B(n685), .Z(G176) );
  INV_X1 U771 ( .A(G166), .ZN(G303) );
  NAND2_X1 U772 ( .A1(G140), .A2(n870), .ZN(n687) );
  NAND2_X1 U773 ( .A1(G104), .A2(n872), .ZN(n686) );
  NAND2_X1 U774 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U775 ( .A(KEYINPUT34), .B(n688), .ZN(n694) );
  NAND2_X1 U776 ( .A1(n866), .A2(G128), .ZN(n689) );
  XOR2_X1 U777 ( .A(KEYINPUT89), .B(n689), .Z(n691) );
  NAND2_X1 U778 ( .A1(n867), .A2(G116), .ZN(n690) );
  NAND2_X1 U779 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U780 ( .A(n692), .B(KEYINPUT35), .Z(n693) );
  NOR2_X1 U781 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U782 ( .A(KEYINPUT36), .B(n695), .Z(n696) );
  XNOR2_X1 U783 ( .A(KEYINPUT90), .B(n696), .ZN(n847) );
  XOR2_X1 U784 ( .A(KEYINPUT37), .B(G2067), .Z(n828) );
  AND2_X1 U785 ( .A1(n847), .A2(n828), .ZN(n969) );
  XNOR2_X1 U786 ( .A(n697), .B(KEYINPUT64), .ZN(n700) );
  NOR2_X1 U787 ( .A1(n700), .A2(n698), .ZN(n829) );
  NAND2_X1 U788 ( .A1(n969), .A2(n829), .ZN(n827) );
  INV_X1 U789 ( .A(KEYINPUT94), .ZN(n699) );
  XNOR2_X1 U790 ( .A(n699), .B(n698), .ZN(n701) );
  NAND2_X1 U791 ( .A1(n701), .A2(n700), .ZN(n738) );
  INV_X1 U792 ( .A(n738), .ZN(n712) );
  NAND2_X1 U793 ( .A1(G1996), .A2(n712), .ZN(n703) );
  XOR2_X1 U794 ( .A(KEYINPUT65), .B(KEYINPUT26), .Z(n702) );
  XNOR2_X1 U795 ( .A(n703), .B(n702), .ZN(n704) );
  NAND2_X1 U796 ( .A1(n704), .A2(n912), .ZN(n707) );
  NAND2_X1 U797 ( .A1(G1341), .A2(n738), .ZN(n705) );
  XOR2_X1 U798 ( .A(KEYINPUT100), .B(n705), .Z(n706) );
  XOR2_X1 U799 ( .A(KEYINPUT66), .B(n708), .Z(n722) );
  NOR2_X1 U800 ( .A1(n722), .A2(n923), .ZN(n709) );
  XNOR2_X1 U801 ( .A(n709), .B(KEYINPUT101), .ZN(n720) );
  BUF_X1 U802 ( .A(n738), .Z(n748) );
  NOR2_X1 U803 ( .A1(n712), .A2(G1348), .ZN(n711) );
  NOR2_X1 U804 ( .A1(G2067), .A2(n748), .ZN(n710) );
  NOR2_X1 U805 ( .A1(n711), .A2(n710), .ZN(n718) );
  NAND2_X1 U806 ( .A1(n712), .A2(G2072), .ZN(n714) );
  NAND2_X1 U807 ( .A1(G1956), .A2(n748), .ZN(n715) );
  NAND2_X1 U808 ( .A1(n716), .A2(n715), .ZN(n725) );
  XOR2_X1 U809 ( .A(KEYINPUT102), .B(n717), .Z(n721) );
  AND2_X1 U810 ( .A1(n718), .A2(n721), .ZN(n719) );
  NAND2_X1 U811 ( .A1(n720), .A2(n719), .ZN(n730) );
  INV_X1 U812 ( .A(n721), .ZN(n724) );
  NAND2_X1 U813 ( .A1(n722), .A2(n923), .ZN(n723) );
  NAND2_X1 U814 ( .A1(G299), .A2(n725), .ZN(n726) );
  XNOR2_X1 U815 ( .A(n726), .B(KEYINPUT28), .ZN(n727) );
  NAND2_X1 U816 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U817 ( .A(KEYINPUT29), .B(n731), .Z(n737) );
  XOR2_X1 U818 ( .A(G2078), .B(KEYINPUT98), .Z(n732) );
  XNOR2_X1 U819 ( .A(KEYINPUT25), .B(n732), .ZN(n938) );
  NOR2_X1 U820 ( .A1(n748), .A2(n938), .ZN(n733) );
  XNOR2_X1 U821 ( .A(n733), .B(KEYINPUT99), .ZN(n735) );
  INV_X1 U822 ( .A(G1961), .ZN(n984) );
  NAND2_X1 U823 ( .A1(n984), .A2(n748), .ZN(n734) );
  NAND2_X1 U824 ( .A1(n735), .A2(n734), .ZN(n743) );
  NAND2_X1 U825 ( .A1(n743), .A2(G171), .ZN(n736) );
  NAND2_X1 U826 ( .A1(n737), .A2(n736), .ZN(n764) );
  NAND2_X1 U827 ( .A1(G8), .A2(n748), .ZN(n789) );
  NOR2_X1 U828 ( .A1(G1966), .A2(n789), .ZN(n766) );
  NOR2_X1 U829 ( .A1(G2084), .A2(n738), .ZN(n739) );
  XNOR2_X1 U830 ( .A(KEYINPUT97), .B(n739), .ZN(n761) );
  NAND2_X1 U831 ( .A1(G8), .A2(n761), .ZN(n740) );
  NOR2_X1 U832 ( .A1(n766), .A2(n740), .ZN(n741) );
  XOR2_X1 U833 ( .A(KEYINPUT30), .B(n741), .Z(n742) );
  NOR2_X1 U834 ( .A1(G168), .A2(n742), .ZN(n745) );
  NOR2_X1 U835 ( .A1(G171), .A2(n743), .ZN(n744) );
  NOR2_X1 U836 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U837 ( .A(KEYINPUT31), .B(n746), .Z(n763) );
  INV_X1 U838 ( .A(G8), .ZN(n754) );
  NOR2_X1 U839 ( .A1(G1971), .A2(n789), .ZN(n747) );
  XNOR2_X1 U840 ( .A(KEYINPUT103), .B(n747), .ZN(n751) );
  NOR2_X1 U841 ( .A1(G2090), .A2(n748), .ZN(n749) );
  NOR2_X1 U842 ( .A1(G166), .A2(n749), .ZN(n750) );
  NAND2_X1 U843 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U844 ( .A(n752), .B(KEYINPUT104), .ZN(n753) );
  OR2_X1 U845 ( .A1(n754), .A2(n753), .ZN(n756) );
  AND2_X1 U846 ( .A1(n763), .A2(n756), .ZN(n755) );
  NAND2_X1 U847 ( .A1(n764), .A2(n755), .ZN(n759) );
  INV_X1 U848 ( .A(n756), .ZN(n757) );
  OR2_X1 U849 ( .A1(n757), .A2(G286), .ZN(n758) );
  NAND2_X1 U850 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U851 ( .A(n760), .B(KEYINPUT32), .ZN(n770) );
  INV_X1 U852 ( .A(n761), .ZN(n762) );
  NAND2_X1 U853 ( .A1(G8), .A2(n762), .ZN(n768) );
  AND2_X1 U854 ( .A1(n764), .A2(n763), .ZN(n765) );
  NOR2_X1 U855 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U856 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U857 ( .A1(n770), .A2(n769), .ZN(n788) );
  NOR2_X1 U858 ( .A1(G1976), .A2(G288), .ZN(n776) );
  NOR2_X1 U859 ( .A1(G1971), .A2(G303), .ZN(n771) );
  NOR2_X1 U860 ( .A1(n776), .A2(n771), .ZN(n927) );
  NAND2_X1 U861 ( .A1(n788), .A2(n927), .ZN(n774) );
  INV_X1 U862 ( .A(n789), .ZN(n772) );
  NAND2_X1 U863 ( .A1(G1976), .A2(G288), .ZN(n926) );
  AND2_X1 U864 ( .A1(n772), .A2(n926), .ZN(n773) );
  AND2_X1 U865 ( .A1(n774), .A2(n773), .ZN(n775) );
  NOR2_X1 U866 ( .A1(KEYINPUT33), .A2(n775), .ZN(n779) );
  NAND2_X1 U867 ( .A1(n776), .A2(KEYINPUT33), .ZN(n777) );
  NOR2_X1 U868 ( .A1(n789), .A2(n777), .ZN(n778) );
  NOR2_X1 U869 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U870 ( .A(G1981), .B(G305), .Z(n918) );
  NAND2_X1 U871 ( .A1(n780), .A2(n918), .ZN(n794) );
  NOR2_X1 U872 ( .A1(G1981), .A2(G305), .ZN(n781) );
  XNOR2_X1 U873 ( .A(KEYINPUT24), .B(n781), .ZN(n782) );
  XNOR2_X1 U874 ( .A(KEYINPUT95), .B(n782), .ZN(n783) );
  NOR2_X1 U875 ( .A1(n789), .A2(n783), .ZN(n784) );
  XOR2_X1 U876 ( .A(n784), .B(KEYINPUT96), .Z(n792) );
  NOR2_X1 U877 ( .A1(G2090), .A2(G303), .ZN(n785) );
  XOR2_X1 U878 ( .A(KEYINPUT105), .B(n785), .Z(n786) );
  NAND2_X1 U879 ( .A1(G8), .A2(n786), .ZN(n787) );
  NAND2_X1 U880 ( .A1(n788), .A2(n787), .ZN(n790) );
  NAND2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n791) );
  AND2_X1 U882 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U883 ( .A1(n794), .A2(n793), .ZN(n816) );
  XNOR2_X1 U884 ( .A(G1986), .B(G290), .ZN(n922) );
  NAND2_X1 U885 ( .A1(n922), .A2(n829), .ZN(n815) );
  NAND2_X1 U886 ( .A1(G119), .A2(n866), .ZN(n796) );
  NAND2_X1 U887 ( .A1(G107), .A2(n867), .ZN(n795) );
  NAND2_X1 U888 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U889 ( .A(KEYINPUT91), .B(n797), .ZN(n802) );
  NAND2_X1 U890 ( .A1(G131), .A2(n870), .ZN(n799) );
  NAND2_X1 U891 ( .A1(G95), .A2(n872), .ZN(n798) );
  NAND2_X1 U892 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U893 ( .A(KEYINPUT92), .B(n800), .Z(n801) );
  NAND2_X1 U894 ( .A1(n802), .A2(n801), .ZN(n859) );
  NAND2_X1 U895 ( .A1(G1991), .A2(n859), .ZN(n803) );
  XNOR2_X1 U896 ( .A(n803), .B(KEYINPUT93), .ZN(n812) );
  NAND2_X1 U897 ( .A1(G129), .A2(n866), .ZN(n805) );
  NAND2_X1 U898 ( .A1(G117), .A2(n867), .ZN(n804) );
  NAND2_X1 U899 ( .A1(n805), .A2(n804), .ZN(n808) );
  NAND2_X1 U900 ( .A1(n872), .A2(G105), .ZN(n806) );
  XOR2_X1 U901 ( .A(KEYINPUT38), .B(n806), .Z(n807) );
  NOR2_X1 U902 ( .A1(n808), .A2(n807), .ZN(n810) );
  NAND2_X1 U903 ( .A1(n870), .A2(G141), .ZN(n809) );
  NAND2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n863) );
  AND2_X1 U905 ( .A1(G1996), .A2(n863), .ZN(n811) );
  NOR2_X1 U906 ( .A1(n812), .A2(n811), .ZN(n970) );
  INV_X1 U907 ( .A(n829), .ZN(n813) );
  NOR2_X1 U908 ( .A1(n970), .A2(n813), .ZN(n819) );
  INV_X1 U909 ( .A(n819), .ZN(n814) );
  NOR2_X1 U910 ( .A1(G1996), .A2(n863), .ZN(n958) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n817) );
  NOR2_X1 U912 ( .A1(G1991), .A2(n859), .ZN(n966) );
  NOR2_X1 U913 ( .A1(n817), .A2(n966), .ZN(n818) );
  NOR2_X1 U914 ( .A1(n819), .A2(n818), .ZN(n820) );
  NOR2_X1 U915 ( .A1(n958), .A2(n820), .ZN(n821) );
  XNOR2_X1 U916 ( .A(n821), .B(KEYINPUT106), .ZN(n822) );
  XNOR2_X1 U917 ( .A(n822), .B(KEYINPUT39), .ZN(n823) );
  NAND2_X1 U918 ( .A1(n823), .A2(n829), .ZN(n824) );
  NAND2_X1 U919 ( .A1(n825), .A2(n824), .ZN(n826) );
  NAND2_X1 U920 ( .A1(n827), .A2(n826), .ZN(n831) );
  NOR2_X1 U921 ( .A1(n828), .A2(n847), .ZN(n973) );
  NAND2_X1 U922 ( .A1(n973), .A2(n829), .ZN(n830) );
  NAND2_X1 U923 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U924 ( .A(n832), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n833), .ZN(G217) );
  AND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U927 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U929 ( .A1(n836), .A2(n835), .ZN(G188) );
  XNOR2_X1 U930 ( .A(G120), .B(KEYINPUT107), .ZN(G236) );
  XOR2_X1 U931 ( .A(G108), .B(KEYINPUT116), .Z(G238) );
  INV_X1 U933 ( .A(G96), .ZN(G221) );
  NOR2_X1 U934 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U935 ( .A(G325), .ZN(G261) );
  NAND2_X1 U936 ( .A1(G112), .A2(n867), .ZN(n840) );
  NAND2_X1 U937 ( .A1(G100), .A2(n872), .ZN(n839) );
  NAND2_X1 U938 ( .A1(n840), .A2(n839), .ZN(n846) );
  NAND2_X1 U939 ( .A1(n866), .A2(G124), .ZN(n841) );
  XNOR2_X1 U940 ( .A(n841), .B(KEYINPUT44), .ZN(n843) );
  NAND2_X1 U941 ( .A1(G136), .A2(n870), .ZN(n842) );
  NAND2_X1 U942 ( .A1(n843), .A2(n842), .ZN(n844) );
  XOR2_X1 U943 ( .A(KEYINPUT111), .B(n844), .Z(n845) );
  NOR2_X1 U944 ( .A1(n846), .A2(n845), .ZN(G162) );
  XOR2_X1 U945 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n849) );
  XOR2_X1 U946 ( .A(n847), .B(G164), .Z(n848) );
  XNOR2_X1 U947 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n965), .B(n850), .ZN(n861) );
  NAND2_X1 U949 ( .A1(G139), .A2(n870), .ZN(n852) );
  NAND2_X1 U950 ( .A1(G103), .A2(n872), .ZN(n851) );
  NAND2_X1 U951 ( .A1(n852), .A2(n851), .ZN(n858) );
  NAND2_X1 U952 ( .A1(n867), .A2(G115), .ZN(n853) );
  XOR2_X1 U953 ( .A(KEYINPUT113), .B(n853), .Z(n855) );
  NAND2_X1 U954 ( .A1(n866), .A2(G127), .ZN(n854) );
  NAND2_X1 U955 ( .A1(n855), .A2(n854), .ZN(n856) );
  XOR2_X1 U956 ( .A(KEYINPUT47), .B(n856), .Z(n857) );
  NOR2_X1 U957 ( .A1(n858), .A2(n857), .ZN(n960) );
  XNOR2_X1 U958 ( .A(n859), .B(n960), .ZN(n860) );
  XNOR2_X1 U959 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U960 ( .A(n862), .B(G162), .Z(n865) );
  XOR2_X1 U961 ( .A(G160), .B(n863), .Z(n864) );
  XNOR2_X1 U962 ( .A(n865), .B(n864), .ZN(n879) );
  NAND2_X1 U963 ( .A1(G130), .A2(n866), .ZN(n869) );
  NAND2_X1 U964 ( .A1(G118), .A2(n867), .ZN(n868) );
  NAND2_X1 U965 ( .A1(n869), .A2(n868), .ZN(n877) );
  NAND2_X1 U966 ( .A1(n870), .A2(G142), .ZN(n871) );
  XNOR2_X1 U967 ( .A(n871), .B(KEYINPUT112), .ZN(n874) );
  NAND2_X1 U968 ( .A1(G106), .A2(n872), .ZN(n873) );
  NAND2_X1 U969 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U970 ( .A(n875), .B(KEYINPUT45), .Z(n876) );
  NOR2_X1 U971 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U972 ( .A(n879), .B(n878), .Z(n880) );
  NOR2_X1 U973 ( .A1(G37), .A2(n880), .ZN(G395) );
  XNOR2_X1 U974 ( .A(G286), .B(n923), .ZN(n882) );
  XNOR2_X1 U975 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U976 ( .A(n883), .B(G301), .ZN(n884) );
  NOR2_X1 U977 ( .A1(G37), .A2(n884), .ZN(G397) );
  XOR2_X1 U978 ( .A(KEYINPUT109), .B(G1986), .Z(n886) );
  XNOR2_X1 U979 ( .A(G1961), .B(G1956), .ZN(n885) );
  XNOR2_X1 U980 ( .A(n886), .B(n885), .ZN(n887) );
  XOR2_X1 U981 ( .A(n887), .B(KEYINPUT41), .Z(n889) );
  XNOR2_X1 U982 ( .A(G1996), .B(G1991), .ZN(n888) );
  XNOR2_X1 U983 ( .A(n889), .B(n888), .ZN(n893) );
  XOR2_X1 U984 ( .A(G1966), .B(G1971), .Z(n891) );
  XNOR2_X1 U985 ( .A(G1981), .B(G1976), .ZN(n890) );
  XNOR2_X1 U986 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U987 ( .A(n893), .B(n892), .Z(n895) );
  XNOR2_X1 U988 ( .A(G2474), .B(KEYINPUT110), .ZN(n894) );
  XNOR2_X1 U989 ( .A(n895), .B(n894), .ZN(G229) );
  XOR2_X1 U990 ( .A(G2096), .B(KEYINPUT108), .Z(n897) );
  XNOR2_X1 U991 ( .A(G2090), .B(KEYINPUT43), .ZN(n896) );
  XNOR2_X1 U992 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U993 ( .A(n898), .B(KEYINPUT42), .Z(n900) );
  XNOR2_X1 U994 ( .A(G2067), .B(G2072), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n900), .B(n899), .ZN(n904) );
  XOR2_X1 U996 ( .A(G2678), .B(G2100), .Z(n902) );
  XNOR2_X1 U997 ( .A(G2078), .B(G2084), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n904), .B(n903), .ZN(G227) );
  NOR2_X1 U1000 ( .A1(G395), .A2(G397), .ZN(n905) );
  XOR2_X1 U1001 ( .A(KEYINPUT115), .B(n905), .Z(n911) );
  NOR2_X1 U1002 ( .A1(G229), .A2(G227), .ZN(n906) );
  XOR2_X1 U1003 ( .A(KEYINPUT49), .B(n906), .Z(n907) );
  NAND2_X1 U1004 ( .A1(G319), .A2(n907), .ZN(n908) );
  NOR2_X1 U1005 ( .A1(G401), .A2(n908), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(KEYINPUT114), .B(n909), .ZN(n910) );
  NAND2_X1 U1007 ( .A1(n911), .A2(n910), .ZN(G225) );
  INV_X1 U1008 ( .A(G225), .ZN(G308) );
  INV_X1 U1009 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1010 ( .A(KEYINPUT125), .B(KEYINPUT126), .ZN(n1016) );
  XNOR2_X1 U1011 ( .A(G171), .B(G1961), .ZN(n916) );
  XOR2_X1 U1012 ( .A(n912), .B(G1341), .Z(n914) );
  XNOR2_X1 U1013 ( .A(G299), .B(G1956), .ZN(n913) );
  NOR2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(n933) );
  XOR2_X1 U1016 ( .A(G1966), .B(G168), .Z(n917) );
  XNOR2_X1 U1017 ( .A(KEYINPUT123), .B(n917), .ZN(n919) );
  NAND2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1019 ( .A(n920), .B(KEYINPUT57), .ZN(n931) );
  AND2_X1 U1020 ( .A1(G303), .A2(G1971), .ZN(n921) );
  NOR2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n925) );
  XOR2_X1 U1022 ( .A(G1348), .B(n923), .Z(n924) );
  NAND2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n929) );
  NAND2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n928) );
  NOR2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1027 ( .A1(n933), .A2(n932), .ZN(n1006) );
  NAND2_X1 U1028 ( .A1(G16), .A2(KEYINPUT56), .ZN(n934) );
  NOR2_X1 U1029 ( .A1(n1006), .A2(n934), .ZN(n1014) );
  XNOR2_X1 U1030 ( .A(G2084), .B(G34), .ZN(n935) );
  XNOR2_X1 U1031 ( .A(n935), .B(KEYINPUT54), .ZN(n953) );
  XNOR2_X1 U1032 ( .A(G2090), .B(G35), .ZN(n950) );
  XNOR2_X1 U1033 ( .A(G2067), .B(G26), .ZN(n937) );
  XNOR2_X1 U1034 ( .A(G33), .B(G2072), .ZN(n936) );
  NOR2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(n942) );
  XNOR2_X1 U1036 ( .A(n938), .B(G27), .ZN(n940) );
  XNOR2_X1 U1037 ( .A(G32), .B(G1996), .ZN(n939) );
  NOR2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(G1991), .B(KEYINPUT119), .ZN(n943) );
  XNOR2_X1 U1041 ( .A(n943), .B(G25), .ZN(n944) );
  NAND2_X1 U1042 ( .A1(G28), .A2(n944), .ZN(n945) );
  XNOR2_X1 U1043 ( .A(KEYINPUT120), .B(n945), .ZN(n946) );
  NOR2_X1 U1044 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1045 ( .A(KEYINPUT53), .B(n948), .ZN(n949) );
  NOR2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1047 ( .A(n951), .B(KEYINPUT121), .ZN(n952) );
  NOR2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(KEYINPUT122), .B(n954), .ZN(n955) );
  NOR2_X1 U1050 ( .A1(G29), .A2(n955), .ZN(n956) );
  XNOR2_X1 U1051 ( .A(n956), .B(KEYINPUT55), .ZN(n983) );
  XOR2_X1 U1052 ( .A(G2090), .B(G162), .Z(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1054 ( .A(KEYINPUT51), .B(n959), .Z(n979) );
  XNOR2_X1 U1055 ( .A(G2072), .B(n960), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(G164), .B(G2078), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(n961), .B(KEYINPUT118), .ZN(n962) );
  NAND2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(n964), .B(KEYINPUT50), .ZN(n977) );
  NOR2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1061 ( .A(KEYINPUT117), .B(n967), .ZN(n968) );
  NOR2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n975) );
  XNOR2_X1 U1063 ( .A(G160), .B(G2084), .ZN(n971) );
  NAND2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1068 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(KEYINPUT52), .B(n980), .ZN(n981) );
  NAND2_X1 U1070 ( .A1(G29), .A2(n981), .ZN(n982) );
  NAND2_X1 U1071 ( .A1(n983), .A2(n982), .ZN(n1011) );
  XNOR2_X1 U1072 ( .A(G5), .B(n984), .ZN(n997) );
  XNOR2_X1 U1073 ( .A(G1348), .B(KEYINPUT59), .ZN(n985) );
  XNOR2_X1 U1074 ( .A(n985), .B(G4), .ZN(n989) );
  XNOR2_X1 U1075 ( .A(G1341), .B(G19), .ZN(n987) );
  XNOR2_X1 U1076 ( .A(G1956), .B(G20), .ZN(n986) );
  NOR2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n992) );
  XNOR2_X1 U1079 ( .A(KEYINPUT124), .B(G1981), .ZN(n990) );
  XNOR2_X1 U1080 ( .A(G6), .B(n990), .ZN(n991) );
  NOR2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1082 ( .A(KEYINPUT60), .B(n993), .Z(n995) );
  XNOR2_X1 U1083 ( .A(G1966), .B(G21), .ZN(n994) );
  NOR2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n1004) );
  XNOR2_X1 U1086 ( .A(G1976), .B(G23), .ZN(n999) );
  XNOR2_X1 U1087 ( .A(G1971), .B(G22), .ZN(n998) );
  NOR2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1001) );
  XOR2_X1 U1089 ( .A(G1986), .B(G24), .Z(n1000) );
  NAND2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1091 ( .A(KEYINPUT58), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(n1005), .B(KEYINPUT61), .ZN(n1008) );
  NOR2_X1 U1094 ( .A1(KEYINPUT56), .A2(n1006), .ZN(n1007) );
  NOR2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1096 ( .A1(G16), .A2(n1009), .ZN(n1010) );
  NOR2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1098 ( .A1(n1012), .A2(G11), .ZN(n1013) );
  NOR2_X1 U1099 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1100 ( .A(n1016), .B(n1015), .ZN(n1017) );
  XNOR2_X1 U1101 ( .A(KEYINPUT62), .B(n1017), .ZN(G150) );
  INV_X1 U1102 ( .A(G150), .ZN(G311) );
endmodule

