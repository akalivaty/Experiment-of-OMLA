//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 0 1 0 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 0 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n556, new_n558, new_n559,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n587, new_n588, new_n589,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n622, new_n624, new_n625, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1210, new_n1211, new_n1212;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT66), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  OR4_X1    g028(.A1(G237), .A2(G236), .A3(G235), .A4(G238), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n454), .A2(G567), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n457), .A2(KEYINPUT68), .ZN(new_n458));
  AOI21_X1  g033(.A(new_n458), .B1(new_n453), .B2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(KEYINPUT68), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT69), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n463), .B(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  AND3_X1   g044(.A1(new_n467), .A2(new_n469), .A3(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(G2105), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n467), .A2(new_n469), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G137), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(G101), .A3(G2104), .ZN(new_n476));
  XOR2_X1   g051(.A(new_n476), .B(KEYINPUT70), .Z(new_n477));
  AND3_X1   g052(.A1(new_n471), .A2(new_n474), .A3(new_n477), .ZN(G160));
  AND3_X1   g053(.A1(new_n467), .A2(new_n469), .A3(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(KEYINPUT71), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT71), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n481), .B1(new_n472), .B2(new_n475), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  AOI22_X1  g058(.A1(new_n483), .A2(G124), .B1(G136), .B2(new_n473), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G112), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n484), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  NAND4_X1  g065(.A1(new_n467), .A2(new_n469), .A3(G138), .A4(new_n475), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  XNOR2_X1  g067(.A(KEYINPUT3), .B(G2104), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n493), .A2(new_n494), .A3(G138), .A4(new_n475), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n479), .A2(G126), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n475), .A2(G114), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT72), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OR2_X1    g075(.A1(G102), .A2(G2105), .ZN(new_n501));
  INV_X1    g076(.A(G114), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G2105), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n501), .A2(new_n503), .A3(new_n504), .A4(G2104), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n497), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n496), .A2(new_n507), .ZN(G164));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n515), .A2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND3_X1  g095(.A1(new_n510), .A2(G51), .A3(G543), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n509), .A2(new_n510), .A3(G89), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n521), .A2(new_n522), .A3(new_n524), .A4(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(G168));
  NAND3_X1  g102(.A1(new_n509), .A2(new_n510), .A3(G90), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n510), .A2(G52), .A3(G543), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT74), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT74), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n528), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(G543), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(KEYINPUT5), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT5), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G543), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G64), .ZN(new_n540));
  INV_X1    g115(.A(G77), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n539), .A2(new_n540), .B1(new_n541), .B2(new_n535), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT73), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI221_X1 g119(.A(KEYINPUT73), .B1(new_n541), .B2(new_n535), .C1(new_n539), .C2(new_n540), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n544), .A2(G651), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n534), .A2(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  INV_X1    g124(.A(G43), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n511), .A2(new_n549), .B1(new_n513), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(new_n517), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(G188));
  NAND3_X1  g135(.A1(new_n536), .A2(new_n538), .A3(G65), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  AND3_X1   g137(.A1(new_n561), .A2(KEYINPUT76), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g138(.A(KEYINPUT76), .B1(new_n561), .B2(new_n562), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT77), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n565), .A2(new_n566), .A3(G651), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n561), .A2(new_n562), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT76), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n561), .A2(KEYINPUT76), .A3(new_n562), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n570), .A2(G651), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(KEYINPUT77), .ZN(new_n573));
  INV_X1    g148(.A(new_n511), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n567), .A2(new_n573), .B1(G91), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT78), .ZN(new_n576));
  AND3_X1   g151(.A1(new_n510), .A2(G53), .A3(G543), .ZN(new_n577));
  NAND2_X1  g152(.A1(KEYINPUT75), .A2(KEYINPUT9), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n577), .B(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n575), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n574), .A2(G91), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n566), .B1(new_n565), .B2(G651), .ZN(new_n582));
  NOR4_X1   g157(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT77), .A4(new_n517), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n581), .B(new_n579), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(KEYINPUT78), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n580), .A2(new_n585), .ZN(G299));
  INV_X1    g161(.A(KEYINPUT79), .ZN(new_n587));
  AND2_X1   g162(.A1(new_n526), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n526), .A2(new_n587), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n588), .A2(new_n589), .ZN(G286));
  NAND2_X1  g165(.A1(new_n574), .A2(G87), .ZN(new_n591));
  INV_X1    g166(.A(new_n513), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G49), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(G288));
  INV_X1    g170(.A(G86), .ZN(new_n596));
  OR3_X1    g171(.A1(new_n511), .A2(KEYINPUT80), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(KEYINPUT80), .B1(new_n511), .B2(new_n596), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(G73), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G61), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n539), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(G48), .A2(new_n592), .B1(new_n602), .B2(G651), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n599), .A2(new_n603), .ZN(G305));
  INV_X1    g179(.A(G85), .ZN(new_n605));
  INV_X1    g180(.A(G47), .ZN(new_n606));
  OAI22_X1  g181(.A1(new_n511), .A2(new_n605), .B1(new_n513), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(new_n517), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n607), .A2(new_n609), .ZN(G290));
  NAND2_X1  g185(.A1(G301), .A2(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n574), .A2(G92), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT10), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n509), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n614));
  INV_X1    g189(.A(G54), .ZN(new_n615));
  OAI22_X1  g190(.A1(new_n614), .A2(new_n517), .B1(new_n615), .B2(new_n513), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n611), .B1(new_n617), .B2(G868), .ZN(G321));
  XNOR2_X1  g193(.A(G321), .B(KEYINPUT81), .ZN(G284));
  MUX2_X1   g194(.A(G299), .B(G286), .S(G868), .Z(G280));
  XOR2_X1   g195(.A(G280), .B(KEYINPUT82), .Z(G297));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n617), .B1(new_n622), .B2(G860), .ZN(G148));
  NAND2_X1  g198(.A1(new_n617), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G868), .B2(new_n554), .ZN(G323));
  XOR2_X1   g201(.A(KEYINPUT83), .B(KEYINPUT11), .Z(new_n627));
  XNOR2_X1  g202(.A(G323), .B(new_n627), .ZN(G282));
  NAND2_X1  g203(.A1(new_n473), .A2(G135), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n475), .A2(G111), .ZN(new_n631));
  NOR3_X1   g206(.A1(new_n472), .A2(new_n481), .A3(new_n475), .ZN(new_n632));
  AOI21_X1  g207(.A(KEYINPUT71), .B1(new_n493), .B2(G2105), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(G123), .ZN(new_n635));
  OAI221_X1 g210(.A(new_n629), .B1(new_n630), .B2(new_n631), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT84), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT85), .B(G2096), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n466), .A2(G2105), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n493), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT13), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2100), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n639), .A2(new_n644), .ZN(G156));
  XNOR2_X1  g220(.A(G2427), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2430), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT15), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n648), .A2(G2435), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(G2435), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(KEYINPUT14), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2443), .B(G2446), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2451), .B(G2454), .Z(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n653), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n659), .A2(G14), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT87), .Z(G401));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  XOR2_X1   g238(.A(G2067), .B(G2678), .Z(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n663), .B1(new_n667), .B2(KEYINPUT18), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2096), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G2100), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n667), .A2(KEYINPUT17), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n665), .A2(new_n666), .ZN(new_n672));
  AOI21_X1  g247(.A(KEYINPUT18), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n670), .B(new_n673), .Z(G227));
  XOR2_X1   g249(.A(G1956), .B(G2474), .Z(new_n675));
  XOR2_X1   g250(.A(G1961), .B(G1966), .Z(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n675), .A2(new_n676), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT20), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n681), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n678), .A2(new_n680), .A3(new_n682), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n685), .B(new_n686), .C1(new_n684), .C2(new_n683), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  INV_X1    g265(.A(G1981), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n689), .B(new_n693), .ZN(G229));
  MUX2_X1   g269(.A(G24), .B(G290), .S(G16), .Z(new_n695));
  XOR2_X1   g270(.A(KEYINPUT88), .B(G1986), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G25), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n473), .A2(G131), .ZN(new_n700));
  OR2_X1    g275(.A1(G95), .A2(G2105), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n701), .B(G2104), .C1(G107), .C2(new_n475), .ZN(new_n702));
  INV_X1    g277(.A(G119), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n700), .B(new_n702), .C1(new_n634), .C2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n699), .B1(new_n705), .B2(new_n698), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT35), .B(G1991), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n706), .B(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n697), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G23), .ZN(new_n713));
  INV_X1    g288(.A(G288), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(new_n712), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT33), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(G1976), .ZN(new_n717));
  NOR2_X1   g292(.A1(G16), .A2(G22), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G166), .B2(G16), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT91), .B(G1971), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT34), .ZN(new_n723));
  MUX2_X1   g298(.A(G6), .B(G305), .S(G16), .Z(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT32), .B(G1981), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT89), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT90), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n724), .B(new_n727), .ZN(new_n728));
  OR3_X1    g303(.A1(new_n722), .A2(new_n723), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n723), .B1(new_n722), .B2(new_n728), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n711), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n732), .ZN(new_n734));
  AOI211_X1 g309(.A(new_n734), .B(new_n711), .C1(new_n729), .C2(new_n730), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(KEYINPUT23), .B1(new_n712), .B2(G20), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G299), .B2(G16), .ZN(new_n738));
  AND3_X1   g313(.A1(new_n712), .A2(KEYINPUT23), .A3(G20), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G1956), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n698), .A2(G35), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G162), .B2(new_n698), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT29), .B(G2090), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n698), .A2(G26), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT28), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n473), .A2(G140), .ZN(new_n751));
  OR2_X1    g326(.A1(G104), .A2(G2105), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n752), .B(G2104), .C1(G116), .C2(new_n475), .ZN(new_n753));
  INV_X1    g328(.A(G128), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n751), .B(new_n753), .C1(new_n634), .C2(new_n754), .ZN(new_n755));
  AND3_X1   g330(.A1(new_n755), .A2(KEYINPUT95), .A3(G29), .ZN(new_n756));
  AOI21_X1  g331(.A(KEYINPUT95), .B1(new_n755), .B2(G29), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n750), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G2067), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n712), .A2(G5), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G171), .B2(new_n712), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(G1961), .Z(new_n763));
  NAND2_X1  g338(.A1(new_n483), .A2(G129), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n473), .A2(G141), .ZN(new_n765));
  NAND3_X1  g340(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT26), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n640), .A2(G105), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT97), .Z(new_n769));
  NAND4_X1  g344(.A1(new_n764), .A2(new_n765), .A3(new_n767), .A4(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n771), .A2(G29), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G29), .B2(G32), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT27), .B(G1996), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT31), .B(G11), .Z(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n773), .B2(new_n774), .ZN(new_n777));
  AND3_X1   g352(.A1(new_n763), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n743), .A2(new_n748), .A3(new_n760), .A4(new_n778), .ZN(new_n779));
  OR2_X1    g354(.A1(G29), .A2(G33), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n640), .A2(G103), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT96), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(KEYINPUT25), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n781), .B(KEYINPUT96), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT25), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(G115), .A2(G2104), .ZN(new_n788));
  INV_X1    g363(.A(G127), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n472), .B2(new_n789), .ZN(new_n790));
  AOI22_X1  g365(.A1(new_n790), .A2(G2105), .B1(new_n473), .B2(G139), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n784), .A2(new_n787), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n780), .B1(new_n792), .B2(new_n698), .ZN(new_n793));
  INV_X1    g368(.A(G2072), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n617), .A2(G16), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G4), .B2(G16), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT93), .B(G1348), .Z(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  OAI221_X1 g374(.A(new_n795), .B1(new_n637), .B2(new_n698), .C1(new_n797), .C2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n698), .A2(G27), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G164), .B2(new_n698), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G2078), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT30), .B(G28), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n803), .B1(new_n698), .B2(new_n804), .ZN(new_n805));
  OR2_X1    g380(.A1(KEYINPUT24), .A2(G34), .ZN(new_n806));
  NAND2_X1  g381(.A1(KEYINPUT24), .A2(G34), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n806), .A2(new_n698), .A3(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G160), .B2(new_n698), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(G2084), .Z(new_n810));
  NOR2_X1   g385(.A1(G16), .A2(G19), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(new_n554), .B2(G16), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT94), .B(G1341), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n805), .A2(new_n810), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(KEYINPUT98), .B1(G16), .B2(G21), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n526), .A2(new_n712), .ZN(new_n817));
  MUX2_X1   g392(.A(new_n816), .B(KEYINPUT98), .S(new_n817), .Z(new_n818));
  INV_X1    g393(.A(G1966), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NOR4_X1   g395(.A1(new_n779), .A2(new_n800), .A3(new_n815), .A4(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n793), .A2(new_n794), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n797), .A2(new_n799), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n821), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n736), .A2(new_n825), .ZN(G311));
  OR2_X1    g401(.A1(new_n736), .A2(new_n825), .ZN(G150));
  INV_X1    g402(.A(G93), .ZN(new_n828));
  INV_X1    g403(.A(G55), .ZN(new_n829));
  OAI22_X1  g404(.A1(new_n511), .A2(new_n828), .B1(new_n513), .B2(new_n829), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n831), .A2(new_n517), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(G860), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT37), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n833), .A2(KEYINPUT99), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT99), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(new_n830), .B2(new_n832), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n837), .A2(new_n554), .A3(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n554), .ZN(new_n841));
  INV_X1    g416(.A(new_n833), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n841), .A2(new_n842), .A3(new_n838), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT38), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n617), .A2(G559), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT39), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT100), .Z(new_n850));
  OAI21_X1  g425(.A(new_n834), .B1(new_n847), .B2(new_n848), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n836), .B1(new_n850), .B2(new_n851), .ZN(G145));
  INV_X1    g427(.A(KEYINPUT103), .ZN(new_n853));
  INV_X1    g428(.A(G130), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n853), .B1(new_n634), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n483), .A2(KEYINPUT103), .A3(G130), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n858));
  INV_X1    g433(.A(G118), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n858), .B1(new_n859), .B2(G2105), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n473), .A2(G142), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT102), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n857), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n642), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n704), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n483), .A2(G119), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n867), .A2(new_n642), .A3(new_n700), .A4(new_n702), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n864), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n860), .B1(new_n855), .B2(new_n856), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n871), .A2(new_n866), .A3(new_n863), .A4(new_n868), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  AOI22_X1  g448(.A1(new_n483), .A2(G128), .B1(G140), .B2(new_n473), .ZN(new_n874));
  AOI22_X1  g449(.A1(G126), .A2(new_n479), .B1(new_n500), .B2(new_n505), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n492), .A2(new_n495), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n874), .A2(new_n877), .A3(new_n753), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n755), .A2(G164), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n878), .A2(new_n879), .A3(new_n770), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n770), .B1(new_n878), .B2(new_n879), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT101), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n792), .A2(new_n882), .ZN(new_n883));
  NOR3_X1   g458(.A1(new_n880), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n784), .A2(new_n787), .A3(KEYINPUT101), .A4(new_n791), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n877), .B1(new_n874), .B2(new_n753), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n755), .A2(G164), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n771), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n878), .A2(new_n879), .A3(new_n770), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n886), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n873), .B1(new_n884), .B2(new_n891), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n870), .A2(new_n872), .ZN(new_n893));
  INV_X1    g468(.A(new_n886), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(new_n880), .B2(new_n881), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n889), .A2(new_n882), .A3(new_n792), .A4(new_n890), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n893), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n892), .A2(KEYINPUT104), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n637), .A2(G162), .ZN(new_n899));
  OR2_X1    g474(.A1(new_n636), .A2(KEYINPUT84), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n636), .A2(KEYINPUT84), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n900), .A2(new_n489), .A3(new_n901), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n899), .A2(new_n902), .A3(G160), .ZN(new_n903));
  AOI21_X1  g478(.A(G160), .B1(new_n899), .B2(new_n902), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT104), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n893), .A2(new_n895), .A3(new_n896), .A4(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n898), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT105), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT105), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n898), .A2(new_n905), .A3(new_n910), .A4(new_n907), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(G37), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n892), .B(new_n897), .C1(new_n903), .C2(new_n904), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT106), .ZN(new_n916));
  AOI21_X1  g491(.A(G37), .B1(new_n909), .B2(new_n911), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(new_n918), .A3(new_n914), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n916), .A2(KEYINPUT40), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT40), .B1(new_n916), .B2(new_n919), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(G395));
  NOR2_X1   g497(.A1(new_n842), .A2(G868), .ZN(new_n923));
  XOR2_X1   g498(.A(G303), .B(G290), .Z(new_n924));
  XNOR2_X1  g499(.A(G305), .B(new_n714), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n924), .B(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(KEYINPUT42), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n580), .A2(new_n585), .A3(new_n617), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n617), .B1(new_n580), .B2(new_n585), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  XOR2_X1   g508(.A(new_n624), .B(new_n844), .Z(new_n934));
  OAI21_X1  g509(.A(KEYINPUT107), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT41), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n930), .B2(new_n931), .ZN(new_n937));
  INV_X1    g512(.A(new_n617), .ZN(new_n938));
  NAND2_X1  g513(.A1(G299), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n580), .A2(new_n585), .A3(new_n617), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n939), .A2(KEYINPUT41), .A3(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n937), .A2(new_n941), .A3(new_n934), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n935), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n937), .A2(new_n941), .A3(new_n934), .A4(KEYINPUT107), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n929), .B1(new_n945), .B2(KEYINPUT108), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n927), .A2(KEYINPUT42), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n946), .B(new_n948), .C1(KEYINPUT108), .C2(new_n945), .ZN(new_n949));
  INV_X1    g524(.A(new_n945), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n950), .B(new_n951), .C1(new_n947), .C2(new_n929), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n923), .B1(new_n953), .B2(G868), .ZN(G295));
  AOI21_X1  g529(.A(new_n923), .B1(new_n953), .B2(G868), .ZN(G331));
  INV_X1    g530(.A(new_n844), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n534), .B(new_n546), .C1(new_n588), .C2(new_n589), .ZN(new_n957));
  NAND2_X1  g532(.A1(G301), .A2(G168), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n959), .B1(new_n957), .B2(new_n958), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n956), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n957), .A2(new_n958), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT110), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n965), .A2(new_n844), .A3(new_n960), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n937), .A2(new_n967), .A3(new_n941), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT112), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n963), .A2(new_n966), .A3(new_n971), .ZN(new_n972));
  OAI211_X1 g547(.A(KEYINPUT111), .B(new_n956), .C1(new_n961), .C2(new_n962), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n932), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n937), .A2(new_n967), .A3(new_n941), .A4(KEYINPUT112), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n970), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n927), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n972), .A2(new_n937), .A3(new_n941), .A4(new_n973), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n932), .A2(new_n963), .A3(new_n966), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n979), .A2(new_n926), .A3(new_n980), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n981), .A2(new_n913), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT43), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n978), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n981), .A2(new_n913), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n926), .B1(new_n979), .B2(new_n980), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT43), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  XOR2_X1   g563(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n985), .A2(KEYINPUT43), .A3(new_n986), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n985), .B1(new_n927), .B2(new_n977), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT44), .B1(new_n992), .B2(new_n983), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n990), .B1(new_n991), .B2(new_n993), .ZN(G397));
  INV_X1    g569(.A(G1384), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(new_n496), .B2(new_n507), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n996), .A2(KEYINPUT113), .ZN(new_n997));
  AOI21_X1  g572(.A(G1384), .B1(new_n875), .B2(new_n876), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n997), .A2(new_n1000), .A3(KEYINPUT45), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n471), .A2(new_n477), .A3(new_n474), .A4(G40), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n1004), .A2(G1986), .A3(G290), .ZN(new_n1005));
  XOR2_X1   g580(.A(new_n1005), .B(KEYINPUT127), .Z(new_n1006));
  XNOR2_X1  g581(.A(new_n1006), .B(KEYINPUT48), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n704), .B(new_n707), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n1008), .B(KEYINPUT114), .ZN(new_n1009));
  INV_X1    g584(.A(G1996), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n770), .B(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n755), .B(new_n759), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1009), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1007), .B1(new_n1004), .B2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1004), .A2(G1996), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n1016), .A2(KEYINPUT46), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(KEYINPUT46), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1004), .B1(new_n771), .B2(new_n1012), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  XOR2_X1   g595(.A(new_n1020), .B(KEYINPUT47), .Z(new_n1021));
  NAND2_X1  g596(.A1(new_n705), .A2(new_n708), .ZN(new_n1022));
  OAI22_X1  g597(.A1(new_n1013), .A2(new_n1022), .B1(G2067), .B2(new_n755), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1023), .A2(new_n1003), .A3(new_n1001), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1015), .A2(new_n1021), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT116), .B1(new_n877), .B2(new_n995), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT116), .ZN(new_n1027));
  AOI211_X1 g602(.A(new_n1027), .B(G1384), .C1(new_n875), .C2(new_n876), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1003), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n1029), .A2(G8), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n603), .B1(new_n596), .B2(new_n511), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(G1981), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n599), .A2(new_n691), .A3(new_n603), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT49), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1032), .A2(KEYINPUT49), .A3(new_n1033), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1030), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G1976), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(new_n1039), .A3(new_n714), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n1033), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n1030), .ZN(new_n1042));
  INV_X1    g617(.A(G1971), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT45), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1003), .B1(new_n996), .B2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n998), .A2(KEYINPUT45), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1043), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT115), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT50), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1050), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1051));
  INV_X1    g626(.A(G2090), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1002), .B1(new_n996), .B2(KEYINPUT50), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1002), .B1(new_n998), .B2(KEYINPUT45), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1055), .B1(KEYINPUT45), .B2(new_n998), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(KEYINPUT115), .A3(new_n1043), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1049), .A2(new_n1054), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(G303), .A2(G8), .ZN(new_n1059));
  XNOR2_X1  g634(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n1059), .B(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1058), .A2(G8), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n714), .A2(G1976), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1029), .A2(G8), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n1066));
  NAND2_X1  g641(.A1(G288), .A2(new_n1039), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1029), .A2(G8), .A3(new_n1063), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT118), .B1(new_n1069), .B2(KEYINPUT52), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1029), .A2(new_n1066), .A3(G8), .A4(new_n1063), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1067), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1068), .B(new_n1038), .C1(new_n1070), .C2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1042), .B1(new_n1062), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT119), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1042), .B(new_n1077), .C1(new_n1062), .C2(new_n1074), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT63), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n996), .A2(new_n1027), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n998), .A2(KEYINPUT116), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1081), .A2(KEYINPUT50), .A3(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT120), .B1(new_n996), .B2(KEYINPUT50), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n998), .A2(new_n1085), .A3(new_n1050), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1083), .A2(new_n1003), .A3(new_n1084), .A4(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1047), .B1(new_n1087), .B2(G2090), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(G8), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1061), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n1071), .A2(KEYINPUT118), .A3(new_n1072), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1065), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1064), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1092), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1091), .A2(new_n1095), .A3(new_n1062), .A4(new_n1038), .ZN(new_n1096));
  INV_X1    g671(.A(G8), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1026), .A2(new_n1028), .A3(KEYINPUT45), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n819), .B1(new_n1098), .B2(new_n1045), .ZN(new_n1099));
  XOR2_X1   g674(.A(KEYINPUT121), .B(G2084), .Z(new_n1100));
  NAND3_X1  g675(.A1(new_n1051), .A2(new_n1053), .A3(new_n1100), .ZN(new_n1101));
  AOI211_X1 g676(.A(new_n1097), .B(G286), .C1(new_n1099), .C2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1080), .B1(new_n1096), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT122), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1095), .A2(new_n1062), .A3(new_n1038), .A4(new_n1102), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1058), .A2(G8), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1080), .B1(new_n1107), .B2(new_n1090), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1105), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n1058), .A2(G8), .A3(new_n1061), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1074), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1112), .A2(KEYINPUT122), .A3(new_n1102), .A4(new_n1108), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1104), .A2(new_n1110), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1079), .A2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1045), .B1(new_n1116), .B2(new_n1044), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1101), .B(G168), .C1(new_n1117), .C2(G1966), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(G8), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT51), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1118), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1121), .A2(KEYINPUT123), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1099), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1101), .ZN(new_n1125));
  OAI21_X1  g700(.A(G8), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  OR2_X1    g701(.A1(new_n1126), .A2(G168), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1119), .A2(new_n1128), .A3(new_n1120), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1123), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT62), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n1056), .A2(G2078), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT53), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1134));
  XOR2_X1   g709(.A(KEYINPUT125), .B(G1961), .Z(new_n1135));
  AOI22_X1  g710(.A1(new_n1132), .A2(new_n1133), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1098), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1045), .A2(G2078), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AND2_X1   g714(.A1(new_n1139), .A2(KEYINPUT124), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT53), .B1(new_n1139), .B2(KEYINPUT124), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1136), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n1142), .A2(G171), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1123), .A2(new_n1144), .A3(new_n1127), .A4(new_n1129), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1131), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT61), .ZN(new_n1147));
  XNOR2_X1  g722(.A(KEYINPUT56), .B(G2072), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1148), .ZN(new_n1149));
  NOR3_X1   g724(.A1(new_n1045), .A2(new_n1046), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT57), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n584), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n567), .A2(new_n573), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1153), .A2(KEYINPUT57), .A3(new_n581), .A4(new_n579), .ZN(new_n1154));
  AOI221_X4 g729(.A(new_n1150), .B1(new_n1152), .B2(new_n1154), .C1(new_n1087), .C2(new_n742), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1087), .A2(new_n742), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1150), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1156), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1147), .B1(new_n1155), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1156), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1002), .B1(new_n1116), .B2(KEYINPUT50), .ZN(new_n1162));
  AND2_X1   g737(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1163));
  AOI21_X1  g738(.A(G1956), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1161), .B1(new_n1164), .B2(new_n1150), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1157), .A2(new_n1156), .A3(new_n1158), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1165), .A2(KEYINPUT61), .A3(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1168));
  XOR2_X1   g743(.A(KEYINPUT58), .B(G1341), .Z(new_n1169));
  AOI22_X1  g744(.A1(new_n1168), .A2(new_n1010), .B1(new_n1029), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(KEYINPUT59), .B1(new_n1170), .B2(new_n841), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT59), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n1029), .A2(new_n1169), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1056), .A2(G1996), .ZN(new_n1174));
  OAI211_X1 g749(.A(new_n1172), .B(new_n554), .C1(new_n1173), .C2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n798), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1176));
  OAI211_X1 g751(.A(new_n759), .B(new_n1003), .C1(new_n1026), .C2(new_n1028), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1177), .ZN(new_n1178));
  NOR3_X1   g753(.A1(new_n1176), .A2(new_n1178), .A3(KEYINPUT60), .ZN(new_n1179));
  AOI22_X1  g754(.A1(new_n1171), .A2(new_n1175), .B1(new_n1179), .B2(new_n617), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1176), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n938), .B1(new_n1181), .B2(new_n1177), .ZN(new_n1182));
  NOR3_X1   g757(.A1(new_n1176), .A2(new_n1178), .A3(new_n617), .ZN(new_n1183));
  OAI21_X1  g758(.A(KEYINPUT60), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1160), .A2(new_n1167), .A3(new_n1180), .A4(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1166), .B1(new_n1159), .B2(new_n1182), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g762(.A(G301), .B(KEYINPUT54), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1142), .A2(new_n1188), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n1001), .A2(new_n1133), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1190), .A2(new_n1138), .ZN(new_n1191));
  XOR2_X1   g766(.A(new_n1191), .B(KEYINPUT126), .Z(new_n1192));
  INV_X1    g767(.A(new_n1188), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1192), .A2(new_n1136), .A3(new_n1193), .ZN(new_n1194));
  NAND4_X1  g769(.A1(new_n1187), .A2(new_n1130), .A3(new_n1189), .A4(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1146), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1096), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1115), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  XOR2_X1   g773(.A(G290), .B(G1986), .Z(new_n1199));
  AOI21_X1  g774(.A(new_n1004), .B1(new_n1014), .B2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1025), .B1(new_n1198), .B2(new_n1200), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g776(.A(G229), .ZN(new_n1203));
  AND3_X1   g777(.A1(new_n917), .A2(new_n918), .A3(new_n914), .ZN(new_n1204));
  AOI21_X1  g778(.A(new_n918), .B1(new_n917), .B2(new_n914), .ZN(new_n1205));
  OAI211_X1 g779(.A(new_n661), .B(new_n1203), .C1(new_n1204), .C2(new_n1205), .ZN(new_n1206));
  INV_X1    g780(.A(G227), .ZN(new_n1207));
  NAND3_X1  g781(.A1(new_n988), .A2(G319), .A3(new_n1207), .ZN(new_n1208));
  NOR2_X1   g782(.A1(new_n1206), .A2(new_n1208), .ZN(G308));
  INV_X1    g783(.A(new_n661), .ZN(new_n1210));
  AOI21_X1  g784(.A(new_n1210), .B1(new_n916), .B2(new_n919), .ZN(new_n1211));
  AOI21_X1  g785(.A(new_n461), .B1(new_n984), .B2(new_n987), .ZN(new_n1212));
  NAND4_X1  g786(.A1(new_n1211), .A2(new_n1207), .A3(new_n1203), .A4(new_n1212), .ZN(G225));
endmodule


