

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U549 ( .A(n517), .B(KEYINPUT65), .ZN(n984) );
  INV_X1 U550 ( .A(n738), .ZN(n729) );
  XNOR2_X1 U551 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U552 ( .A(G2104), .B(KEYINPUT64), .Z(n514) );
  NOR2_X1 U553 ( .A1(n730), .A2(n729), .ZN(n515) );
  OR2_X1 U554 ( .A1(n695), .A2(n694), .ZN(n516) );
  INV_X1 U555 ( .A(KEYINPUT87), .ZN(n640) );
  NAND2_X1 U556 ( .A1(n642), .A2(G8), .ZN(n643) );
  XNOR2_X1 U557 ( .A(n643), .B(KEYINPUT30), .ZN(n644) );
  INV_X1 U558 ( .A(KEYINPUT29), .ZN(n634) );
  NOR2_X1 U559 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U560 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U561 ( .A(n665), .B(KEYINPUT89), .ZN(n666) );
  INV_X1 U562 ( .A(KEYINPUT17), .ZN(n518) );
  XNOR2_X1 U563 ( .A(n518), .B(KEYINPUT66), .ZN(n519) );
  BUF_X1 U564 ( .A(n527), .Z(n988) );
  INV_X1 U565 ( .A(KEYINPUT23), .ZN(n528) );
  INV_X1 U566 ( .A(KEYINPUT40), .ZN(n747) );
  NOR2_X1 U567 ( .A1(G651), .A2(n572), .ZN(n781) );
  XNOR2_X1 U568 ( .A(n747), .B(KEYINPUT97), .ZN(n748) );
  NAND2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n517) );
  NAND2_X1 U570 ( .A1(G114), .A2(n984), .ZN(n522) );
  NOR2_X1 U571 ( .A1(G2105), .A2(G2104), .ZN(n520) );
  XNOR2_X2 U572 ( .A(n520), .B(n519), .ZN(n698) );
  NAND2_X1 U573 ( .A1(G138), .A2(n698), .ZN(n521) );
  NAND2_X1 U574 ( .A1(n522), .A2(n521), .ZN(n526) );
  AND2_X1 U575 ( .A1(n514), .A2(G2105), .ZN(n985) );
  NAND2_X1 U576 ( .A1(G126), .A2(n985), .ZN(n524) );
  NOR2_X1 U577 ( .A1(n514), .A2(G2105), .ZN(n527) );
  NAND2_X1 U578 ( .A1(G102), .A2(n988), .ZN(n523) );
  NAND2_X1 U579 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X1 U580 ( .A1(n526), .A2(n525), .ZN(G164) );
  NAND2_X1 U581 ( .A1(n984), .A2(G113), .ZN(n531) );
  NAND2_X1 U582 ( .A1(G101), .A2(n527), .ZN(n529) );
  NAND2_X1 U583 ( .A1(n531), .A2(n530), .ZN(n535) );
  NAND2_X1 U584 ( .A1(n985), .A2(G125), .ZN(n533) );
  NAND2_X1 U585 ( .A1(G137), .A2(n698), .ZN(n532) );
  NAND2_X1 U586 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X2 U587 ( .A1(n535), .A2(n534), .ZN(G160) );
  NOR2_X1 U588 ( .A1(G543), .A2(G651), .ZN(n778) );
  NAND2_X1 U589 ( .A1(n778), .A2(G89), .ZN(n536) );
  XNOR2_X1 U590 ( .A(n536), .B(KEYINPUT4), .ZN(n538) );
  XOR2_X1 U591 ( .A(G543), .B(KEYINPUT0), .Z(n572) );
  INV_X1 U592 ( .A(G651), .ZN(n540) );
  NOR2_X1 U593 ( .A1(n572), .A2(n540), .ZN(n782) );
  NAND2_X1 U594 ( .A1(G76), .A2(n782), .ZN(n537) );
  NAND2_X1 U595 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U596 ( .A(n539), .B(KEYINPUT5), .ZN(n546) );
  NOR2_X1 U597 ( .A1(G543), .A2(n540), .ZN(n541) );
  XOR2_X1 U598 ( .A(KEYINPUT1), .B(n541), .Z(n777) );
  NAND2_X1 U599 ( .A1(G63), .A2(n777), .ZN(n543) );
  NAND2_X1 U600 ( .A1(G51), .A2(n781), .ZN(n542) );
  NAND2_X1 U601 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U602 ( .A(KEYINPUT6), .B(n544), .Z(n545) );
  NAND2_X1 U603 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U604 ( .A(n547), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U605 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U606 ( .A1(G78), .A2(n782), .ZN(n549) );
  NAND2_X1 U607 ( .A1(G91), .A2(n778), .ZN(n548) );
  NAND2_X1 U608 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U609 ( .A(KEYINPUT70), .B(n550), .ZN(n553) );
  NAND2_X1 U610 ( .A1(G53), .A2(n781), .ZN(n551) );
  XNOR2_X1 U611 ( .A(KEYINPUT71), .B(n551), .ZN(n552) );
  NOR2_X1 U612 ( .A1(n553), .A2(n552), .ZN(n555) );
  NAND2_X1 U613 ( .A1(n777), .A2(G65), .ZN(n554) );
  NAND2_X1 U614 ( .A1(n555), .A2(n554), .ZN(G299) );
  NAND2_X1 U615 ( .A1(G64), .A2(n777), .ZN(n557) );
  NAND2_X1 U616 ( .A1(G52), .A2(n781), .ZN(n556) );
  NAND2_X1 U617 ( .A1(n557), .A2(n556), .ZN(n562) );
  NAND2_X1 U618 ( .A1(G77), .A2(n782), .ZN(n559) );
  NAND2_X1 U619 ( .A1(G90), .A2(n778), .ZN(n558) );
  NAND2_X1 U620 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U621 ( .A(KEYINPUT9), .B(n560), .Z(n561) );
  NOR2_X1 U622 ( .A1(n562), .A2(n561), .ZN(G171) );
  INV_X1 U623 ( .A(G171), .ZN(G301) );
  NAND2_X1 U624 ( .A1(G75), .A2(n782), .ZN(n564) );
  NAND2_X1 U625 ( .A1(G88), .A2(n778), .ZN(n563) );
  NAND2_X1 U626 ( .A1(n564), .A2(n563), .ZN(n568) );
  NAND2_X1 U627 ( .A1(G62), .A2(n777), .ZN(n566) );
  NAND2_X1 U628 ( .A1(G50), .A2(n781), .ZN(n565) );
  NAND2_X1 U629 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U630 ( .A1(n568), .A2(n567), .ZN(G166) );
  INV_X1 U631 ( .A(G166), .ZN(G303) );
  NAND2_X1 U632 ( .A1(G49), .A2(n781), .ZN(n570) );
  NAND2_X1 U633 ( .A1(G74), .A2(G651), .ZN(n569) );
  NAND2_X1 U634 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U635 ( .A1(n777), .A2(n571), .ZN(n574) );
  NAND2_X1 U636 ( .A1(n572), .A2(G87), .ZN(n573) );
  NAND2_X1 U637 ( .A1(n574), .A2(n573), .ZN(G288) );
  NAND2_X1 U638 ( .A1(G61), .A2(n777), .ZN(n576) );
  NAND2_X1 U639 ( .A1(G86), .A2(n778), .ZN(n575) );
  NAND2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n579) );
  NAND2_X1 U641 ( .A1(n782), .A2(G73), .ZN(n577) );
  XOR2_X1 U642 ( .A(KEYINPUT2), .B(n577), .Z(n578) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n581) );
  NAND2_X1 U644 ( .A1(n781), .A2(G48), .ZN(n580) );
  NAND2_X1 U645 ( .A1(n581), .A2(n580), .ZN(G305) );
  NAND2_X1 U646 ( .A1(n782), .A2(G72), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(KEYINPUT68), .ZN(n590) );
  NAND2_X1 U648 ( .A1(G60), .A2(n777), .ZN(n584) );
  NAND2_X1 U649 ( .A1(G47), .A2(n781), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U651 ( .A(KEYINPUT69), .B(n585), .Z(n588) );
  NAND2_X1 U652 ( .A1(G85), .A2(n778), .ZN(n586) );
  XNOR2_X1 U653 ( .A(KEYINPUT67), .B(n586), .ZN(n587) );
  NOR2_X1 U654 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U655 ( .A1(n590), .A2(n589), .ZN(G290) );
  NOR2_X2 U656 ( .A1(G164), .A2(G1384), .ZN(n714) );
  NAND2_X1 U657 ( .A1(G160), .A2(G40), .ZN(n715) );
  INV_X1 U658 ( .A(n715), .ZN(n591) );
  NAND2_X2 U659 ( .A1(n714), .A2(n591), .ZN(n653) );
  INV_X1 U660 ( .A(n653), .ZN(n592) );
  NAND2_X1 U661 ( .A1(n592), .A2(G1996), .ZN(n593) );
  XNOR2_X1 U662 ( .A(n593), .B(KEYINPUT26), .ZN(n595) );
  NAND2_X1 U663 ( .A1(G1341), .A2(n653), .ZN(n594) );
  NAND2_X1 U664 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U665 ( .A(KEYINPUT85), .B(n596), .Z(n607) );
  NAND2_X1 U666 ( .A1(n777), .A2(G56), .ZN(n597) );
  XNOR2_X1 U667 ( .A(KEYINPUT14), .B(n597), .ZN(n603) );
  NAND2_X1 U668 ( .A1(n778), .A2(G81), .ZN(n598) );
  XNOR2_X1 U669 ( .A(n598), .B(KEYINPUT12), .ZN(n600) );
  NAND2_X1 U670 ( .A1(G68), .A2(n782), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U672 ( .A(KEYINPUT13), .B(n601), .ZN(n602) );
  NAND2_X1 U673 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U674 ( .A(n604), .B(KEYINPUT73), .ZN(n606) );
  NAND2_X1 U675 ( .A1(n781), .A2(G43), .ZN(n605) );
  NAND2_X1 U676 ( .A1(n606), .A2(n605), .ZN(n907) );
  NOR2_X1 U677 ( .A1(n607), .A2(n907), .ZN(n621) );
  NAND2_X1 U678 ( .A1(G54), .A2(n781), .ZN(n609) );
  NAND2_X1 U679 ( .A1(G79), .A2(n782), .ZN(n608) );
  NAND2_X1 U680 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U681 ( .A(KEYINPUT74), .B(n610), .ZN(n614) );
  NAND2_X1 U682 ( .A1(G66), .A2(n777), .ZN(n612) );
  NAND2_X1 U683 ( .A1(G92), .A2(n778), .ZN(n611) );
  NAND2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U685 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U686 ( .A(KEYINPUT15), .B(n615), .Z(n1009) );
  NAND2_X1 U687 ( .A1(n621), .A2(n1009), .ZN(n620) );
  NAND2_X1 U688 ( .A1(G1348), .A2(n653), .ZN(n617) );
  NAND2_X1 U689 ( .A1(G2067), .A2(n592), .ZN(n616) );
  NAND2_X1 U690 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U691 ( .A(KEYINPUT86), .B(n618), .ZN(n619) );
  NAND2_X1 U692 ( .A1(n620), .A2(n619), .ZN(n623) );
  OR2_X1 U693 ( .A1(n1009), .A2(n621), .ZN(n622) );
  NAND2_X1 U694 ( .A1(n623), .A2(n622), .ZN(n629) );
  INV_X1 U695 ( .A(G299), .ZN(n794) );
  NAND2_X1 U696 ( .A1(G2072), .A2(n592), .ZN(n624) );
  XNOR2_X1 U697 ( .A(n624), .B(KEYINPUT84), .ZN(n625) );
  XNOR2_X1 U698 ( .A(KEYINPUT27), .B(n625), .ZN(n627) );
  AND2_X1 U699 ( .A1(n653), .A2(G1956), .ZN(n626) );
  NOR2_X1 U700 ( .A1(n627), .A2(n626), .ZN(n630) );
  NAND2_X1 U701 ( .A1(n794), .A2(n630), .ZN(n628) );
  NAND2_X1 U702 ( .A1(n629), .A2(n628), .ZN(n633) );
  NOR2_X1 U703 ( .A1(n794), .A2(n630), .ZN(n631) );
  XOR2_X1 U704 ( .A(n631), .B(KEYINPUT28), .Z(n632) );
  NAND2_X1 U705 ( .A1(n633), .A2(n632), .ZN(n635) );
  XNOR2_X1 U706 ( .A(n635), .B(n634), .ZN(n639) );
  NAND2_X1 U707 ( .A1(G1961), .A2(n653), .ZN(n637) );
  XOR2_X1 U708 ( .A(G2078), .B(KEYINPUT25), .Z(n833) );
  NAND2_X1 U709 ( .A1(n592), .A2(n833), .ZN(n636) );
  NAND2_X1 U710 ( .A1(n637), .A2(n636), .ZN(n645) );
  OR2_X1 U711 ( .A1(G301), .A2(n645), .ZN(n638) );
  NAND2_X1 U712 ( .A1(n639), .A2(n638), .ZN(n651) );
  NOR2_X1 U713 ( .A1(G2084), .A2(n653), .ZN(n661) );
  NAND2_X1 U714 ( .A1(G8), .A2(n653), .ZN(n694) );
  NOR2_X1 U715 ( .A1(G1966), .A2(n694), .ZN(n662) );
  NOR2_X1 U716 ( .A1(n661), .A2(n662), .ZN(n641) );
  XNOR2_X1 U717 ( .A(n641), .B(n640), .ZN(n642) );
  NOR2_X1 U718 ( .A1(G168), .A2(n644), .ZN(n648) );
  NAND2_X1 U719 ( .A1(G301), .A2(n645), .ZN(n646) );
  XOR2_X1 U720 ( .A(KEYINPUT88), .B(n646), .Z(n647) );
  XOR2_X1 U721 ( .A(KEYINPUT31), .B(n649), .Z(n650) );
  NAND2_X1 U722 ( .A1(n651), .A2(n650), .ZN(n664) );
  NAND2_X1 U723 ( .A1(n664), .A2(G286), .ZN(n658) );
  NOR2_X1 U724 ( .A1(G1971), .A2(n694), .ZN(n652) );
  XNOR2_X1 U725 ( .A(n652), .B(KEYINPUT90), .ZN(n655) );
  NOR2_X1 U726 ( .A1(n653), .A2(G2090), .ZN(n654) );
  NOR2_X1 U727 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U728 ( .A1(n656), .A2(G303), .ZN(n657) );
  NAND2_X1 U729 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U730 ( .A1(n659), .A2(G8), .ZN(n660) );
  XNOR2_X1 U731 ( .A(n660), .B(KEYINPUT32), .ZN(n669) );
  NAND2_X1 U732 ( .A1(G8), .A2(n661), .ZN(n667) );
  INV_X1 U733 ( .A(n662), .ZN(n663) );
  NAND2_X1 U734 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U735 ( .A1(n669), .A2(n668), .ZN(n685) );
  NOR2_X1 U736 ( .A1(G1976), .A2(G288), .ZN(n679) );
  NOR2_X1 U737 ( .A1(G1971), .A2(G303), .ZN(n670) );
  NOR2_X1 U738 ( .A1(n679), .A2(n670), .ZN(n895) );
  INV_X1 U739 ( .A(KEYINPUT33), .ZN(n671) );
  AND2_X1 U740 ( .A1(n895), .A2(n671), .ZN(n672) );
  NAND2_X1 U741 ( .A1(n685), .A2(n672), .ZN(n676) );
  INV_X1 U742 ( .A(n694), .ZN(n673) );
  NAND2_X1 U743 ( .A1(G1976), .A2(G288), .ZN(n894) );
  AND2_X1 U744 ( .A1(n673), .A2(n894), .ZN(n674) );
  OR2_X1 U745 ( .A1(KEYINPUT33), .A2(n674), .ZN(n675) );
  NAND2_X1 U746 ( .A1(n676), .A2(n675), .ZN(n678) );
  INV_X1 U747 ( .A(KEYINPUT91), .ZN(n677) );
  XNOR2_X1 U748 ( .A(n678), .B(n677), .ZN(n682) );
  NAND2_X1 U749 ( .A1(n679), .A2(KEYINPUT33), .ZN(n680) );
  NOR2_X1 U750 ( .A1(n694), .A2(n680), .ZN(n681) );
  NOR2_X2 U751 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U752 ( .A(n683), .B(KEYINPUT92), .ZN(n684) );
  XOR2_X1 U753 ( .A(G1981), .B(G305), .Z(n890) );
  NAND2_X1 U754 ( .A1(n684), .A2(n890), .ZN(n690) );
  NOR2_X1 U755 ( .A1(G2090), .A2(G303), .ZN(n686) );
  NAND2_X1 U756 ( .A1(G8), .A2(n686), .ZN(n687) );
  NAND2_X1 U757 ( .A1(n685), .A2(n687), .ZN(n688) );
  NAND2_X1 U758 ( .A1(n688), .A2(n694), .ZN(n689) );
  NAND2_X1 U759 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U760 ( .A(n691), .B(KEYINPUT93), .ZN(n696) );
  NOR2_X1 U761 ( .A1(G1981), .A2(G305), .ZN(n692) );
  XNOR2_X1 U762 ( .A(n692), .B(KEYINPUT24), .ZN(n693) );
  XNOR2_X1 U763 ( .A(n693), .B(KEYINPUT83), .ZN(n695) );
  NAND2_X1 U764 ( .A1(n696), .A2(n516), .ZN(n731) );
  NAND2_X1 U765 ( .A1(G105), .A2(n988), .ZN(n697) );
  XNOR2_X1 U766 ( .A(n697), .B(KEYINPUT38), .ZN(n705) );
  NAND2_X1 U767 ( .A1(n985), .A2(G129), .ZN(n700) );
  NAND2_X1 U768 ( .A1(G141), .A2(n698), .ZN(n699) );
  NAND2_X1 U769 ( .A1(n700), .A2(n699), .ZN(n703) );
  NAND2_X1 U770 ( .A1(G117), .A2(n984), .ZN(n701) );
  XNOR2_X1 U771 ( .A(KEYINPUT81), .B(n701), .ZN(n702) );
  NOR2_X1 U772 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U773 ( .A1(n705), .A2(n704), .ZN(n979) );
  NAND2_X1 U774 ( .A1(G1996), .A2(n979), .ZN(n713) );
  NAND2_X1 U775 ( .A1(G107), .A2(n984), .ZN(n707) );
  NAND2_X1 U776 ( .A1(G119), .A2(n985), .ZN(n706) );
  NAND2_X1 U777 ( .A1(n707), .A2(n706), .ZN(n711) );
  NAND2_X1 U778 ( .A1(n988), .A2(G95), .ZN(n709) );
  NAND2_X1 U779 ( .A1(G131), .A2(n698), .ZN(n708) );
  NAND2_X1 U780 ( .A1(n709), .A2(n708), .ZN(n710) );
  OR2_X1 U781 ( .A1(n711), .A2(n710), .ZN(n994) );
  NAND2_X1 U782 ( .A1(G1991), .A2(n994), .ZN(n712) );
  NAND2_X1 U783 ( .A1(n713), .A2(n712), .ZN(n854) );
  NOR2_X1 U784 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U785 ( .A(n716), .B(KEYINPUT80), .ZN(n743) );
  NAND2_X1 U786 ( .A1(n854), .A2(n743), .ZN(n717) );
  XNOR2_X1 U787 ( .A(n717), .B(KEYINPUT82), .ZN(n719) );
  XNOR2_X1 U788 ( .A(G1986), .B(G290), .ZN(n899) );
  NAND2_X1 U789 ( .A1(n899), .A2(n743), .ZN(n718) );
  NAND2_X1 U790 ( .A1(n719), .A2(n718), .ZN(n730) );
  NAND2_X1 U791 ( .A1(n988), .A2(G104), .ZN(n721) );
  NAND2_X1 U792 ( .A1(G140), .A2(n698), .ZN(n720) );
  NAND2_X1 U793 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U794 ( .A(KEYINPUT34), .B(n722), .ZN(n727) );
  NAND2_X1 U795 ( .A1(G116), .A2(n984), .ZN(n724) );
  NAND2_X1 U796 ( .A1(G128), .A2(n985), .ZN(n723) );
  NAND2_X1 U797 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U798 ( .A(KEYINPUT35), .B(n725), .Z(n726) );
  NOR2_X1 U799 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U800 ( .A(KEYINPUT36), .B(n728), .ZN(n1003) );
  XNOR2_X1 U801 ( .A(G2067), .B(KEYINPUT37), .ZN(n741) );
  NOR2_X1 U802 ( .A1(n1003), .A2(n741), .ZN(n874) );
  NAND2_X1 U803 ( .A1(n874), .A2(n743), .ZN(n738) );
  NAND2_X1 U804 ( .A1(n731), .A2(n515), .ZN(n746) );
  NOR2_X1 U805 ( .A1(G1996), .A2(n979), .ZN(n851) );
  NOR2_X1 U806 ( .A1(G1986), .A2(G290), .ZN(n732) );
  NOR2_X1 U807 ( .A1(G1991), .A2(n994), .ZN(n873) );
  NOR2_X1 U808 ( .A1(n732), .A2(n873), .ZN(n733) );
  XNOR2_X1 U809 ( .A(n733), .B(KEYINPUT94), .ZN(n734) );
  NOR2_X1 U810 ( .A1(n854), .A2(n734), .ZN(n735) );
  XOR2_X1 U811 ( .A(KEYINPUT95), .B(n735), .Z(n736) );
  NOR2_X1 U812 ( .A1(n851), .A2(n736), .ZN(n737) );
  XNOR2_X1 U813 ( .A(KEYINPUT39), .B(n737), .ZN(n739) );
  NAND2_X1 U814 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U815 ( .A(n740), .B(KEYINPUT96), .ZN(n742) );
  NAND2_X1 U816 ( .A1(n1003), .A2(n741), .ZN(n855) );
  NAND2_X1 U817 ( .A1(n742), .A2(n855), .ZN(n744) );
  NAND2_X1 U818 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U819 ( .A1(n746), .A2(n745), .ZN(n749) );
  XNOR2_X1 U820 ( .A(n749), .B(n748), .ZN(G329) );
  AND2_X1 U821 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U822 ( .A(G57), .ZN(G237) );
  INV_X1 U823 ( .A(G132), .ZN(G219) );
  INV_X1 U824 ( .A(G82), .ZN(G220) );
  NAND2_X1 U825 ( .A1(G7), .A2(G661), .ZN(n750) );
  XNOR2_X1 U826 ( .A(n750), .B(KEYINPUT10), .ZN(n751) );
  XNOR2_X1 U827 ( .A(KEYINPUT72), .B(n751), .ZN(G223) );
  INV_X1 U828 ( .A(G223), .ZN(n814) );
  NAND2_X1 U829 ( .A1(n814), .A2(G567), .ZN(n752) );
  XOR2_X1 U830 ( .A(KEYINPUT11), .B(n752), .Z(G234) );
  INV_X1 U831 ( .A(G860), .ZN(n757) );
  OR2_X1 U832 ( .A1(n907), .A2(n757), .ZN(G153) );
  NAND2_X1 U833 ( .A1(G868), .A2(G301), .ZN(n754) );
  OR2_X1 U834 ( .A1(n1009), .A2(G868), .ZN(n753) );
  NAND2_X1 U835 ( .A1(n754), .A2(n753), .ZN(G284) );
  INV_X1 U836 ( .A(G868), .ZN(n797) );
  NOR2_X1 U837 ( .A1(G286), .A2(n797), .ZN(n756) );
  NOR2_X1 U838 ( .A1(G868), .A2(G299), .ZN(n755) );
  NOR2_X1 U839 ( .A1(n756), .A2(n755), .ZN(G297) );
  NAND2_X1 U840 ( .A1(n757), .A2(G559), .ZN(n758) );
  NAND2_X1 U841 ( .A1(n758), .A2(n1009), .ZN(n759) );
  XNOR2_X1 U842 ( .A(n759), .B(KEYINPUT16), .ZN(n760) );
  XOR2_X1 U843 ( .A(KEYINPUT75), .B(n760), .Z(G148) );
  NOR2_X1 U844 ( .A1(G868), .A2(n907), .ZN(n763) );
  NAND2_X1 U845 ( .A1(G868), .A2(n1009), .ZN(n761) );
  NOR2_X1 U846 ( .A1(G559), .A2(n761), .ZN(n762) );
  NOR2_X1 U847 ( .A1(n763), .A2(n762), .ZN(G282) );
  NAND2_X1 U848 ( .A1(G123), .A2(n985), .ZN(n764) );
  XNOR2_X1 U849 ( .A(n764), .B(KEYINPUT76), .ZN(n765) );
  XNOR2_X1 U850 ( .A(KEYINPUT18), .B(n765), .ZN(n770) );
  NAND2_X1 U851 ( .A1(G111), .A2(n984), .ZN(n767) );
  NAND2_X1 U852 ( .A1(G99), .A2(n988), .ZN(n766) );
  NAND2_X1 U853 ( .A1(n767), .A2(n766), .ZN(n768) );
  XOR2_X1 U854 ( .A(KEYINPUT78), .B(n768), .Z(n769) );
  NAND2_X1 U855 ( .A1(n770), .A2(n769), .ZN(n773) );
  NAND2_X1 U856 ( .A1(G135), .A2(n698), .ZN(n771) );
  XNOR2_X1 U857 ( .A(KEYINPUT77), .B(n771), .ZN(n772) );
  NOR2_X1 U858 ( .A1(n773), .A2(n772), .ZN(n977) );
  XNOR2_X1 U859 ( .A(n977), .B(G2096), .ZN(n775) );
  INV_X1 U860 ( .A(G2100), .ZN(n774) );
  NAND2_X1 U861 ( .A1(n775), .A2(n774), .ZN(G156) );
  NAND2_X1 U862 ( .A1(n1009), .A2(G559), .ZN(n795) );
  XNOR2_X1 U863 ( .A(n907), .B(n795), .ZN(n776) );
  NOR2_X1 U864 ( .A1(n776), .A2(G860), .ZN(n787) );
  NAND2_X1 U865 ( .A1(G67), .A2(n777), .ZN(n780) );
  NAND2_X1 U866 ( .A1(G93), .A2(n778), .ZN(n779) );
  NAND2_X1 U867 ( .A1(n780), .A2(n779), .ZN(n786) );
  NAND2_X1 U868 ( .A1(G55), .A2(n781), .ZN(n784) );
  NAND2_X1 U869 ( .A1(G80), .A2(n782), .ZN(n783) );
  NAND2_X1 U870 ( .A1(n784), .A2(n783), .ZN(n785) );
  OR2_X1 U871 ( .A1(n786), .A2(n785), .ZN(n798) );
  XOR2_X1 U872 ( .A(n787), .B(n798), .Z(G145) );
  XOR2_X1 U873 ( .A(n798), .B(G290), .Z(n788) );
  XNOR2_X1 U874 ( .A(n788), .B(G288), .ZN(n789) );
  XNOR2_X1 U875 ( .A(KEYINPUT19), .B(n789), .ZN(n791) );
  XNOR2_X1 U876 ( .A(G305), .B(G166), .ZN(n790) );
  XNOR2_X1 U877 ( .A(n791), .B(n790), .ZN(n792) );
  XNOR2_X1 U878 ( .A(n792), .B(n907), .ZN(n793) );
  XNOR2_X1 U879 ( .A(n794), .B(n793), .ZN(n1007) );
  XNOR2_X1 U880 ( .A(n795), .B(n1007), .ZN(n796) );
  NAND2_X1 U881 ( .A1(n796), .A2(G868), .ZN(n800) );
  NAND2_X1 U882 ( .A1(n798), .A2(n797), .ZN(n799) );
  NAND2_X1 U883 ( .A1(n800), .A2(n799), .ZN(G295) );
  NAND2_X1 U884 ( .A1(G2084), .A2(G2078), .ZN(n801) );
  XOR2_X1 U885 ( .A(KEYINPUT20), .B(n801), .Z(n802) );
  NAND2_X1 U886 ( .A1(G2090), .A2(n802), .ZN(n803) );
  XNOR2_X1 U887 ( .A(KEYINPUT21), .B(n803), .ZN(n804) );
  NAND2_X1 U888 ( .A1(n804), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U889 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U890 ( .A1(G220), .A2(G219), .ZN(n805) );
  XOR2_X1 U891 ( .A(KEYINPUT22), .B(n805), .Z(n806) );
  NOR2_X1 U892 ( .A1(G218), .A2(n806), .ZN(n807) );
  NAND2_X1 U893 ( .A1(G96), .A2(n807), .ZN(n944) );
  NAND2_X1 U894 ( .A1(n944), .A2(G2106), .ZN(n811) );
  NAND2_X1 U895 ( .A1(G120), .A2(G108), .ZN(n808) );
  NOR2_X1 U896 ( .A1(G237), .A2(n808), .ZN(n809) );
  NAND2_X1 U897 ( .A1(G69), .A2(n809), .ZN(n945) );
  NAND2_X1 U898 ( .A1(n945), .A2(G567), .ZN(n810) );
  NAND2_X1 U899 ( .A1(n811), .A2(n810), .ZN(n956) );
  NAND2_X1 U900 ( .A1(G483), .A2(G661), .ZN(n812) );
  NOR2_X1 U901 ( .A1(n956), .A2(n812), .ZN(n818) );
  NAND2_X1 U902 ( .A1(n818), .A2(G36), .ZN(n813) );
  XOR2_X1 U903 ( .A(KEYINPUT79), .B(n813), .Z(G176) );
  NAND2_X1 U904 ( .A1(G2106), .A2(n814), .ZN(G217) );
  NAND2_X1 U905 ( .A1(G15), .A2(G2), .ZN(n816) );
  INV_X1 U906 ( .A(G661), .ZN(n815) );
  NOR2_X1 U907 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U908 ( .A(n817), .B(KEYINPUT99), .ZN(G259) );
  NAND2_X1 U909 ( .A1(G3), .A2(G1), .ZN(n819) );
  NAND2_X1 U910 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U911 ( .A(n820), .B(KEYINPUT100), .ZN(G188) );
  XOR2_X1 U912 ( .A(G108), .B(KEYINPUT114), .Z(G238) );
  NAND2_X1 U914 ( .A1(G124), .A2(n985), .ZN(n821) );
  XNOR2_X1 U915 ( .A(n821), .B(KEYINPUT44), .ZN(n824) );
  NAND2_X1 U916 ( .A1(n698), .A2(G136), .ZN(n822) );
  XNOR2_X1 U917 ( .A(n822), .B(KEYINPUT104), .ZN(n823) );
  NAND2_X1 U918 ( .A1(n824), .A2(n823), .ZN(n828) );
  NAND2_X1 U919 ( .A1(G112), .A2(n984), .ZN(n826) );
  NAND2_X1 U920 ( .A1(G100), .A2(n988), .ZN(n825) );
  NAND2_X1 U921 ( .A1(n826), .A2(n825), .ZN(n827) );
  NOR2_X1 U922 ( .A1(n828), .A2(n827), .ZN(G162) );
  XOR2_X1 U923 ( .A(G1996), .B(G32), .Z(n829) );
  NAND2_X1 U924 ( .A1(n829), .A2(G28), .ZN(n832) );
  XNOR2_X1 U925 ( .A(G25), .B(G1991), .ZN(n830) );
  XNOR2_X1 U926 ( .A(KEYINPUT120), .B(n830), .ZN(n831) );
  NOR2_X1 U927 ( .A1(n832), .A2(n831), .ZN(n840) );
  XNOR2_X1 U928 ( .A(n833), .B(G27), .ZN(n838) );
  XNOR2_X1 U929 ( .A(G2067), .B(G26), .ZN(n835) );
  XNOR2_X1 U930 ( .A(G2072), .B(G33), .ZN(n834) );
  NOR2_X1 U931 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U932 ( .A(KEYINPUT121), .B(n836), .ZN(n837) );
  NOR2_X1 U933 ( .A1(n838), .A2(n837), .ZN(n839) );
  NAND2_X1 U934 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U935 ( .A(n841), .B(KEYINPUT53), .ZN(n844) );
  XOR2_X1 U936 ( .A(G2084), .B(G34), .Z(n842) );
  XNOR2_X1 U937 ( .A(KEYINPUT54), .B(n842), .ZN(n843) );
  NAND2_X1 U938 ( .A1(n844), .A2(n843), .ZN(n846) );
  XNOR2_X1 U939 ( .A(G35), .B(G2090), .ZN(n845) );
  NOR2_X1 U940 ( .A1(n846), .A2(n845), .ZN(n847) );
  XNOR2_X1 U941 ( .A(KEYINPUT122), .B(n847), .ZN(n848) );
  NOR2_X1 U942 ( .A1(G29), .A2(n848), .ZN(n849) );
  XNOR2_X1 U943 ( .A(n849), .B(KEYINPUT55), .ZN(n888) );
  XOR2_X1 U944 ( .A(G2090), .B(G162), .Z(n850) );
  NOR2_X1 U945 ( .A1(n851), .A2(n850), .ZN(n852) );
  XOR2_X1 U946 ( .A(KEYINPUT51), .B(n852), .Z(n853) );
  XNOR2_X1 U947 ( .A(KEYINPUT116), .B(n853), .ZN(n883) );
  INV_X1 U948 ( .A(n854), .ZN(n856) );
  NAND2_X1 U949 ( .A1(n856), .A2(n855), .ZN(n881) );
  XNOR2_X1 U950 ( .A(G164), .B(G2078), .ZN(n857) );
  XNOR2_X1 U951 ( .A(n857), .B(KEYINPUT117), .ZN(n869) );
  NAND2_X1 U952 ( .A1(n988), .A2(G103), .ZN(n859) );
  NAND2_X1 U953 ( .A1(G139), .A2(n698), .ZN(n858) );
  NAND2_X1 U954 ( .A1(n859), .A2(n858), .ZN(n866) );
  NAND2_X1 U955 ( .A1(n984), .A2(G115), .ZN(n860) );
  XNOR2_X1 U956 ( .A(n860), .B(KEYINPUT106), .ZN(n862) );
  NAND2_X1 U957 ( .A1(G127), .A2(n985), .ZN(n861) );
  NAND2_X1 U958 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U959 ( .A(KEYINPUT107), .B(n863), .ZN(n864) );
  XNOR2_X1 U960 ( .A(KEYINPUT47), .B(n864), .ZN(n865) );
  NOR2_X1 U961 ( .A1(n866), .A2(n865), .ZN(n867) );
  XOR2_X1 U962 ( .A(KEYINPUT108), .B(n867), .Z(n1001) );
  XNOR2_X1 U963 ( .A(n1001), .B(G2072), .ZN(n868) );
  NOR2_X1 U964 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U965 ( .A(KEYINPUT118), .B(n870), .ZN(n871) );
  XNOR2_X1 U966 ( .A(n871), .B(KEYINPUT50), .ZN(n879) );
  XOR2_X1 U967 ( .A(G160), .B(G2084), .Z(n872) );
  NOR2_X1 U968 ( .A1(n873), .A2(n872), .ZN(n876) );
  NOR2_X1 U969 ( .A1(n874), .A2(n977), .ZN(n875) );
  NAND2_X1 U970 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U971 ( .A(KEYINPUT115), .B(n877), .ZN(n878) );
  NAND2_X1 U972 ( .A1(n879), .A2(n878), .ZN(n880) );
  NOR2_X1 U973 ( .A1(n881), .A2(n880), .ZN(n882) );
  NAND2_X1 U974 ( .A1(n883), .A2(n882), .ZN(n884) );
  XNOR2_X1 U975 ( .A(n884), .B(KEYINPUT119), .ZN(n885) );
  XOR2_X1 U976 ( .A(KEYINPUT52), .B(n885), .Z(n886) );
  NAND2_X1 U977 ( .A1(G29), .A2(n886), .ZN(n887) );
  NAND2_X1 U978 ( .A1(n888), .A2(n887), .ZN(n941) );
  XNOR2_X1 U979 ( .A(G16), .B(KEYINPUT56), .ZN(n913) );
  XNOR2_X1 U980 ( .A(n1009), .B(G1348), .ZN(n911) );
  XOR2_X1 U981 ( .A(G1966), .B(G168), .Z(n889) );
  XNOR2_X1 U982 ( .A(KEYINPUT123), .B(n889), .ZN(n891) );
  NAND2_X1 U983 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U984 ( .A(n892), .B(KEYINPUT57), .ZN(n906) );
  INV_X1 U985 ( .A(G1971), .ZN(n893) );
  NOR2_X1 U986 ( .A1(G166), .A2(n893), .ZN(n897) );
  NAND2_X1 U987 ( .A1(n895), .A2(n894), .ZN(n896) );
  NOR2_X1 U988 ( .A1(n897), .A2(n896), .ZN(n901) );
  XNOR2_X1 U989 ( .A(G1956), .B(G299), .ZN(n898) );
  NOR2_X1 U990 ( .A1(n899), .A2(n898), .ZN(n900) );
  NAND2_X1 U991 ( .A1(n901), .A2(n900), .ZN(n904) );
  XOR2_X1 U992 ( .A(G1961), .B(G171), .Z(n902) );
  XNOR2_X1 U993 ( .A(KEYINPUT124), .B(n902), .ZN(n903) );
  NOR2_X1 U994 ( .A1(n904), .A2(n903), .ZN(n905) );
  NAND2_X1 U995 ( .A1(n906), .A2(n905), .ZN(n909) );
  XNOR2_X1 U996 ( .A(G1341), .B(n907), .ZN(n908) );
  NOR2_X1 U997 ( .A1(n909), .A2(n908), .ZN(n910) );
  NAND2_X1 U998 ( .A1(n911), .A2(n910), .ZN(n912) );
  NAND2_X1 U999 ( .A1(n913), .A2(n912), .ZN(n938) );
  INV_X1 U1000 ( .A(G16), .ZN(n936) );
  XNOR2_X1 U1001 ( .A(G1348), .B(KEYINPUT59), .ZN(n914) );
  XNOR2_X1 U1002 ( .A(n914), .B(G4), .ZN(n918) );
  XNOR2_X1 U1003 ( .A(G1981), .B(G6), .ZN(n916) );
  XNOR2_X1 U1004 ( .A(G1956), .B(G20), .ZN(n915) );
  NOR2_X1 U1005 ( .A1(n916), .A2(n915), .ZN(n917) );
  NAND2_X1 U1006 ( .A1(n918), .A2(n917), .ZN(n921) );
  XOR2_X1 U1007 ( .A(KEYINPUT125), .B(G1341), .Z(n919) );
  XNOR2_X1 U1008 ( .A(G19), .B(n919), .ZN(n920) );
  NOR2_X1 U1009 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1010 ( .A(KEYINPUT60), .B(n922), .ZN(n926) );
  XNOR2_X1 U1011 ( .A(G1966), .B(G21), .ZN(n924) );
  XNOR2_X1 U1012 ( .A(G5), .B(G1961), .ZN(n923) );
  NOR2_X1 U1013 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1014 ( .A1(n926), .A2(n925), .ZN(n933) );
  XNOR2_X1 U1015 ( .A(G1976), .B(G23), .ZN(n928) );
  XNOR2_X1 U1016 ( .A(G1971), .B(G22), .ZN(n927) );
  NOR2_X1 U1017 ( .A1(n928), .A2(n927), .ZN(n930) );
  XOR2_X1 U1018 ( .A(G1986), .B(G24), .Z(n929) );
  NAND2_X1 U1019 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1020 ( .A(KEYINPUT58), .B(n931), .ZN(n932) );
  NOR2_X1 U1021 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1022 ( .A(KEYINPUT61), .B(n934), .ZN(n935) );
  NAND2_X1 U1023 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1024 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1025 ( .A(n939), .B(KEYINPUT126), .ZN(n940) );
  NOR2_X1 U1026 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1027 ( .A1(n942), .A2(G11), .ZN(n943) );
  XOR2_X1 U1028 ( .A(KEYINPUT62), .B(n943), .Z(G311) );
  XNOR2_X1 U1029 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1030 ( .A(G120), .ZN(G236) );
  INV_X1 U1031 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1032 ( .A1(n945), .A2(n944), .ZN(G325) );
  INV_X1 U1033 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U1034 ( .A(G1348), .B(G2454), .ZN(n946) );
  XNOR2_X1 U1035 ( .A(n946), .B(G2430), .ZN(n947) );
  XNOR2_X1 U1036 ( .A(n947), .B(G1341), .ZN(n953) );
  XOR2_X1 U1037 ( .A(G2443), .B(G2427), .Z(n949) );
  XNOR2_X1 U1038 ( .A(G2438), .B(G2446), .ZN(n948) );
  XNOR2_X1 U1039 ( .A(n949), .B(n948), .ZN(n951) );
  XOR2_X1 U1040 ( .A(G2451), .B(G2435), .Z(n950) );
  XNOR2_X1 U1041 ( .A(n951), .B(n950), .ZN(n952) );
  XNOR2_X1 U1042 ( .A(n953), .B(n952), .ZN(n954) );
  NAND2_X1 U1043 ( .A1(n954), .A2(G14), .ZN(n955) );
  XOR2_X1 U1044 ( .A(KEYINPUT98), .B(n955), .Z(G401) );
  INV_X1 U1045 ( .A(n956), .ZN(G319) );
  XOR2_X1 U1046 ( .A(KEYINPUT42), .B(G2078), .Z(n958) );
  XNOR2_X1 U1047 ( .A(G2067), .B(G2084), .ZN(n957) );
  XNOR2_X1 U1048 ( .A(n958), .B(n957), .ZN(n959) );
  XOR2_X1 U1049 ( .A(n959), .B(G2678), .Z(n961) );
  XNOR2_X1 U1050 ( .A(G2072), .B(KEYINPUT101), .ZN(n960) );
  XNOR2_X1 U1051 ( .A(n961), .B(n960), .ZN(n965) );
  XOR2_X1 U1052 ( .A(G2100), .B(G2096), .Z(n963) );
  XNOR2_X1 U1053 ( .A(G2090), .B(KEYINPUT43), .ZN(n962) );
  XNOR2_X1 U1054 ( .A(n963), .B(n962), .ZN(n964) );
  XOR2_X1 U1055 ( .A(n965), .B(n964), .Z(G227) );
  XOR2_X1 U1056 ( .A(KEYINPUT102), .B(G2474), .Z(n967) );
  XNOR2_X1 U1057 ( .A(G1981), .B(G1976), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(n967), .B(n966), .ZN(n968) );
  XOR2_X1 U1059 ( .A(n968), .B(KEYINPUT103), .Z(n970) );
  XNOR2_X1 U1060 ( .A(G1956), .B(KEYINPUT41), .ZN(n969) );
  XNOR2_X1 U1061 ( .A(n970), .B(n969), .ZN(n974) );
  XOR2_X1 U1062 ( .A(G1961), .B(G1966), .Z(n972) );
  XNOR2_X1 U1063 ( .A(G1986), .B(G1971), .ZN(n971) );
  XNOR2_X1 U1064 ( .A(n972), .B(n971), .ZN(n973) );
  XOR2_X1 U1065 ( .A(n974), .B(n973), .Z(n976) );
  XNOR2_X1 U1066 ( .A(G1996), .B(G1991), .ZN(n975) );
  XNOR2_X1 U1067 ( .A(n976), .B(n975), .ZN(G229) );
  XOR2_X1 U1068 ( .A(n977), .B(G162), .Z(n978) );
  XNOR2_X1 U1069 ( .A(n979), .B(n978), .ZN(n983) );
  XOR2_X1 U1070 ( .A(KEYINPUT105), .B(KEYINPUT46), .Z(n981) );
  XNOR2_X1 U1071 ( .A(KEYINPUT48), .B(KEYINPUT109), .ZN(n980) );
  XNOR2_X1 U1072 ( .A(n981), .B(n980), .ZN(n982) );
  XOR2_X1 U1073 ( .A(n983), .B(n982), .Z(n999) );
  NAND2_X1 U1074 ( .A1(G118), .A2(n984), .ZN(n987) );
  NAND2_X1 U1075 ( .A1(G130), .A2(n985), .ZN(n986) );
  NAND2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n993) );
  NAND2_X1 U1077 ( .A1(n988), .A2(G106), .ZN(n990) );
  NAND2_X1 U1078 ( .A1(G142), .A2(n698), .ZN(n989) );
  NAND2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1080 ( .A(n991), .B(KEYINPUT45), .Z(n992) );
  NOR2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n995) );
  XNOR2_X1 U1082 ( .A(n995), .B(n994), .ZN(n996) );
  XOR2_X1 U1083 ( .A(G160), .B(n996), .Z(n997) );
  XNOR2_X1 U1084 ( .A(G164), .B(n997), .ZN(n998) );
  XNOR2_X1 U1085 ( .A(n999), .B(n998), .ZN(n1000) );
  XOR2_X1 U1086 ( .A(n1001), .B(n1000), .Z(n1002) );
  XNOR2_X1 U1087 ( .A(n1003), .B(n1002), .ZN(n1004) );
  NOR2_X1 U1088 ( .A1(G37), .A2(n1004), .ZN(G395) );
  XOR2_X1 U1089 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n1006) );
  XNOR2_X1 U1090 ( .A(G171), .B(KEYINPUT110), .ZN(n1005) );
  XNOR2_X1 U1091 ( .A(n1006), .B(n1005), .ZN(n1008) );
  XNOR2_X1 U1092 ( .A(n1008), .B(n1007), .ZN(n1011) );
  XOR2_X1 U1093 ( .A(G286), .B(n1009), .Z(n1010) );
  XNOR2_X1 U1094 ( .A(n1011), .B(n1010), .ZN(n1012) );
  NOR2_X1 U1095 ( .A1(G37), .A2(n1012), .ZN(G397) );
  NOR2_X1 U1096 ( .A1(G227), .A2(G229), .ZN(n1013) );
  XOR2_X1 U1097 ( .A(KEYINPUT49), .B(n1013), .Z(n1014) );
  NAND2_X1 U1098 ( .A1(G319), .A2(n1014), .ZN(n1015) );
  NOR2_X1 U1099 ( .A1(G401), .A2(n1015), .ZN(n1018) );
  NOR2_X1 U1100 ( .A1(G395), .A2(G397), .ZN(n1016) );
  XOR2_X1 U1101 ( .A(KEYINPUT113), .B(n1016), .Z(n1017) );
  NAND2_X1 U1102 ( .A1(n1018), .A2(n1017), .ZN(G225) );
  INV_X1 U1103 ( .A(G225), .ZN(G308) );
  INV_X1 U1104 ( .A(G69), .ZN(G235) );
endmodule

