//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 1 1 1 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 1 1 1 1 1 0 1 0 1 0 0 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953;
  INV_X1    g000(.A(G143), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT1), .B1(new_n187), .B2(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT69), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT69), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(KEYINPUT1), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n189), .A2(G128), .A3(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(G143), .B(G146), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n187), .A2(G146), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT1), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n191), .A2(new_n198), .A3(new_n199), .A4(G128), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT68), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT68), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n195), .A2(new_n202), .A3(new_n199), .A4(G128), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n197), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n206));
  INV_X1    g020(.A(G134), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G137), .ZN(new_n209));
  NAND2_X1  g023(.A1(KEYINPUT64), .A2(G134), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n211), .B(KEYINPUT66), .C1(G134), .C2(new_n209), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n208), .A2(new_n213), .A3(new_n209), .A4(new_n210), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n212), .A2(KEYINPUT67), .A3(G131), .A4(new_n214), .ZN(new_n215));
  AND2_X1   g029(.A1(KEYINPUT64), .A2(G134), .ZN(new_n216));
  NOR2_X1   g030(.A1(KEYINPUT64), .A2(G134), .ZN(new_n217));
  NOR3_X1   g031(.A1(new_n216), .A2(new_n217), .A3(G137), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT66), .B1(new_n209), .B2(G134), .ZN(new_n219));
  OAI211_X1 g033(.A(G131), .B(new_n214), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n215), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT11), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n218), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g039(.A1(G134), .A2(G137), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n216), .A2(new_n217), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n226), .B1(new_n227), .B2(G137), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n225), .B1(new_n228), .B2(new_n224), .ZN(new_n229));
  INV_X1    g043(.A(G131), .ZN(new_n230));
  AOI21_X1  g044(.A(KEYINPUT65), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n208), .A2(G137), .A3(new_n210), .ZN(new_n232));
  INV_X1    g046(.A(new_n226), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n224), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n211), .A2(KEYINPUT11), .ZN(new_n235));
  OAI211_X1 g049(.A(KEYINPUT65), .B(new_n230), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n205), .B(new_n223), .C1(new_n231), .C2(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n230), .B1(new_n234), .B2(new_n235), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT65), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n234), .A2(new_n235), .ZN(new_n242));
  AOI22_X1  g056(.A1(new_n241), .A2(new_n236), .B1(G131), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(KEYINPUT0), .A2(G128), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n195), .A2(new_n244), .ZN(new_n245));
  XOR2_X1   g059(.A(KEYINPUT0), .B(G128), .Z(new_n246));
  OAI21_X1  g060(.A(new_n245), .B1(new_n246), .B2(new_n195), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n238), .B1(new_n243), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT30), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(G116), .B(G119), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(KEYINPUT70), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT2), .B(G113), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n253), .B(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n242), .A2(G131), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n256), .B1(new_n231), .B2(new_n237), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n247), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT30), .A3(new_n238), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n251), .A2(new_n255), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n255), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n238), .B(new_n261), .C1(new_n243), .C2(new_n248), .ZN(new_n262));
  OR2_X1    g076(.A1(KEYINPUT71), .A2(G953), .ZN(new_n263));
  NAND2_X1  g077(.A1(KEYINPUT71), .A2(G953), .ZN(new_n264));
  AOI21_X1  g078(.A(G237), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G210), .ZN(new_n266));
  XOR2_X1   g080(.A(KEYINPUT26), .B(G101), .Z(new_n267));
  XNOR2_X1  g081(.A(new_n266), .B(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT72), .B(KEYINPUT27), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n268), .B(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n260), .A2(new_n262), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT31), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT28), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n249), .A2(new_n255), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n274), .B1(new_n275), .B2(new_n262), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n262), .A2(new_n274), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n270), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT31), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n260), .A2(new_n280), .A3(new_n262), .A4(new_n271), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n273), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(G472), .A2(G902), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT32), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G902), .ZN(new_n287));
  INV_X1    g101(.A(new_n262), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n261), .B1(new_n258), .B2(new_n238), .ZN(new_n289));
  OAI21_X1  g103(.A(KEYINPUT28), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n290), .A2(KEYINPUT29), .A3(new_n277), .A4(new_n271), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(new_n277), .A3(new_n271), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT29), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n271), .B1(new_n260), .B2(new_n262), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n287), .B(new_n291), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G472), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n282), .A2(KEYINPUT32), .A3(new_n283), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n286), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G217), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n300), .B1(G234), .B2(new_n287), .ZN(new_n301));
  XNOR2_X1  g115(.A(G125), .B(G140), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT16), .ZN(new_n303));
  INV_X1    g117(.A(G140), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G125), .ZN(new_n305));
  OR2_X1    g119(.A1(new_n305), .A2(KEYINPUT16), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n303), .A2(G146), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G119), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G128), .ZN(new_n309));
  INV_X1    g123(.A(G128), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G119), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(KEYINPUT73), .ZN(new_n313));
  XOR2_X1   g127(.A(KEYINPUT24), .B(G110), .Z(new_n314));
  NAND2_X1  g128(.A1(new_n311), .A2(KEYINPUT75), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT23), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT23), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n311), .A2(KEYINPUT75), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n316), .A2(new_n309), .A3(new_n318), .ZN(new_n319));
  OAI22_X1  g133(.A1(new_n313), .A2(new_n314), .B1(new_n319), .B2(G110), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT76), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n307), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT77), .ZN(new_n323));
  INV_X1    g137(.A(G125), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G140), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n323), .B1(new_n305), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n302), .A2(new_n323), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(new_n328), .A3(new_n190), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n322), .B(new_n329), .C1(new_n321), .C2(new_n320), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n313), .A2(new_n314), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT74), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n331), .B(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(G146), .B1(new_n303), .B2(new_n306), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n307), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n335), .B1(G110), .B2(new_n319), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n330), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n263), .A2(new_n264), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(G221), .A3(G234), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n340), .B(KEYINPUT22), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(new_n209), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n338), .B(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT25), .B1(new_n344), .B2(new_n287), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT25), .ZN(new_n346));
  NOR3_X1   g160(.A1(new_n343), .A2(new_n346), .A3(G902), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n301), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n301), .A2(G902), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G475), .ZN(new_n352));
  AOI21_X1  g166(.A(G143), .B1(new_n265), .B2(G214), .ZN(new_n353));
  INV_X1    g167(.A(G237), .ZN(new_n354));
  AND2_X1   g168(.A1(KEYINPUT71), .A2(G953), .ZN(new_n355));
  NOR2_X1   g169(.A1(KEYINPUT71), .A2(G953), .ZN(new_n356));
  OAI211_X1 g170(.A(G214), .B(new_n354), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n357), .A2(new_n187), .ZN(new_n358));
  OAI21_X1  g172(.A(G131), .B1(new_n353), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT17), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n265), .A2(G143), .A3(G214), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n357), .A2(new_n187), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n230), .A3(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n359), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n361), .A2(new_n362), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(KEYINPUT17), .A3(G131), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n364), .A2(new_n335), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n365), .A2(KEYINPUT18), .A3(G131), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n329), .B1(new_n190), .B2(new_n302), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT18), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n361), .B(new_n362), .C1(new_n370), .C2(new_n230), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n368), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  XNOR2_X1  g186(.A(G113), .B(G122), .ZN(new_n373));
  INV_X1    g187(.A(G104), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n373), .B(new_n374), .ZN(new_n375));
  XOR2_X1   g189(.A(new_n375), .B(KEYINPUT84), .Z(new_n376));
  AND3_X1   g190(.A1(new_n367), .A2(new_n372), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT19), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n378), .B1(new_n326), .B2(KEYINPUT82), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT77), .B1(new_n378), .B2(KEYINPUT82), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n302), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(G146), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT83), .B1(new_n382), .B2(new_n307), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n359), .A2(new_n363), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT83), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n303), .A2(G146), .A3(new_n306), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT82), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n387), .B1(new_n302), .B2(new_n323), .ZN(new_n388));
  AOI22_X1  g202(.A1(new_n388), .A2(new_n378), .B1(new_n302), .B2(new_n380), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n385), .B(new_n386), .C1(new_n389), .C2(G146), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n383), .A2(new_n384), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n375), .B1(new_n391), .B2(new_n372), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n352), .B(new_n287), .C1(new_n377), .C2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT20), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n367), .A2(new_n372), .A3(new_n376), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n368), .A2(new_n369), .A3(new_n371), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n379), .A2(new_n381), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n307), .B1(new_n398), .B2(new_n190), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n399), .A2(new_n385), .B1(new_n359), .B2(new_n363), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n397), .B1(new_n400), .B2(new_n383), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n396), .B1(new_n401), .B2(new_n375), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n402), .A2(KEYINPUT20), .A3(new_n352), .A4(new_n287), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n375), .B1(new_n367), .B2(new_n372), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n287), .B1(new_n377), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G475), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n395), .A2(new_n403), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT85), .ZN(new_n408));
  INV_X1    g222(.A(G478), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n409), .A2(KEYINPUT15), .ZN(new_n410));
  INV_X1    g224(.A(G122), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G116), .ZN(new_n412));
  INV_X1    g226(.A(G116), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G122), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(KEYINPUT78), .B(G107), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n415), .B(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n310), .A2(G143), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n187), .A2(G128), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OR2_X1    g234(.A1(new_n420), .A2(new_n227), .ZN(new_n421));
  AOI21_X1  g235(.A(KEYINPUT13), .B1(new_n187), .B2(G128), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n187), .A2(G128), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT86), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT86), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n310), .A2(G143), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n425), .B(new_n418), .C1(new_n426), .C2(KEYINPUT13), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(KEYINPUT13), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n424), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n417), .B(new_n421), .C1(new_n429), .C2(new_n207), .ZN(new_n430));
  XNOR2_X1  g244(.A(KEYINPUT9), .B(G234), .ZN(new_n431));
  NOR3_X1   g245(.A1(new_n431), .A2(new_n300), .A3(G953), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n420), .B(new_n227), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n415), .A2(new_n416), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT87), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n414), .A2(KEYINPUT14), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n412), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n414), .A2(KEYINPUT14), .ZN(new_n439));
  OAI21_X1  g253(.A(G107), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n415), .A2(KEYINPUT87), .A3(new_n416), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n433), .A2(new_n436), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n430), .A2(new_n432), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT88), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n430), .A2(new_n442), .ZN(new_n445));
  INV_X1    g259(.A(new_n432), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT88), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n430), .A2(new_n448), .A3(new_n432), .A4(new_n442), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n444), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n287), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT89), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n410), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n452), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n450), .A2(KEYINPUT89), .A3(new_n287), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n453), .B1(new_n456), .B2(new_n410), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT85), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n395), .A2(new_n403), .A3(new_n458), .A4(new_n406), .ZN(new_n459));
  INV_X1    g273(.A(G952), .ZN(new_n460));
  AOI211_X1 g274(.A(G953), .B(new_n460), .C1(G234), .C2(G237), .ZN(new_n461));
  AOI211_X1 g275(.A(new_n287), .B(new_n339), .C1(G234), .C2(G237), .ZN(new_n462));
  XOR2_X1   g276(.A(KEYINPUT21), .B(G898), .Z(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n461), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n408), .A2(new_n457), .A3(new_n459), .A4(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G469), .ZN(new_n468));
  OR2_X1    g282(.A1(new_n374), .A2(G107), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n469), .B1(new_n416), .B2(G104), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(G101), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT3), .ZN(new_n472));
  AND2_X1   g286(.A1(KEYINPUT78), .A2(G107), .ZN(new_n473));
  NOR2_X1   g287(.A1(KEYINPUT78), .A2(G107), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n472), .B(G104), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G101), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n374), .A2(G107), .ZN(new_n477));
  OAI21_X1  g291(.A(KEYINPUT3), .B1(new_n374), .B2(G107), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n475), .A2(new_n476), .A3(new_n477), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n471), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n188), .A2(G128), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n201), .A2(new_n203), .B1(new_n196), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  OR2_X1    g297(.A1(new_n483), .A2(KEYINPUT10), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n475), .A2(new_n477), .A3(new_n478), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(G101), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(KEYINPUT4), .A3(new_n479), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT4), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n485), .A2(new_n488), .A3(G101), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n487), .A2(new_n247), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n480), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(KEYINPUT10), .A3(new_n205), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n484), .A2(new_n243), .A3(new_n490), .A4(new_n492), .ZN(new_n493));
  AOI22_X1  g307(.A1(new_n196), .A2(new_n194), .B1(new_n201), .B2(new_n203), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n483), .B1(new_n494), .B2(new_n480), .ZN(new_n495));
  OAI21_X1  g309(.A(KEYINPUT12), .B1(new_n495), .B2(new_n243), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT12), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n491), .A2(new_n205), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n257), .B(new_n497), .C1(new_n483), .C2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n339), .A2(G227), .ZN(new_n500));
  XNOR2_X1  g314(.A(G110), .B(G140), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n500), .B(new_n501), .ZN(new_n502));
  AND4_X1   g316(.A1(new_n493), .A2(new_n496), .A3(new_n499), .A4(new_n502), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n492), .B(new_n490), .C1(KEYINPUT10), .C2(new_n483), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n257), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n502), .B1(new_n505), .B2(new_n493), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n468), .B(new_n287), .C1(new_n503), .C2(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n468), .A2(new_n287), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n496), .A2(new_n493), .A3(new_n499), .ZN(new_n510));
  INV_X1    g324(.A(new_n502), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n505), .A2(new_n493), .A3(new_n502), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(G469), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n507), .A2(new_n509), .A3(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(G221), .B1(new_n431), .B2(G902), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n487), .A2(new_n255), .A3(new_n489), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n252), .A2(KEYINPUT5), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n413), .A2(KEYINPUT5), .A3(G119), .ZN(new_n520));
  INV_X1    g334(.A(G113), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n254), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n519), .A2(new_n522), .B1(new_n523), .B2(new_n252), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n491), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n518), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(G110), .B(G122), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(KEYINPUT79), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n518), .A2(new_n525), .A3(new_n528), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(KEYINPUT6), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(G224), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(G953), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n494), .A2(G125), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n247), .A2(G125), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n535), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n534), .B(new_n537), .C1(new_n494), .C2(G125), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT6), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n526), .A2(new_n542), .A3(new_n529), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n532), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT80), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n519), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n252), .A2(KEYINPUT80), .A3(KEYINPUT5), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n522), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n523), .A2(new_n252), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n491), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT8), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n480), .A2(new_n524), .B1(new_n552), .B2(new_n528), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n529), .A2(KEYINPUT8), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n551), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT7), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n556), .B(new_n537), .C1(new_n494), .C2(G125), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g372(.A(KEYINPUT7), .B(new_n535), .C1(new_n536), .C2(new_n538), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n558), .A2(new_n531), .A3(new_n559), .A4(new_n540), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n544), .A2(new_n287), .A3(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(G210), .B1(G237), .B2(G902), .ZN(new_n562));
  XOR2_X1   g376(.A(new_n562), .B(KEYINPUT81), .Z(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(G214), .B1(G237), .B2(G902), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n544), .A2(new_n560), .A3(new_n287), .A4(new_n563), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n467), .A2(new_n517), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n299), .A2(new_n351), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(G101), .ZN(G3));
  NAND2_X1  g385(.A1(new_n282), .A2(new_n287), .ZN(new_n572));
  AOI22_X1  g386(.A1(new_n572), .A2(G472), .B1(new_n282), .B2(new_n283), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n348), .A2(new_n350), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n574), .A2(new_n575), .A3(new_n517), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n408), .A2(new_n459), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT33), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n450), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n445), .A2(KEYINPUT90), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(new_n446), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n579), .B1(KEYINPUT33), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n409), .A2(G902), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n451), .A2(new_n409), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n577), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n565), .A2(new_n566), .A3(new_n567), .A4(new_n466), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n576), .A2(new_n589), .ZN(new_n590));
  XOR2_X1   g404(.A(KEYINPUT34), .B(G104), .Z(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(G6));
  INV_X1    g406(.A(new_n457), .ZN(new_n593));
  INV_X1    g407(.A(new_n407), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(new_n588), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n576), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g411(.A(KEYINPUT35), .B(G107), .Z(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(G9));
  NOR2_X1   g413(.A1(new_n342), .A2(KEYINPUT36), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n338), .B(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n349), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n348), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n569), .A2(new_n573), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(KEYINPUT91), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(KEYINPUT37), .ZN(new_n606));
  XOR2_X1   g420(.A(new_n606), .B(G110), .Z(G12));
  INV_X1    g421(.A(new_n517), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n299), .A2(new_n608), .A3(new_n603), .ZN(new_n609));
  INV_X1    g423(.A(new_n568), .ZN(new_n610));
  INV_X1    g424(.A(G900), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n461), .B1(new_n462), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n595), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n609), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(G128), .ZN(G30));
  AND3_X1   g429(.A1(new_n282), .A2(KEYINPUT32), .A3(new_n283), .ZN(new_n616));
  AOI21_X1  g430(.A(KEYINPUT32), .B1(new_n282), .B2(new_n283), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n270), .B1(new_n288), .B2(new_n289), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n272), .A2(G472), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(G472), .A2(G902), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT92), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n620), .A2(KEYINPUT92), .A3(new_n621), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(KEYINPUT93), .B1(new_n618), .B2(new_n626), .ZN(new_n627));
  AND4_X1   g441(.A1(KEYINPUT93), .A2(new_n286), .A3(new_n626), .A4(new_n298), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(new_n612), .B(KEYINPUT39), .Z(new_n631));
  NAND2_X1  g445(.A1(new_n608), .A2(new_n631), .ZN(new_n632));
  OR2_X1    g446(.A1(new_n632), .A2(KEYINPUT40), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(KEYINPUT40), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n577), .A2(new_n593), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n565), .A2(new_n567), .ZN(new_n637));
  XOR2_X1   g451(.A(new_n637), .B(KEYINPUT38), .Z(new_n638));
  NAND4_X1  g452(.A1(new_n633), .A2(new_n634), .A3(new_n636), .A4(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n603), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n630), .A2(new_n640), .A3(new_n566), .A4(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G143), .ZN(G45));
  AOI22_X1  g457(.A1(new_n408), .A2(new_n459), .B1(new_n584), .B2(new_n585), .ZN(new_n644));
  INV_X1    g458(.A(new_n612), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OR3_X1    g460(.A1(new_n646), .A2(KEYINPUT94), .A3(new_n568), .ZN(new_n647));
  OAI21_X1  g461(.A(KEYINPUT94), .B1(new_n646), .B2(new_n568), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n609), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G146), .ZN(G48));
  AOI21_X1  g464(.A(new_n575), .B1(new_n618), .B2(new_n297), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n503), .A2(new_n506), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n468), .B1(new_n652), .B2(new_n287), .ZN(new_n653));
  INV_X1    g467(.A(new_n516), .ZN(new_n654));
  INV_X1    g468(.A(new_n507), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n651), .A2(new_n589), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT41), .B(G113), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G15));
  NAND3_X1  g473(.A1(new_n651), .A2(new_n596), .A3(new_n656), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G116), .ZN(G18));
  INV_X1    g475(.A(new_n656), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(new_n568), .ZN(new_n663));
  INV_X1    g477(.A(new_n467), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n663), .A2(new_n299), .A3(new_n664), .A4(new_n603), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G119), .ZN(G21));
  NOR2_X1   g480(.A1(new_n662), .A2(new_n465), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT95), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n668), .B1(new_n276), .B2(new_n278), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n290), .A2(KEYINPUT95), .A3(new_n277), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n669), .A2(new_n670), .A3(new_n270), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n671), .A2(new_n273), .A3(new_n281), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n283), .ZN(new_n673));
  AOI21_X1  g487(.A(KEYINPUT96), .B1(new_n572), .B2(G472), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT96), .ZN(new_n675));
  INV_X1    g489(.A(G472), .ZN(new_n676));
  AOI211_X1 g490(.A(new_n675), .B(new_n676), .C1(new_n282), .C2(new_n287), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n351), .B(new_n673), .C1(new_n674), .C2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT97), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n635), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n577), .A2(KEYINPUT97), .A3(new_n593), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n681), .A2(new_n610), .A3(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT98), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AOI211_X1 g499(.A(new_n680), .B(new_n457), .C1(new_n408), .C2(new_n459), .ZN(new_n686));
  AOI21_X1  g500(.A(KEYINPUT97), .B1(new_n577), .B2(new_n593), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(KEYINPUT98), .B1(new_n688), .B2(new_n610), .ZN(new_n689));
  OAI211_X1 g503(.A(new_n667), .B(new_n679), .C1(new_n685), .C2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(KEYINPUT99), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n683), .B(new_n684), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT99), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n692), .A2(new_n693), .A3(new_n667), .A4(new_n679), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G122), .ZN(G24));
  OAI211_X1 g510(.A(new_n603), .B(new_n673), .C1(new_n674), .C2(new_n677), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n646), .A2(KEYINPUT100), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT100), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n644), .A2(new_n700), .A3(new_n645), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n698), .A2(new_n663), .A3(new_n702), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT101), .B(G125), .Z(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G27));
  NAND2_X1  g519(.A1(new_n637), .A2(new_n566), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT103), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n507), .A2(new_n509), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT102), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n513), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n513), .A2(new_n710), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n711), .A2(G469), .A3(new_n512), .A4(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n654), .B1(new_n709), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n637), .A2(KEYINPUT103), .A3(new_n566), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n708), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(KEYINPUT104), .ZN(new_n717));
  AOI21_X1  g531(.A(KEYINPUT103), .B1(new_n637), .B2(new_n566), .ZN(new_n718));
  INV_X1    g532(.A(new_n566), .ZN(new_n719));
  AOI211_X1 g533(.A(new_n707), .B(new_n719), .C1(new_n565), .C2(new_n567), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT104), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n722), .A3(new_n714), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n717), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n724), .A2(new_n651), .A3(new_n702), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT42), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n726), .B1(new_n717), .B2(new_n723), .ZN(new_n728));
  OAI21_X1  g542(.A(KEYINPUT105), .B1(new_n616), .B2(new_n617), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT105), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n286), .A2(new_n730), .A3(new_n298), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n729), .A2(new_n731), .A3(new_n297), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n728), .A2(new_n351), .A3(new_n702), .A4(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n727), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G131), .ZN(G33));
  NOR2_X1   g549(.A1(new_n716), .A2(KEYINPUT104), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n722), .B1(new_n721), .B2(new_n714), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n651), .B(new_n613), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT106), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT106), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n724), .A2(new_n740), .A3(new_n651), .A4(new_n613), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G134), .ZN(G36));
  NAND4_X1  g557(.A1(new_n711), .A2(KEYINPUT45), .A3(new_n512), .A4(new_n712), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n744), .A2(KEYINPUT107), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(KEYINPUT107), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n468), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n512), .A2(new_n513), .ZN(new_n748));
  OR2_X1    g562(.A1(new_n748), .A2(KEYINPUT45), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n750), .A2(KEYINPUT46), .A3(new_n509), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT108), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n751), .A2(new_n752), .A3(new_n507), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n752), .B1(new_n751), .B2(new_n507), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT46), .B1(new_n750), .B2(new_n509), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(new_n654), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n586), .A2(new_n408), .A3(new_n459), .ZN(new_n758));
  XOR2_X1   g572(.A(new_n758), .B(KEYINPUT43), .Z(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(new_n574), .A3(new_n603), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT44), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n757), .A2(new_n631), .A3(new_n721), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(KEYINPUT109), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G137), .ZN(G39));
  INV_X1    g578(.A(KEYINPUT110), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n765), .A2(KEYINPUT47), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n765), .A2(KEYINPUT47), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n757), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI22_X1  g582(.A1(new_n756), .A2(new_n654), .B1(new_n765), .B2(KEYINPUT47), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n299), .A2(new_n351), .ZN(new_n770));
  INV_X1    g584(.A(new_n721), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(new_n646), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n768), .A2(new_n769), .A3(new_n770), .A4(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G140), .ZN(G42));
  INV_X1    g588(.A(new_n638), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n775), .A2(new_n351), .A3(new_n566), .A4(new_n516), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n653), .A2(new_n655), .ZN(new_n777));
  XOR2_X1   g591(.A(new_n777), .B(KEYINPUT49), .Z(new_n778));
  OR4_X1    g592(.A1(new_n630), .A2(new_n758), .A3(new_n776), .A4(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT112), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n593), .A2(new_n612), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n609), .A2(new_n594), .A3(new_n721), .A4(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n593), .A2(new_n408), .A3(new_n459), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n588), .B1(new_n587), .B2(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n784), .A2(new_n351), .A3(new_n608), .A4(new_n573), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n785), .A2(new_n570), .A3(new_n604), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n698), .A2(new_n724), .A3(new_n702), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n782), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n788), .A2(new_n734), .A3(new_n742), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n657), .A2(new_n660), .A3(new_n665), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n790), .B1(new_n691), .B2(new_n694), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n641), .B1(new_n685), .B2(new_n689), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n645), .B(new_n714), .C1(new_n627), .C2(new_n628), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n649), .A2(new_n703), .A3(new_n614), .ZN(new_n795));
  OAI21_X1  g609(.A(KEYINPUT52), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n714), .ZN(new_n797));
  INV_X1    g611(.A(new_n628), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n618), .A2(new_n626), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT93), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n797), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n802), .A2(new_n692), .A3(new_n641), .A4(new_n645), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n703), .A2(new_n614), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n803), .A2(new_n804), .A3(new_n805), .A4(new_n649), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n789), .A2(new_n791), .A3(new_n796), .A4(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n780), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n807), .A2(new_n808), .ZN(new_n810));
  AOI22_X1  g624(.A1(new_n727), .A2(new_n733), .B1(new_n739), .B2(new_n741), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n791), .A2(new_n811), .A3(new_n788), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n806), .A2(new_n796), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n812), .A2(new_n813), .A3(KEYINPUT112), .A4(KEYINPUT53), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n809), .A2(new_n810), .A3(new_n814), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n815), .A2(KEYINPUT54), .ZN(new_n816));
  INV_X1    g630(.A(new_n807), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT53), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(KEYINPUT111), .A3(new_n810), .ZN(new_n819));
  OR3_X1    g633(.A1(new_n807), .A2(KEYINPUT111), .A3(new_n808), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n819), .A2(KEYINPUT54), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n816), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n768), .A2(new_n769), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n777), .B(KEYINPUT113), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n654), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n759), .A2(new_n461), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(new_n678), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n827), .A2(new_n721), .A3(new_n829), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n828), .A2(new_n662), .A3(new_n771), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n698), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n771), .A2(new_n662), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n629), .A2(new_n351), .A3(new_n461), .A4(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT114), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n577), .A2(new_n586), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n829), .A2(new_n719), .A3(new_n775), .A4(new_n656), .ZN(new_n838));
  XOR2_X1   g652(.A(new_n838), .B(KEYINPUT50), .Z(new_n839));
  NAND4_X1  g653(.A1(new_n830), .A2(new_n832), .A3(new_n837), .A4(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT51), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n831), .A2(new_n351), .A3(new_n732), .ZN(new_n843));
  XOR2_X1   g657(.A(KEYINPUT116), .B(KEYINPUT48), .Z(new_n844));
  XNOR2_X1  g658(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n460), .A2(G953), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n835), .A2(new_n644), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n848), .B1(new_n840), .B2(new_n841), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n829), .A2(new_n663), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT115), .ZN(new_n851));
  AND4_X1   g665(.A1(new_n823), .A2(new_n842), .A3(new_n849), .A4(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(G952), .A2(G953), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(KEYINPUT117), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n779), .B1(new_n852), .B2(new_n854), .ZN(G75));
  NOR2_X1   g669(.A1(new_n339), .A2(G952), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n815), .A2(G902), .A3(new_n563), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT56), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n532), .A2(new_n543), .ZN(new_n861));
  XOR2_X1   g675(.A(new_n861), .B(KEYINPUT118), .Z(new_n862));
  XOR2_X1   g676(.A(new_n862), .B(new_n541), .Z(new_n863));
  XOR2_X1   g677(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n864));
  XNOR2_X1  g678(.A(new_n863), .B(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n860), .A2(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n858), .A2(new_n857), .A3(new_n859), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n868), .A2(new_n860), .ZN(new_n869));
  AOI211_X1 g683(.A(new_n856), .B(new_n867), .C1(new_n869), .C2(new_n866), .ZN(G51));
  NAND2_X1  g684(.A1(new_n815), .A2(KEYINPUT54), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n816), .A2(KEYINPUT121), .A3(new_n871), .ZN(new_n872));
  OR3_X1    g686(.A1(new_n815), .A2(KEYINPUT121), .A3(KEYINPUT54), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n508), .B(KEYINPUT57), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n652), .B(KEYINPUT122), .Z(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n815), .A2(G902), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n878), .A2(new_n749), .A3(new_n747), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n856), .B1(new_n877), .B2(new_n879), .ZN(G54));
  NAND3_X1  g694(.A1(new_n878), .A2(KEYINPUT58), .A3(G475), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(new_n402), .Z(new_n882));
  NOR2_X1   g696(.A1(new_n882), .A2(new_n856), .ZN(G60));
  NAND2_X1  g697(.A1(G478), .A2(G902), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT59), .ZN(new_n885));
  AND4_X1   g699(.A1(new_n582), .A2(new_n872), .A3(new_n873), .A4(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n582), .B1(new_n822), .B2(new_n885), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n886), .A2(new_n856), .A3(new_n887), .ZN(G63));
  NAND2_X1  g702(.A1(G217), .A2(G902), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(KEYINPUT60), .Z(new_n890));
  NAND2_X1  g704(.A1(new_n815), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n856), .B1(new_n891), .B2(new_n343), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT123), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n815), .A2(new_n601), .A3(new_n890), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n893), .B1(new_n892), .B2(new_n894), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT61), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n891), .A2(new_n343), .ZN(new_n899));
  INV_X1    g713(.A(new_n856), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n899), .A2(new_n900), .A3(new_n894), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT123), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT61), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n898), .A2(new_n904), .ZN(G66));
  AND2_X1   g719(.A1(new_n791), .A2(new_n786), .ZN(new_n906));
  INV_X1    g720(.A(new_n339), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT124), .ZN(new_n909));
  OAI21_X1  g723(.A(G953), .B1(new_n464), .B2(new_n533), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n862), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n912), .B1(G898), .B2(new_n339), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n911), .B(new_n913), .ZN(G69));
  NAND2_X1  g728(.A1(new_n251), .A2(new_n259), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(new_n389), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n773), .A2(new_n762), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n771), .A2(new_n632), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n587), .A2(new_n783), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n651), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(KEYINPUT125), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n642), .A2(new_n804), .A3(new_n649), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT62), .Z(new_n924));
  OR2_X1    g738(.A1(new_n921), .A2(KEYINPUT125), .ZN(new_n925));
  AND4_X1   g739(.A1(new_n918), .A2(new_n922), .A3(new_n924), .A4(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n917), .B1(new_n926), .B2(new_n907), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(KEYINPUT126), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT126), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n929), .B(new_n917), .C1(new_n926), .C2(new_n907), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n757), .A2(new_n631), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n692), .A2(new_n351), .A3(new_n732), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n795), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n811), .B(KEYINPUT127), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n918), .A2(new_n339), .A3(new_n933), .A4(new_n934), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n935), .B(new_n916), .C1(new_n611), .C2(new_n339), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n928), .A2(new_n930), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n339), .B1(G227), .B2(G900), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n938), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n928), .A2(new_n930), .A3(new_n940), .A4(new_n936), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n939), .A2(new_n941), .ZN(G72));
  NAND2_X1  g756(.A1(new_n260), .A2(new_n262), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n271), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n926), .A2(new_n906), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n621), .B(KEYINPUT63), .Z(new_n946));
  AOI21_X1  g760(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n918), .A2(new_n906), .A3(new_n933), .A4(new_n934), .ZN(new_n948));
  AOI211_X1 g762(.A(new_n271), .B(new_n943), .C1(new_n948), .C2(new_n946), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n819), .A2(new_n820), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n943), .A2(new_n271), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n944), .A2(new_n946), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NOR4_X1   g767(.A1(new_n947), .A2(new_n949), .A3(new_n856), .A4(new_n953), .ZN(G57));
endmodule


